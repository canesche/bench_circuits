module top ( clock, 
    pcount_3_, pkey_5_, pkey_131_, pkey_144_, pkey_157_, pkey_230_,
    pkey_243_, pcount_2_, pkey_4_, pkey_132_, pkey_158_, pkey_169_,
    pkey_242_, pcount_1_, pkey_146_, pkey_168_, pkey_245_, pcount_0_,
    pkey_6_, pkey_130_, pkey_145_, pkey_244_, pkey_9_, pkey_16_, pkey_27_,
    pkey_38_, pkey_49_, pkey_122_, pkey_148_, pkey_153_, pkey_166_,
    pkey_221_, pkey_252_, pkey_8_, pkey_17_, pkey_26_, pkey_48_, pkey_110_,
    pkey_121_, pkey_147_, pkey_154_, pkey_165_, pkey_220_, pkey_246_,
    pkey_253_, pkey_18_, pkey_29_, pkey_36_, pkey_120_, pkey_155_,
    pkey_164_, pkey_210_, pkey_249_, pkey_254_, pkey_19_, pkey_28_,
    pkey_37_, pkey_46_, pkey_112_, pkey_149_, pkey_156_, pkey_163_,
    pkey_211_, pkey_248_, pkey_56_, pkey_67_, pkey_78_, pkey_89_,
    pkey_113_, pkey_126_, pkey_139_, pkey_162_, pkey_212_, pkey_225_,
    pkey_238_, pkey_57_, pkey_66_, pkey_88_, pkey_114_, pkey_125_,
    pkey_150_, pkey_161_, pkey_213_, pkey_224_, pkey_58_, pkey_69_,
    pkey_76_, pkey_115_, pkey_124_, pkey_137_, pkey_160_, pkey_214_,
    pkey_250_, pkey_59_, pkey_68_, pkey_77_, pkey_86_, pkey_116_,
    pkey_123_, pkey_138_, pkey_152_, pkey_222_, pkey_237_, pkey_251_,
    pkey_1_, pkey_96_, pkey_117_, pkey_140_, pkey_216_, pkey_229_,
    pkey_234_, pkey_0_, pkey_97_, pkey_118_, pkey_129_, pkey_136_,
    pkey_217_, pkey_228_, pkey_235_, pkey_3_, pkey_98_, pkey_128_,
    pkey_133_, pkey_142_, pkey_218_, pkey_227_, pkey_232_, pkey_241_,
    pkey_2_, pkey_99_, pkey_134_, pkey_141_, pkey_219_, pkey_226_,
    pkey_233_, pkey_240_, pkey_70_, pkey_81_, pkey_92_, pkey_180_,
    pkey_193_, pkey_80_, pkey_93_, pkey_107_, pkey_194_, pkey_206_, pclk,
    pkey_50_, pkey_61_, pkey_94_, pkey_182_, pkey_195_, pkey_209_,
    pstart_0_, pkey_51_, pkey_60_, pkey_109_, pkey_181_, pkey_196_,
    pkey_208_, pkey_52_, pkey_74_, pkey_85_, pkey_104_, pkey_171_,
    pkey_197_, pkey_203_, pencrypt_0_, pkey_53_, pkey_62_, pkey_75_,
    pkey_84_, pkey_172_, pkey_198_, pkey_202_, pkey_54_, pkey_65_,
    pkey_72_, pkey_83_, pkey_90_, pkey_106_, pkey_205_, pkey_64_, pkey_73_,
    pkey_82_, pkey_91_, pkey_105_, pkey_170_, pkey_204_, pkey_12_,
    pkey_34_, pkey_45_, pkey_100_, pkey_188_, pkey_13_, pkey_22_, pkey_35_,
    pkey_44_, pkey_176_, pkey_187_, pkey_14_, pkey_25_, pkey_32_, pkey_43_,
    pkey_102_, pkey_173_, pkey_201_, pkey_24_, pkey_33_, pkey_42_,
    pkey_101_, pkey_174_, pkey_189_, pkey_200_, pkey_30_, pkey_41_,
    pkey_179_, pkey_184_, pkey_40_, pkey_190_, pkey_10_, pkey_21_,
    pkey_177_, pkey_186_, pkey_11_, pkey_20_, pkey_178_, pkey_185_,
    pkey_192_,
    pksi_50_, pksi_61_, pksi_72_, pksi_83_, pksi_94_, pksi_102_, pksi_115_,
    pksi_128_, pdata_ready_0_, pksi_51_, pksi_60_, pksi_73_, pksi_82_,
    pksi_95_, pksi_101_, pksi_116_, pksi_127_, pksi_52_, pksi_63_,
    pksi_70_, pksi_81_, pksi_96_, pksi_100_, pksi_113_, pksi_53_, pksi_62_,
    pksi_71_, pksi_80_, pksi_97_, pksi_114_, pksi_129_, pksi_54_, pksi_65_,
    pksi_76_, pksi_87_, pksi_90_, pksi_119_, pksi_124_, pksi_191_,
    pksi_55_, pksi_64_, pksi_77_, pksi_86_, pksi_91_, pksi_123_, pksi_56_,
    pksi_67_, pksi_74_, pksi_85_, pksi_92_, pksi_117_, pksi_126_, pksi_57_,
    pksi_66_, pksi_75_, pksi_84_, pksi_93_, pksi_118_, pksi_125_,
    pksi_190_, pksi_14_, pksi_25_, pksi_36_, pksi_47_, pksi_120_, pksi_15_,
    pksi_24_, pksi_37_, pksi_46_, pksi_109_, pnew_count_3_, pksi_16_,
    pksi_27_, pksi_34_, pksi_45_, pksi_108_, pksi_122_, pksi_17_, pksi_26_,
    pksi_35_, pksi_44_, pksi_107_, pksi_121_, pksi_10_, pksi_21_, pksi_32_,
    pksi_43_, pksi_106_, pksi_111_, pnew_count_0_, pksi_11_, pksi_20_,
    pksi_33_, pksi_42_, pksi_105_, pksi_112_, pksi_12_, pksi_23_, pksi_30_,
    pksi_41_, pksi_104_, pnew_count_2_, pksi_13_, pksi_22_, pksi_31_,
    pksi_40_, pksi_103_, pksi_110_, pnew_count_1_, pksi_3_, pksi_151_,
    pksi_164_, pksi_177_, pksi_2_, pksi_152_, pksi_163_, pksi_178_,
    pksi_189_, pksi_1_, pksi_166_, pksi_179_, pksi_188_, pksi_0_,
    pksi_150_, pksi_165_, pksi_187_, pksi_18_, pksi_29_, pksi_142_,
    pksi_168_, pksi_173_, pksi_186_, pksi_19_, pksi_28_, pksi_130_,
    pksi_141_, pksi_167_, pksi_174_, pksi_185_, pksi_38_, pksi_49_,
    pksi_131_, pksi_140_, pksi_175_, pksi_184_, pksi_39_, pksi_48_,
    pksi_132_, pksi_169_, pksi_176_, pksi_183_, pksi_58_, pksi_69_,
    pksi_133_, pksi_146_, pksi_159_, pksi_182_, pksi_59_, pksi_68_,
    pksi_134_, pksi_145_, pksi_170_, pksi_181_, pksi_9_, pksi_78_,
    pksi_89_, pksi_135_, pksi_144_, pksi_157_, pksi_171_, pksi_180_,
    pksi_8_, pksi_79_, pksi_88_, pksi_136_, pksi_143_, pksi_158_,
    pksi_172_, pksi_7_, pksi_98_, pksi_137_, pksi_155_, pksi_160_, pksi_6_,
    pksi_99_, pksi_138_, pksi_149_, pksi_156_, pksi_5_, pksi_139_,
    pksi_148_, pksi_153_, pksi_162_, pksi_4_, pksi_147_, pksi_154_,
    pksi_161_  );
  input  clock;
  input  pcount_3_, pkey_5_, pkey_131_, pkey_144_, pkey_157_, pkey_230_,
    pkey_243_, pcount_2_, pkey_4_, pkey_132_, pkey_158_, pkey_169_,
    pkey_242_, pcount_1_, pkey_146_, pkey_168_, pkey_245_, pcount_0_,
    pkey_6_, pkey_130_, pkey_145_, pkey_244_, pkey_9_, pkey_16_, pkey_27_,
    pkey_38_, pkey_49_, pkey_122_, pkey_148_, pkey_153_, pkey_166_,
    pkey_221_, pkey_252_, pkey_8_, pkey_17_, pkey_26_, pkey_48_, pkey_110_,
    pkey_121_, pkey_147_, pkey_154_, pkey_165_, pkey_220_, pkey_246_,
    pkey_253_, pkey_18_, pkey_29_, pkey_36_, pkey_120_, pkey_155_,
    pkey_164_, pkey_210_, pkey_249_, pkey_254_, pkey_19_, pkey_28_,
    pkey_37_, pkey_46_, pkey_112_, pkey_149_, pkey_156_, pkey_163_,
    pkey_211_, pkey_248_, pkey_56_, pkey_67_, pkey_78_, pkey_89_,
    pkey_113_, pkey_126_, pkey_139_, pkey_162_, pkey_212_, pkey_225_,
    pkey_238_, pkey_57_, pkey_66_, pkey_88_, pkey_114_, pkey_125_,
    pkey_150_, pkey_161_, pkey_213_, pkey_224_, pkey_58_, pkey_69_,
    pkey_76_, pkey_115_, pkey_124_, pkey_137_, pkey_160_, pkey_214_,
    pkey_250_, pkey_59_, pkey_68_, pkey_77_, pkey_86_, pkey_116_,
    pkey_123_, pkey_138_, pkey_152_, pkey_222_, pkey_237_, pkey_251_,
    pkey_1_, pkey_96_, pkey_117_, pkey_140_, pkey_216_, pkey_229_,
    pkey_234_, pkey_0_, pkey_97_, pkey_118_, pkey_129_, pkey_136_,
    pkey_217_, pkey_228_, pkey_235_, pkey_3_, pkey_98_, pkey_128_,
    pkey_133_, pkey_142_, pkey_218_, pkey_227_, pkey_232_, pkey_241_,
    pkey_2_, pkey_99_, pkey_134_, pkey_141_, pkey_219_, pkey_226_,
    pkey_233_, pkey_240_, pkey_70_, pkey_81_, pkey_92_, pkey_180_,
    pkey_193_, pkey_80_, pkey_93_, pkey_107_, pkey_194_, pkey_206_, pclk,
    pkey_50_, pkey_61_, pkey_94_, pkey_182_, pkey_195_, pkey_209_,
    pstart_0_, pkey_51_, pkey_60_, pkey_109_, pkey_181_, pkey_196_,
    pkey_208_, pkey_52_, pkey_74_, pkey_85_, pkey_104_, pkey_171_,
    pkey_197_, pkey_203_, pencrypt_0_, pkey_53_, pkey_62_, pkey_75_,
    pkey_84_, pkey_172_, pkey_198_, pkey_202_, pkey_54_, pkey_65_,
    pkey_72_, pkey_83_, pkey_90_, pkey_106_, pkey_205_, pkey_64_, pkey_73_,
    pkey_82_, pkey_91_, pkey_105_, pkey_170_, pkey_204_, pkey_12_,
    pkey_34_, pkey_45_, pkey_100_, pkey_188_, pkey_13_, pkey_22_, pkey_35_,
    pkey_44_, pkey_176_, pkey_187_, pkey_14_, pkey_25_, pkey_32_, pkey_43_,
    pkey_102_, pkey_173_, pkey_201_, pkey_24_, pkey_33_, pkey_42_,
    pkey_101_, pkey_174_, pkey_189_, pkey_200_, pkey_30_, pkey_41_,
    pkey_179_, pkey_184_, pkey_40_, pkey_190_, pkey_10_, pkey_21_,
    pkey_177_, pkey_186_, pkey_11_, pkey_20_, pkey_178_, pkey_185_,
    pkey_192_;
  output pksi_50_, pksi_61_, pksi_72_, pksi_83_, pksi_94_, pksi_102_,
    pksi_115_, pksi_128_, pdata_ready_0_, pksi_51_, pksi_60_, pksi_73_,
    pksi_82_, pksi_95_, pksi_101_, pksi_116_, pksi_127_, pksi_52_,
    pksi_63_, pksi_70_, pksi_81_, pksi_96_, pksi_100_, pksi_113_, pksi_53_,
    pksi_62_, pksi_71_, pksi_80_, pksi_97_, pksi_114_, pksi_129_, pksi_54_,
    pksi_65_, pksi_76_, pksi_87_, pksi_90_, pksi_119_, pksi_124_,
    pksi_191_, pksi_55_, pksi_64_, pksi_77_, pksi_86_, pksi_91_, pksi_123_,
    pksi_56_, pksi_67_, pksi_74_, pksi_85_, pksi_92_, pksi_117_, pksi_126_,
    pksi_57_, pksi_66_, pksi_75_, pksi_84_, pksi_93_, pksi_118_, pksi_125_,
    pksi_190_, pksi_14_, pksi_25_, pksi_36_, pksi_47_, pksi_120_, pksi_15_,
    pksi_24_, pksi_37_, pksi_46_, pksi_109_, pnew_count_3_, pksi_16_,
    pksi_27_, pksi_34_, pksi_45_, pksi_108_, pksi_122_, pksi_17_, pksi_26_,
    pksi_35_, pksi_44_, pksi_107_, pksi_121_, pksi_10_, pksi_21_, pksi_32_,
    pksi_43_, pksi_106_, pksi_111_, pnew_count_0_, pksi_11_, pksi_20_,
    pksi_33_, pksi_42_, pksi_105_, pksi_112_, pksi_12_, pksi_23_, pksi_30_,
    pksi_41_, pksi_104_, pnew_count_2_, pksi_13_, pksi_22_, pksi_31_,
    pksi_40_, pksi_103_, pksi_110_, pnew_count_1_, pksi_3_, pksi_151_,
    pksi_164_, pksi_177_, pksi_2_, pksi_152_, pksi_163_, pksi_178_,
    pksi_189_, pksi_1_, pksi_166_, pksi_179_, pksi_188_, pksi_0_,
    pksi_150_, pksi_165_, pksi_187_, pksi_18_, pksi_29_, pksi_142_,
    pksi_168_, pksi_173_, pksi_186_, pksi_19_, pksi_28_, pksi_130_,
    pksi_141_, pksi_167_, pksi_174_, pksi_185_, pksi_38_, pksi_49_,
    pksi_131_, pksi_140_, pksi_175_, pksi_184_, pksi_39_, pksi_48_,
    pksi_132_, pksi_169_, pksi_176_, pksi_183_, pksi_58_, pksi_69_,
    pksi_133_, pksi_146_, pksi_159_, pksi_182_, pksi_59_, pksi_68_,
    pksi_134_, pksi_145_, pksi_170_, pksi_181_, pksi_9_, pksi_78_,
    pksi_89_, pksi_135_, pksi_144_, pksi_157_, pksi_171_, pksi_180_,
    pksi_8_, pksi_79_, pksi_88_, pksi_136_, pksi_143_, pksi_158_,
    pksi_172_, pksi_7_, pksi_98_, pksi_137_, pksi_155_, pksi_160_, pksi_6_,
    pksi_99_, pksi_138_, pksi_149_, pksi_156_, pksi_5_, pksi_139_,
    pksi_148_, pksi_153_, pksi_162_, pksi_4_, pksi_147_, pksi_154_,
    pksi_161_;
  reg n_n95, n_n105, n_n2410, n_n122, n_n132, n_n141, n_n178, n_n2513,
    n_n96, n_n2396, n_n2412, n_n121, n_n133, n_n2448, n_n179, n_n187,
    n_n97, n_n107, n_n114, n_n120, n_n149, n_n159, n_n180, n_n189, n_n195,
    n_n98, n_n106, n_n2408, n_n119, n_n150, n_n158, n_n181, n_n188, n_n15,
    n_n92, n_n102, n_n112, n_n2420, n_n165, n_n174, n_n184, n_n193, n_n93,
    n_n101, n_n113, n_n118, n_n2485, n_n2495, n_n175, n_n194, n_n94,
    n_n104, n_n110, n_n117, n_n176, n_n186, n_n2384, n_n103, n_n111,
    n_n2416, n_n177, n_n185, n_n192, n_n12, n_n125, n_n2440, n_n143,
    n_n153, n_n162, n_n171, n_n2272, n_n126, n_n134, n_n144, n_n152,
    n_n163, n_n170, n_n13, n_n2430, n_n136, n_n142, n_n151, n_n2481,
    n_n173, n_n14, n_n127, n_n135, n_n2452, n_n2462, n_n164, n_n172, n_n9,
    n_n99, n_n109, n_n128, n_n138, n_n147, n_n157, n_n160, n_n167, n_n182,
    n_n190, n_n10, n_n100, n_n108, n_n129, n_n137, n_n148, n_n156, n_n2474,
    n_n166, n_n183, n_n2517, n_n2268, n_n115, n_n124, n_n130, n_n140,
    n_n145, n_n155, n_n2476, n_n169, n_n2507, n_n11, n_n116, n_n123,
    n_n131, n_n139, n_n146, n_n154, n_n161, n_n168, n_n191, n_n49, n_n59,
    n_n68, n_n78, n_n2374, n_n50, n_n58, n_n69, n_n77, n_n87, n_n51, n_n60,
    n_n66, n_n76, n_n88, n_n8, n_n52, n_n2337, n_n67, n_n75, n_n89,
    n_n2277, n_n24, n_n34, n_n43, n_n90, n_n16, n_n23, n_n35, n_n42, n_n91,
    n_n2280, n_n26, n_n33, n_n41, n_n17, n_n25, n_n2301, n_n40, n_n18,
    n_n28, n_n37, n_n2320, n_n57, n_n65, n_n19, n_n27, n_n38, n_n46,
    n_n2333, n_n64, n_n20, n_n30, n_n2305, n_n45, n_n73, n_n83, n_n21,
    n_n29, n_n36, n_n44, n_n74, n_n82, n_n22, n_n32, n_n53, n_n62, n_n71,
    n_n2365, n_n2369, n_n2288, n_n31, n_n54, n_n61, n_n72, n_n81, n_n84,
    n_n2310, n_n48, n_n55, n_n63, n_n70, n_n80, n_n85, n_n39, n_n47, n_n56,
    n_n2342, n_n2352, n_n79, n_n86;
  wire new_n1099_1_, new_n1100_, new_n1101_, new_n1102_, new_n1103_,
    new_n1104_1_, new_n1105_, new_n1106_, new_n1107_, new_n1108_,
    new_n1109_1_, new_n1110_, new_n1111_, new_n1112_, new_n1113_,
    new_n1114_1_, new_n1115_, new_n1116_, new_n1117_, new_n1118_,
    new_n1119_1_, new_n1120_, new_n1121_, new_n1122_, new_n1123_,
    new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_1_,
    new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_1_,
    new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1140_, new_n1142_,
    new_n1143_, new_n1144_1_, new_n1145_, new_n1146_, new_n1147_,
    new_n1148_, new_n1150_, new_n1151_, new_n1152_, new_n1153_,
    new_n1154_1_, new_n1155_, new_n1157_, new_n1158_, new_n1159_1_,
    new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_1_,
    new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_1_,
    new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_1_,
    new_n1176_, new_n1177_, new_n1178_, new_n1179_1_, new_n1180_,
    new_n1181_, new_n1182_, new_n1183_, new_n1184_1_, new_n1185_,
    new_n1187_, new_n1188_, new_n1189_1_, new_n1190_, new_n1191_,
    new_n1192_, new_n1193_, new_n1194_1_, new_n1195_, new_n1196_,
    new_n1198_, new_n1199_1_, new_n1200_, new_n1201_, new_n1202_,
    new_n1203_, new_n1204_1_, new_n1205_, new_n1206_, new_n1207_,
    new_n1209_1_, new_n1210_, new_n1211_, new_n1212_, new_n1213_,
    new_n1214_1_, new_n1215_, new_n1216_, new_n1217_, new_n1218_,
    new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_1_,
    new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_1_,
    new_n1231_, new_n1232_, new_n1233_, new_n1234_1_, new_n1235_,
    new_n1236_, new_n1237_, new_n1238_, new_n1239_1_, new_n1240_,
    new_n1242_, new_n1243_, new_n1244_1_, new_n1245_, new_n1246_,
    new_n1247_, new_n1248_, new_n1249_1_, new_n1250_, new_n1251_,
    new_n1253_, new_n1254_1_, new_n1255_, new_n1256_, new_n1257_,
    new_n1258_, new_n1259_1_, new_n1260_, new_n1261_, new_n1262_,
    new_n1264_1_, new_n1265_, new_n1266_, new_n1267_, new_n1268_,
    new_n1269_1_, new_n1270_, new_n1271_, new_n1272_, new_n1273_,
    new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_1_,
    new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_1_,
    new_n1286_, new_n1287_, new_n1288_, new_n1289_1_, new_n1290_,
    new_n1291_, new_n1292_, new_n1293_, new_n1294_1_, new_n1295_,
    new_n1297_, new_n1298_, new_n1299_1_, new_n1300_, new_n1301_,
    new_n1302_, new_n1303_, new_n1304_1_, new_n1305_, new_n1306_,
    new_n1308_, new_n1309_1_, new_n1310_, new_n1311_, new_n1312_,
    new_n1313_, new_n1314_1_, new_n1315_, new_n1316_, new_n1317_,
    new_n1319_1_, new_n1320_, new_n1321_, new_n1322_, new_n1323_,
    new_n1324_1_, new_n1325_, new_n1326_, new_n1327_, new_n1328_,
    new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_1_,
    new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1339_1_,
    new_n1341_, new_n1342_, new_n1343_, new_n1344_1_, new_n1345_,
    new_n1346_, new_n1347_, new_n1348_, new_n1349_1_, new_n1350_,
    new_n1352_, new_n1353_, new_n1354_1_, new_n1355_, new_n1356_,
    new_n1357_, new_n1358_, new_n1359_1_, new_n1360_, new_n1361_,
    new_n1363_, new_n1364_1_, new_n1365_, new_n1366_, new_n1367_,
    new_n1368_, new_n1369_1_, new_n1370_, new_n1371_, new_n1372_,
    new_n1374_1_, new_n1375_, new_n1376_, new_n1377_, new_n1378_,
    new_n1379_1_, new_n1380_, new_n1381_, new_n1382_, new_n1383_,
    new_n1385_, new_n1386_, new_n1387_, new_n1388_, new_n1389_1_,
    new_n1390_, new_n1391_, new_n1392_, new_n1393_, new_n1394_1_,
    new_n1396_, new_n1397_, new_n1398_, new_n1399_1_, new_n1400_,
    new_n1401_, new_n1402_, new_n1403_, new_n1404_1_, new_n1405_,
    new_n1407_, new_n1408_, new_n1409_1_, new_n1410_, new_n1411_,
    new_n1412_, new_n1413_, new_n1414_1_, new_n1415_, new_n1416_,
    new_n1418_, new_n1419_1_, new_n1420_, new_n1421_, new_n1422_,
    new_n1423_, new_n1424_1_, new_n1425_, new_n1426_, new_n1427_,
    new_n1429_1_, new_n1430_, new_n1431_, new_n1432_, new_n1433_,
    new_n1434_1_, new_n1435_, new_n1436_, new_n1437_, new_n1438_,
    new_n1440_, new_n1441_, new_n1442_, new_n1443_, new_n1444_1_,
    new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_1_,
    new_n1451_, new_n1452_, new_n1453_, new_n1454_1_, new_n1455_,
    new_n1456_, new_n1457_, new_n1458_, new_n1459_1_, new_n1460_,
    new_n1462_, new_n1463_, new_n1464_1_, new_n1465_, new_n1466_,
    new_n1467_, new_n1468_, new_n1469_1_, new_n1470_, new_n1471_,
    new_n1473_, new_n1474_1_, new_n1475_, new_n1476_, new_n1477_,
    new_n1478_, new_n1479_1_, new_n1480_, new_n1481_, new_n1482_,
    new_n1484_1_, new_n1485_, new_n1486_, new_n1487_, new_n1488_,
    new_n1489_1_, new_n1490_, new_n1491_, new_n1492_, new_n1493_,
    new_n1495_, new_n1496_, new_n1497_, new_n1498_, new_n1499_1_,
    new_n1500_, new_n1501_, new_n1502_, new_n1503_, new_n1504_1_,
    new_n1506_, new_n1507_, new_n1508_, new_n1509_1_, new_n1510_,
    new_n1511_, new_n1512_, new_n1513_, new_n1514_1_, new_n1516_,
    new_n1517_, new_n1518_, new_n1519_1_, new_n1520_, new_n1521_,
    new_n1522_, new_n1523_, new_n1524_1_, new_n1525_, new_n1527_,
    new_n1528_, new_n1529_1_, new_n1530_, new_n1531_, new_n1532_,
    new_n1533_, new_n1534_1_, new_n1535_, new_n1536_, new_n1538_,
    new_n1539_1_, new_n1540_, new_n1541_, new_n1542_, new_n1543_,
    new_n1544_1_, new_n1545_, new_n1546_, new_n1547_, new_n1549_1_,
    new_n1550_, new_n1551_, new_n1552_, new_n1553_, new_n1554_1_,
    new_n1555_, new_n1556_, new_n1557_, new_n1558_, new_n1560_, new_n1561_,
    new_n1562_, new_n1563_, new_n1564_1_, new_n1565_, new_n1566_,
    new_n1567_, new_n1568_, new_n1569_1_, new_n1571_, new_n1572_,
    new_n1573_, new_n1574_1_, new_n1575_, new_n1576_, new_n1577_,
    new_n1578_, new_n1579_1_, new_n1580_, new_n1582_, new_n1583_,
    new_n1584_1_, new_n1585_, new_n1586_, new_n1587_, new_n1588_,
    new_n1589_1_, new_n1590_, new_n1591_, new_n1593_, new_n1594_1_,
    new_n1595_, new_n1596_, new_n1597_, new_n1598_, new_n1599_1_,
    new_n1600_, new_n1601_, new_n1602_, new_n1604_1_, new_n1605_,
    new_n1606_, new_n1607_, new_n1608_, new_n1609_1_, new_n1610_,
    new_n1611_, new_n1612_, new_n1613_, new_n1615_, new_n1616_, new_n1617_,
    new_n1618_, new_n1619_1_, new_n1620_, new_n1621_, new_n1622_,
    new_n1623_, new_n1624_1_, new_n1626_, new_n1627_, new_n1628_,
    new_n1629_1_, new_n1630_, new_n1631_, new_n1632_, new_n1633_,
    new_n1634_1_, new_n1635_, new_n1637_, new_n1638_, new_n1639_1_,
    new_n1640_, new_n1641_, new_n1642_, new_n1643_, new_n1644_1_,
    new_n1645_, new_n1646_, new_n1648_, new_n1649_1_, new_n1650_,
    new_n1651_, new_n1652_, new_n1653_, new_n1654_1_, new_n1655_,
    new_n1656_, new_n1657_, new_n1659_1_, new_n1660_, new_n1661_,
    new_n1662_, new_n1663_, new_n1664_1_, new_n1665_, new_n1666_,
    new_n1667_, new_n1668_, new_n1670_, new_n1671_, new_n1672_, new_n1673_,
    new_n1674_1_, new_n1675_, new_n1676_, new_n1677_, new_n1678_,
    new_n1679_1_, new_n1681_, new_n1682_, new_n1683_, new_n1684_1_,
    new_n1685_, new_n1686_, new_n1687_, new_n1688_, new_n1689_1_,
    new_n1690_, new_n1692_, new_n1693_, new_n1694_1_, new_n1695_,
    new_n1696_, new_n1697_, new_n1698_, new_n1699_1_, new_n1700_,
    new_n1701_, new_n1703_, new_n1704_1_, new_n1705_, new_n1706_,
    new_n1707_, new_n1708_, new_n1709_1_, new_n1710_, new_n1711_,
    new_n1712_, new_n1714_1_, new_n1715_, new_n1716_, new_n1717_,
    new_n1718_, new_n1719_1_, new_n1720_, new_n1721_, new_n1722_,
    new_n1723_, new_n1725_, new_n1726_, new_n1727_, new_n1728_,
    new_n1729_1_, new_n1730_, new_n1731_, new_n1732_, new_n1733_,
    new_n1734_1_, new_n1736_, new_n1737_, new_n1738_, new_n1739_1_,
    new_n1740_, new_n1741_, new_n1742_, new_n1743_, new_n1744_1_,
    new_n1745_, new_n1747_, new_n1748_, new_n1749_1_, new_n1750_,
    new_n1751_, new_n1752_, new_n1753_, new_n1754_1_, new_n1755_,
    new_n1756_, new_n1758_, new_n1759_1_, new_n1760_, new_n1761_,
    new_n1762_, new_n1763_, new_n1764_1_, new_n1765_, new_n1766_,
    new_n1767_, new_n1769_1_, new_n1770_, new_n1771_, new_n1772_,
    new_n1773_, new_n1774_1_, new_n1775_, new_n1776_, new_n1777_,
    new_n1778_, new_n1780_, new_n1781_, new_n1782_, new_n1783_,
    new_n1784_1_, new_n1785_, new_n1786_, new_n1787_, new_n1788_,
    new_n1789_1_, new_n1791_, new_n1792_, new_n1793_, new_n1794_1_,
    new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1799_1_,
    new_n1800_, new_n1802_, new_n1803_, new_n1804_1_, new_n1805_,
    new_n1806_, new_n1807_, new_n1808_, new_n1809_1_, new_n1810_,
    new_n1812_, new_n1813_, new_n1814_1_, new_n1815_, new_n1816_,
    new_n1817_, new_n1818_, new_n1819_1_, new_n1820_, new_n1821_,
    new_n1823_, new_n1824_1_, new_n1825_, new_n1826_, new_n1827_,
    new_n1828_, new_n1829_1_, new_n1830_, new_n1831_, new_n1832_,
    new_n1834_1_, new_n1835_, new_n1836_, new_n1837_, new_n1838_,
    new_n1839_1_, new_n1840_, new_n1841_, new_n1842_, new_n1843_,
    new_n1845_, new_n1846_, new_n1847_, new_n1848_, new_n1849_1_,
    new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1854_1_,
    new_n1856_, new_n1857_, new_n1858_, new_n1859_1_, new_n1860_,
    new_n1861_, new_n1862_, new_n1863_, new_n1864_1_, new_n1865_,
    new_n1867_, new_n1868_, new_n1869_1_, new_n1870_, new_n1871_,
    new_n1872_, new_n1873_, new_n1874_1_, new_n1875_, new_n1876_,
    new_n1878_, new_n1879_1_, new_n1880_, new_n1881_, new_n1882_,
    new_n1883_, new_n1884_1_, new_n1885_, new_n1886_, new_n1887_,
    new_n1889_1_, new_n1890_, new_n1891_, new_n1892_, new_n1893_,
    new_n1894_1_, new_n1895_, new_n1896_, new_n1897_, new_n1898_,
    new_n1900_, new_n1901_, new_n1902_, new_n1903_, new_n1904_1_,
    new_n1905_, new_n1906_, new_n1907_, new_n1908_, new_n1909_1_,
    new_n1911_, new_n1912_, new_n1913_, new_n1914_1_, new_n1915_,
    new_n1916_, new_n1917_, new_n1918_, new_n1919_1_, new_n1920_,
    new_n1922_, new_n1923_, new_n1924_1_, new_n1925_, new_n1926_,
    new_n1927_, new_n1928_, new_n1929_1_, new_n1930_, new_n1931_,
    new_n1933_, new_n1934_1_, new_n1935_, new_n1936_, new_n1937_,
    new_n1938_, new_n1939_1_, new_n1940_, new_n1941_, new_n1942_,
    new_n1944_1_, new_n1945_, new_n1946_, new_n1947_, new_n1948_,
    new_n1949_1_, new_n1950_, new_n1951_, new_n1952_, new_n1953_,
    new_n1955_, new_n1956_, new_n1957_, new_n1958_, new_n1959_1_,
    new_n1960_, new_n1961_, new_n1962_, new_n1963_, new_n1965_, new_n1966_,
    new_n1967_, new_n1968_, new_n1969_1_, new_n1970_, new_n1971_,
    new_n1972_, new_n1973_, new_n1974_, new_n1976_, new_n1977_, new_n1978_,
    new_n1979_, new_n1980_, new_n1981_, new_n1982_, new_n1983_, new_n1984_,
    new_n1985_, new_n1987_, new_n1988_, new_n1989_, new_n1990_, new_n1991_,
    new_n1992_, new_n1993_, new_n1994_, new_n1995_, new_n1996_, new_n1998_,
    new_n1999_, new_n2000_, new_n2001_, new_n2002_, new_n2003_, new_n2004_,
    new_n2005_, new_n2006_, new_n2007_, new_n2009_, new_n2010_, new_n2011_,
    new_n2012_, new_n2013_, new_n2014_, new_n2015_, new_n2016_, new_n2017_,
    new_n2018_, new_n2020_, new_n2021_, new_n2022_, new_n2023_, new_n2024_,
    new_n2025_, new_n2026_, new_n2027_, new_n2028_, new_n2029_, new_n2031_,
    new_n2032_, new_n2033_, new_n2034_, new_n2035_, new_n2036_, new_n2037_,
    new_n2038_, new_n2039_, new_n2040_, new_n2042_, new_n2043_, new_n2044_,
    new_n2045_, new_n2046_, new_n2047_, new_n2048_, new_n2049_, new_n2050_,
    new_n2051_, new_n2053_, new_n2054_, new_n2055_, new_n2056_, new_n2057_,
    new_n2058_, new_n2059_, new_n2060_, new_n2061_, new_n2062_, new_n2064_,
    new_n2065_, new_n2066_, new_n2067_, new_n2068_, new_n2069_, new_n2070_,
    new_n2071_, new_n2072_, new_n2073_, new_n2075_, new_n2076_, new_n2077_,
    new_n2078_, new_n2079_, new_n2080_, new_n2081_, new_n2082_, new_n2083_,
    new_n2084_, new_n2086_, new_n2087_, new_n2088_, new_n2089_, new_n2090_,
    new_n2091_, new_n2092_, new_n2093_, new_n2094_, new_n2095_, new_n2097_,
    new_n2098_, new_n2099_, new_n2100_, new_n2101_, new_n2102_, new_n2103_,
    new_n2104_, new_n2105_, new_n2106_, new_n2108_, new_n2109_, new_n2110_,
    new_n2111_, new_n2112_, new_n2113_, new_n2114_, new_n2115_, new_n2116_,
    new_n2117_, new_n2119_, new_n2120_, new_n2121_, new_n2122_, new_n2123_,
    new_n2124_, new_n2125_, new_n2126_, new_n2127_, new_n2128_, new_n2130_,
    new_n2131_, new_n2132_, new_n2133_, new_n2134_, new_n2135_, new_n2136_,
    new_n2137_, new_n2138_, new_n2139_, new_n2141_, new_n2142_, new_n2143_,
    new_n2144_, new_n2145_, new_n2146_, new_n2147_, new_n2148_, new_n2149_,
    new_n2150_, new_n2152_, new_n2153_, new_n2154_, new_n2155_, new_n2156_,
    new_n2157_, new_n2158_, new_n2159_, new_n2160_, new_n2161_, new_n2163_,
    new_n2164_, new_n2165_, new_n2166_, new_n2167_, new_n2168_, new_n2169_,
    new_n2170_, new_n2171_, new_n2172_, new_n2174_, new_n2175_, new_n2176_,
    new_n2177_, new_n2178_, new_n2179_, new_n2180_, new_n2181_, new_n2182_,
    new_n2183_, new_n2185_, new_n2186_, new_n2187_, new_n2188_, new_n2189_,
    new_n2190_, new_n2191_, new_n2192_, new_n2193_, new_n2194_, new_n2196_,
    new_n2197_, new_n2198_, new_n2199_, new_n2200_, new_n2201_, new_n2202_,
    new_n2203_, new_n2204_, new_n2205_, new_n2207_, new_n2208_, new_n2209_,
    new_n2210_, new_n2211_, new_n2212_, new_n2213_, new_n2214_, new_n2215_,
    new_n2216_, new_n2218_, new_n2219_, new_n2220_, new_n2221_, new_n2222_,
    new_n2223_, new_n2224_, new_n2225_, new_n2226_, new_n2227_, new_n2229_,
    new_n2230_, new_n2231_, new_n2232_, new_n2233_, new_n2234_, new_n2235_,
    new_n2236_, new_n2237_, new_n2239_, new_n2240_, new_n2241_, new_n2242_,
    new_n2243_, new_n2244_, new_n2245_, new_n2246_, new_n2247_, new_n2248_,
    new_n2250_, new_n2251_, new_n2252_, new_n2253_, new_n2254_, new_n2255_,
    new_n2256_, new_n2257_, new_n2258_, new_n2259_, new_n2261_, new_n2262_,
    new_n2263_, new_n2264_, new_n2265_, new_n2266_, new_n2267_, new_n2268_,
    new_n2269_, new_n2270_, new_n2272_, new_n2273_, new_n2274_, new_n2275_,
    new_n2276_, new_n2277_, new_n2278_, new_n2279_, new_n2280_, new_n2281_,
    new_n2283_, new_n2284_, new_n2285_, new_n2286_, new_n2287_, new_n2288_,
    new_n2289_, new_n2290_, new_n2291_, new_n2292_, new_n2294_, new_n2295_,
    new_n2296_, new_n2297_, new_n2298_, new_n2299_, new_n2300_, new_n2301_,
    new_n2302_, new_n2303_, new_n2305_, new_n2306_, new_n2307_, new_n2308_,
    new_n2309_, new_n2310_, new_n2311_, new_n2312_, new_n2313_, new_n2314_,
    new_n2316_, new_n2317_, new_n2318_, new_n2319_, new_n2320_, new_n2321_,
    new_n2322_, new_n2323_, new_n2324_, new_n2325_, new_n2327_, new_n2328_,
    new_n2329_, new_n2330_, new_n2331_, new_n2332_, new_n2333_, new_n2334_,
    new_n2335_, new_n2336_, new_n2338_, new_n2339_, new_n2340_, new_n2341_,
    new_n2342_, new_n2343_, new_n2344_, new_n2345_, new_n2346_, new_n2347_,
    new_n2349_, new_n2350_, new_n2351_, new_n2352_, new_n2353_, new_n2354_,
    new_n2355_, new_n2356_, new_n2357_, new_n2358_, new_n2360_, new_n2361_,
    new_n2362_, new_n2363_, new_n2364_, new_n2365_, new_n2366_, new_n2367_,
    new_n2368_, new_n2369_, new_n2371_, new_n2372_, new_n2373_, new_n2374_,
    new_n2375_, new_n2376_, new_n2377_, new_n2378_, new_n2379_, new_n2380_,
    new_n2382_, new_n2383_, new_n2384_, new_n2385_, new_n2386_, new_n2387_,
    new_n2388_, new_n2389_, new_n2390_, new_n2391_, new_n2393_, new_n2394_,
    new_n2395_, new_n2396_, new_n2397_, new_n2398_, new_n2399_, new_n2400_,
    new_n2401_, new_n2402_, new_n2404_, new_n2405_, new_n2406_, new_n2407_,
    new_n2408_, new_n2409_, new_n2410_, new_n2411_, new_n2412_, new_n2413_,
    new_n2415_, new_n2416_, new_n2417_, new_n2418_, new_n2419_, new_n2420_,
    new_n2421_, new_n2422_, new_n2423_, new_n2424_, new_n2426_, new_n2427_,
    new_n2428_, new_n2429_, new_n2430_, new_n2431_, new_n2432_, new_n2433_,
    new_n2434_, new_n2435_, new_n2437_, new_n2438_, new_n2439_, new_n2440_,
    new_n2441_, new_n2442_, new_n2443_, new_n2444_, new_n2445_, new_n2446_,
    new_n2448_, new_n2449_, new_n2450_, new_n2451_, new_n2452_, new_n2453_,
    new_n2454_, new_n2455_, new_n2456_, new_n2457_, new_n2459_, new_n2460_,
    new_n2461_, new_n2462_, new_n2463_, new_n2464_, new_n2465_, new_n2466_,
    new_n2467_, new_n2468_, new_n2470_, new_n2471_, new_n2472_, new_n2473_,
    new_n2474_, new_n2475_, new_n2476_, new_n2477_, new_n2478_, new_n2479_,
    new_n2481_, new_n2482_, new_n2483_, new_n2484_, new_n2485_, new_n2486_,
    new_n2487_, new_n2488_, new_n2489_, new_n2490_, new_n2492_, new_n2493_,
    new_n2494_, new_n2495_, new_n2496_, new_n2497_, new_n2498_, new_n2499_,
    new_n2500_, new_n2501_, new_n2503_, new_n2504_, new_n2505_, new_n2506_,
    new_n2507_, new_n2508_, new_n2509_, new_n2510_, new_n2511_, new_n2512_,
    new_n2514_, new_n2515_, new_n2516_, new_n2517_, new_n2518_, new_n2519_,
    new_n2520_, new_n2521_, new_n2522_, new_n2523_, new_n2525_, new_n2526_,
    new_n2527_, new_n2528_, new_n2529_, new_n2530_, new_n2531_, new_n2532_,
    new_n2533_, new_n2534_, new_n2536_, new_n2537_, new_n2538_, new_n2539_,
    new_n2540_, new_n2541_, new_n2542_, new_n2543_, new_n2544_, new_n2545_,
    new_n2547_, new_n2548_, new_n2549_, new_n2550_, new_n2551_, new_n2552_,
    new_n2553_, new_n2554_, new_n2555_, new_n2556_, new_n2558_, new_n2559_,
    new_n2560_, new_n2561_, new_n2562_, new_n2563_, new_n2564_, new_n2565_,
    new_n2566_, new_n2567_, new_n2569_, new_n2570_, new_n2571_, new_n2572_,
    new_n2573_, new_n2574_, new_n2575_, new_n2576_, new_n2577_, new_n2578_,
    new_n2580_, new_n2581_, new_n2582_, new_n2583_, new_n2584_, new_n2585_,
    new_n2586_, new_n2587_, new_n2588_, new_n2589_, new_n2591_, new_n2592_,
    new_n2593_, new_n2594_, new_n2595_, new_n2596_, new_n2597_, new_n2598_,
    new_n2599_, new_n2600_, new_n2602_, new_n2603_, new_n2604_, new_n2605_,
    new_n2606_, new_n2607_, new_n2608_, new_n2609_, new_n2610_, new_n2611_,
    new_n2613_, new_n2614_, new_n2615_, new_n2616_, new_n2617_, new_n2618_,
    new_n2619_, new_n2620_, new_n2621_, new_n2622_, new_n2624_, new_n2625_,
    new_n2626_, new_n2627_, new_n2628_, new_n2629_, new_n2630_, new_n2631_,
    new_n2632_, new_n2633_, new_n2635_, new_n2636_, new_n2637_, new_n2638_,
    new_n2639_, new_n2640_, new_n2641_, new_n2642_, new_n2643_, new_n2644_,
    new_n2646_, new_n2647_, new_n2648_, new_n2649_, new_n2650_, new_n2651_,
    new_n2652_, new_n2653_, new_n2654_, new_n2655_, new_n2657_, new_n2658_,
    new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2663_, new_n2664_,
    new_n2665_, new_n2666_, new_n2668_, new_n2669_, new_n2670_, new_n2671_,
    new_n2672_, new_n2673_, new_n2674_, new_n2675_, new_n2676_, new_n2677_,
    new_n2679_, new_n2680_, new_n2681_, new_n2682_, new_n2683_, new_n2684_,
    new_n2685_, new_n2686_, new_n2687_, new_n2688_, new_n2690_, new_n2691_,
    new_n2692_, new_n2693_, new_n2694_, new_n2695_, new_n2696_, new_n2697_,
    new_n2698_, new_n2699_, new_n2701_, new_n2702_, new_n2703_, new_n2704_,
    new_n2705_, new_n2706_, new_n2707_, new_n2708_, new_n2709_, new_n2710_,
    new_n2712_, new_n2713_, new_n2714_, new_n2715_, new_n2716_, new_n2717_,
    new_n2718_, new_n2719_, new_n2720_, new_n2721_, new_n2723_, new_n2724_,
    new_n2725_, new_n2726_, new_n2727_, new_n2728_, new_n2729_, new_n2730_,
    new_n2731_, new_n2732_, new_n2734_, new_n2735_, new_n2736_, new_n2737_,
    new_n2738_, new_n2739_, new_n2740_, new_n2741_, new_n2742_, new_n2743_,
    new_n2745_, new_n2746_, new_n2747_, new_n2748_, new_n2749_, new_n2750_,
    new_n2751_, new_n2752_, new_n2753_, new_n2754_, new_n2756_, new_n2757_,
    new_n2758_, new_n2759_, new_n2760_, new_n2761_, new_n2762_, new_n2763_,
    new_n2764_, new_n2765_, new_n2767_, new_n2768_, new_n2769_, new_n2770_,
    new_n2771_, new_n2772_, new_n2773_, new_n2774_, new_n2775_, new_n2776_,
    new_n2778_, new_n2779_, new_n2780_, new_n2781_, new_n2782_, new_n2783_,
    new_n2784_, new_n2785_, new_n2786_, new_n2787_, new_n2789_, new_n2790_,
    new_n2791_, new_n2792_, new_n2793_, new_n2794_, new_n2795_, new_n2796_,
    new_n2797_, new_n2798_, new_n2800_, new_n2801_, new_n2802_, new_n2803_,
    new_n2804_, new_n2805_, new_n2806_, new_n2807_, new_n2808_, new_n2809_,
    new_n2811_, new_n2812_, new_n2813_, new_n2814_, new_n2815_, new_n2816_,
    new_n2817_, new_n2818_, new_n2819_, new_n2820_, new_n2822_, new_n2823_,
    new_n2824_, new_n2825_, new_n2826_, new_n2827_, new_n2828_, new_n2829_,
    new_n2830_, new_n2831_, new_n2833_, new_n2834_, new_n2835_, new_n2836_,
    new_n2837_, new_n2838_, new_n2839_, new_n2840_, new_n2841_, new_n2842_,
    new_n2844_, new_n2845_, new_n2846_, new_n2847_, new_n2848_, new_n2849_,
    new_n2850_, new_n2851_, new_n2852_, new_n2853_, new_n2855_, new_n2856_,
    new_n2857_, new_n2858_, new_n2859_, new_n2860_, new_n2861_, new_n2862_,
    new_n2863_, new_n2864_, new_n2866_, new_n2867_, new_n2868_, new_n2869_,
    new_n2870_, new_n2871_, new_n2872_, new_n2873_, new_n2874_, new_n2875_,
    new_n2877_, new_n2878_, new_n2879_, new_n2880_, new_n2881_, new_n2882_,
    new_n2883_, new_n2884_, new_n2885_, new_n2886_, new_n2888_, new_n2889_,
    new_n2890_, new_n2891_, new_n2892_, new_n2893_, new_n2894_, new_n2895_,
    new_n2896_, new_n2897_, new_n2899_, new_n2900_, new_n2901_, new_n2902_,
    new_n2903_, new_n2904_, new_n2905_, new_n2906_, new_n2907_, new_n2908_,
    new_n2910_, new_n2911_, new_n2912_, new_n2913_, new_n2914_, new_n2915_,
    new_n2916_, new_n2917_, new_n2918_, new_n2919_, new_n2921_, new_n2922_,
    new_n2923_, new_n2924_, new_n2925_, new_n2926_, new_n2927_, new_n2928_,
    new_n2929_, new_n2930_, new_n2932_, new_n2933_, new_n2934_, new_n2935_,
    new_n2936_, new_n2937_, new_n2938_, new_n2939_, new_n2940_, new_n2941_,
    new_n2943_, new_n2944_, new_n2945_, new_n2946_, new_n2947_, new_n2948_,
    new_n2949_, new_n2950_, new_n2951_, new_n2952_, new_n2954_, new_n2955_,
    new_n2956_, new_n2957_, new_n2958_, new_n2959_, new_n2960_, new_n2961_,
    new_n2962_, new_n2963_, new_n2965_, new_n2966_, new_n2967_, new_n2968_,
    new_n2969_, new_n2970_, new_n2971_, new_n2972_, new_n2973_, new_n2974_,
    new_n2976_, new_n2977_, new_n2978_, new_n2979_, new_n2980_, new_n2981_,
    new_n2982_, new_n2983_, new_n2984_, new_n2985_, new_n2987_, new_n2988_,
    new_n2989_, new_n2990_, new_n2991_, new_n2992_, new_n2993_, new_n2994_,
    new_n2995_, new_n2996_, new_n2998_, new_n2999_, new_n3000_, new_n3001_,
    new_n3002_, new_n3003_, new_n3004_, new_n3005_, new_n3006_, new_n3007_,
    new_n3009_, new_n3010_, new_n3011_, new_n3012_, new_n3013_, new_n3014_,
    new_n3015_, new_n3016_, new_n3017_, new_n3018_, new_n3020_, new_n3021_,
    new_n3022_, new_n3023_, new_n3024_, new_n3025_, new_n3026_, new_n3027_,
    new_n3028_, new_n3029_, new_n3031_, new_n3032_, new_n3033_, new_n3034_,
    new_n3035_, new_n3036_, new_n3037_, new_n3038_, new_n3039_, new_n3040_,
    new_n3042_, new_n3043_, new_n3044_, new_n3045_, new_n3046_, new_n3047_,
    new_n3048_, new_n3049_, new_n3050_, new_n3051_, new_n3053_, new_n3054_,
    new_n3055_, new_n3056_, new_n3057_, new_n3058_, new_n3059_, new_n3060_,
    new_n3061_, new_n3062_, new_n3064_, new_n3065_, new_n3066_, new_n3067_,
    new_n3068_, new_n3069_, new_n3070_, new_n3071_, new_n3072_, new_n3073_,
    new_n3075_, new_n3076_, new_n3077_, new_n3078_, new_n3079_, new_n3080_,
    new_n3081_, new_n3082_, new_n3083_, new_n3084_, new_n3086_, new_n3087_,
    new_n3088_, new_n3089_, new_n3090_, new_n3091_, new_n3092_, new_n3093_,
    new_n3094_, new_n3095_, new_n3097_, new_n3098_, new_n3099_, new_n3100_,
    new_n3101_, new_n3102_, new_n3103_, new_n3104_, new_n3105_, new_n3106_,
    new_n3108_, new_n3109_, new_n3110_, new_n3111_, new_n3112_, new_n3113_,
    new_n3114_, new_n3115_, new_n3116_, new_n3117_, new_n3119_, new_n3120_,
    new_n3121_, new_n3122_, new_n3123_, new_n3124_, new_n3125_, new_n3126_,
    new_n3127_, new_n3128_, new_n3130_, new_n3131_, new_n3132_, new_n3133_,
    new_n3134_, new_n3135_, new_n3136_, new_n3137_, new_n3138_, new_n3139_,
    new_n3141_, new_n3142_, new_n3143_, new_n3144_, new_n3145_, new_n3146_,
    new_n3147_, new_n3148_, new_n3149_, new_n3150_, new_n3152_, new_n3153_,
    new_n3154_, new_n3155_, new_n3156_, new_n3157_, new_n3158_, new_n3159_,
    new_n3160_, new_n3161_, new_n3163_, new_n3164_, new_n3165_, new_n3166_,
    new_n3167_, new_n3168_, new_n3169_, new_n3170_, new_n3171_, new_n3172_,
    new_n3174_, new_n3175_, new_n3176_, new_n3177_, new_n3178_, new_n3179_,
    new_n3180_, new_n3181_, new_n3182_, new_n3183_, new_n3185_, new_n3186_,
    new_n3187_, new_n3188_, new_n3189_, new_n3190_, new_n3191_, new_n3192_,
    new_n3193_, new_n3194_, new_n3196_, new_n3197_, new_n3198_, new_n3199_,
    new_n3200_, new_n3201_, new_n3202_, new_n3203_, new_n3204_, new_n3205_,
    new_n3207_, new_n3208_, new_n3209_, new_n3210_, new_n3211_, new_n3212_,
    new_n3213_, new_n3214_, new_n3215_, new_n3216_, new_n3218_, new_n3219_,
    new_n3220_, new_n3221_, new_n3222_, new_n3223_, new_n3224_, new_n3225_,
    new_n3226_, new_n3227_, new_n3229_, new_n3230_, new_n3231_, new_n3232_,
    new_n3233_, new_n3234_, new_n3235_, new_n3236_, new_n3237_, new_n3238_,
    new_n3240_, new_n3241_, new_n3242_, new_n3243_, new_n3244_, new_n3245_,
    new_n3246_, new_n3247_, new_n3248_, new_n3249_, new_n3251_, new_n3252_,
    new_n3253_, new_n3254_, new_n3255_, new_n3256_, new_n3257_, new_n3258_,
    new_n3259_, new_n3260_, new_n3262_, new_n3263_, new_n3264_, new_n3265_,
    new_n3266_, new_n3267_, new_n3268_, new_n3269_, new_n3270_, new_n3271_,
    new_n3273_, new_n3274_, new_n3275_, new_n3276_, new_n3277_, new_n3278_,
    new_n3279_, new_n3280_, new_n3281_, new_n3282_, new_n3284_, new_n3285_,
    new_n3286_, new_n3287_, new_n3288_, new_n3289_, new_n3290_, new_n3291_,
    new_n3292_, new_n3293_, new_n3295_, new_n3296_, new_n3297_, new_n3298_,
    new_n3299_, new_n3300_, new_n3301_, new_n3302_, new_n3303_, new_n3304_,
    new_n3306_, new_n3307_, new_n3308_, new_n3309_, new_n3310_, new_n3311_,
    new_n3312_, new_n3313_, new_n3314_, new_n3315_, new_n3317_, new_n3318_,
    new_n3319_, new_n3320_, new_n3321_, new_n3322_, new_n3323_, new_n3324_,
    new_n3325_, new_n3326_, new_n3328_, new_n3329_, new_n3330_, new_n3331_,
    new_n3332_, new_n3333_, new_n3334_, new_n3335_, new_n3336_, new_n3337_,
    new_n3339_, new_n3340_, new_n3341_, new_n3342_, new_n3343_, new_n3344_,
    new_n3345_, new_n3346_, new_n3347_, new_n3348_, new_n3350_, new_n3351_,
    new_n3352_, new_n3353_, new_n3354_, new_n3355_, new_n3356_, new_n3357_,
    new_n3358_, new_n3359_, new_n3361_, new_n3362_, new_n3363_, new_n3364_,
    new_n3365_, new_n3366_, new_n3367_, new_n3368_, new_n3369_, new_n3370_,
    new_n3372_, new_n3373_, new_n3374_, new_n3375_, new_n3376_, new_n3377_,
    new_n3378_, new_n3379_, new_n3380_, new_n3381_, new_n3383_, new_n3384_,
    new_n3385_, new_n3386_, new_n3387_, new_n3388_, new_n3389_, new_n3390_,
    new_n3391_, new_n3392_, new_n3394_, new_n3395_, new_n3396_, new_n3397_,
    new_n3398_, new_n3399_, new_n3400_, new_n3401_, new_n3402_, new_n3403_,
    new_n3405_, new_n3406_, new_n3407_, new_n3408_, new_n3409_, new_n3410_,
    new_n3411_, new_n3412_, new_n3413_, new_n3414_, new_n3416_, new_n3417_,
    new_n3418_, new_n3419_, new_n3420_, new_n3421_, new_n3422_, new_n3423_,
    new_n3424_, new_n3425_, new_n3427_, new_n3428_, new_n3429_, new_n3430_,
    new_n3431_, new_n3432_, new_n3433_, new_n3434_, new_n3435_, new_n3436_,
    new_n3438_, new_n3439_, new_n3440_, new_n3441_, new_n3442_, new_n3443_,
    new_n3444_, new_n3445_, new_n3446_, new_n3447_, new_n3449_, new_n3450_,
    new_n3451_, new_n3452_, new_n3453_, new_n3454_, new_n3455_, new_n3456_,
    new_n3457_, new_n3458_, new_n3460_, new_n3461_, new_n3462_, new_n3463_,
    new_n3464_, new_n3465_, new_n3466_, new_n3467_, new_n3468_, new_n3469_,
    new_n3471_, new_n3472_, new_n3473_, new_n3474_, new_n3475_, new_n3476_,
    new_n3477_, new_n3478_, new_n3479_, new_n3480_, new_n3482_, new_n3483_,
    new_n3484_, new_n3485_, new_n3486_, new_n3487_, new_n3488_, new_n3489_,
    new_n3490_, new_n3491_, new_n3493_, new_n3494_, new_n3495_, new_n3496_,
    new_n3497_, new_n3498_, new_n3499_, new_n3500_, new_n3501_, new_n3502_,
    new_n3504_, new_n3505_, new_n3506_, new_n3507_, new_n3508_, new_n3509_,
    new_n3510_, new_n3511_, new_n3512_, new_n3513_, new_n3515_, new_n3516_,
    new_n3517_, new_n3518_, new_n3519_, new_n3520_, new_n3521_, new_n3522_,
    new_n3523_, new_n3524_, new_n3526_, new_n3527_, new_n3528_, new_n3529_,
    new_n3530_, new_n3531_, new_n3532_, new_n3533_, new_n3534_, new_n3535_,
    new_n3537_, new_n3538_, new_n3539_, new_n3540_, new_n3541_, new_n3542_,
    new_n3543_, new_n3544_, new_n3545_, new_n3546_, new_n3548_, new_n3549_,
    new_n3550_, new_n3551_, new_n3552_, new_n3553_, new_n3554_, new_n3555_,
    new_n3556_, new_n3557_, new_n3559_, new_n3560_, new_n3561_, new_n3562_,
    new_n3563_, new_n3564_, new_n3565_, new_n3566_, new_n3567_, new_n3568_,
    new_n3570_, new_n3571_, new_n3572_, new_n3573_, new_n3574_, new_n3575_,
    new_n3576_, new_n3577_, new_n3578_, new_n3579_, new_n3581_, new_n3582_,
    new_n3583_, new_n3584_, new_n3585_, new_n3586_, new_n3587_, new_n3588_,
    new_n3589_, new_n3590_, new_n3592_, new_n3593_, new_n3594_, new_n3595_,
    new_n3596_, new_n3597_, new_n3598_, new_n3599_, new_n3600_, new_n3601_,
    new_n3603_, new_n3604_, new_n3605_, new_n3606_, new_n3607_, new_n3608_,
    new_n3609_, new_n3610_, new_n3611_, new_n3612_, new_n3614_, new_n3615_,
    new_n3616_, new_n3617_, new_n3618_, new_n3619_, new_n3620_, new_n3621_,
    new_n3622_, new_n3623_, n854, n859, n864, n869, n874, n879, n884, n889,
    n894, n899, n904, n909, n914, n919, n924, n929, n934, n939, n944, n949,
    n954, n959, n964, n969, n974, n979, n984, n989, n994, n999, n1004,
    n1009, n1014, n1019, n1024, n1029, n1034, n1039, n1044, n1049, n1054,
    n1059, n1064, n1069, n1074, n1079, n1084, n1089, n1094, n1099, n1104,
    n1109, n1114, n1119, n1124, n1129, n1134, n1139, n1144, n1149, n1154,
    n1159, n1164, n1169, n1174, n1179, n1184, n1189, n1194, n1199, n1204,
    n1209, n1214, n1219, n1224, n1229, n1234, n1239, n1244, n1249, n1254,
    n1259, n1264, n1269, n1274, n1279, n1284, n1289, n1294, n1299, n1304,
    n1309, n1314, n1319, n1324, n1329, n1334, n1339, n1344, n1349, n1354,
    n1359, n1364, n1369, n1374, n1379, n1384, n1389, n1394, n1399, n1404,
    n1409, n1414, n1419, n1424, n1429, n1434, n1439, n1444, n1449, n1454,
    n1459, n1464, n1469, n1474, n1479, n1484, n1489, n1494, n1499, n1504,
    n1509, n1514, n1519, n1524, n1529, n1534, n1539, n1544, n1549, n1554,
    n1559, n1564, n1569, n1574, n1579, n1584, n1589, n1594, n1599, n1604,
    n1609, n1614, n1619, n1624, n1629, n1634, n1639, n1644, n1649, n1654,
    n1659, n1664, n1669, n1674, n1679, n1684, n1689, n1694, n1699, n1704,
    n1709, n1714, n1719, n1724, n1729, n1734, n1739, n1744, n1749, n1754,
    n1759, n1764, n1769, n1774, n1779, n1784, n1789, n1794, n1799, n1804,
    n1809, n1814, n1819, n1824, n1829, n1834, n1839, n1844, n1849, n1854,
    n1859, n1864, n1869, n1874, n1879, n1884, n1889, n1894, n1899, n1904,
    n1909, n1914, n1919, n1924, n1929, n1934, n1939, n1944, n1949, n1954,
    n1959, n1964, n1969;
  assign new_n1099_1_ = ~pstart_0_ & ~pencrypt_0_;
  assign new_n1100_ = pcount_3_ & ~pcount_0_;
  assign new_n1101_ = pcount_2_ & pcount_1_;
  assign new_n1102_ = new_n1100_ & new_n1101_;
  assign new_n1103_ = pcount_1_ & pcount_0_;
  assign new_n1104_1_ = ~pcount_3_ & new_n1103_;
  assign new_n1105_ = pcount_2_ & new_n1104_1_;
  assign new_n1106_ = ~pcount_2_ & ~pcount_0_;
  assign new_n1107_ = ~pcount_1_ & new_n1106_;
  assign new_n1108_ = ~pcount_3_ & new_n1107_;
  assign new_n1109_1_ = ~new_n1102_ & ~new_n1105_;
  assign new_n1110_ = ~new_n1108_ & new_n1109_1_;
  assign new_n1111_ = ~pcount_0_ & ~new_n1110_;
  assign new_n1112_ = ~pcount_1_ & new_n1111_;
  assign new_n1113_ = new_n1099_1_ & new_n1112_;
  assign new_n1114_1_ = ~pstart_0_ & pencrypt_0_;
  assign new_n1115_ = ~pcount_3_ & ~pcount_1_;
  assign new_n1116_ = ~pcount_2_ & new_n1115_;
  assign new_n1117_ = ~new_n1103_ & ~new_n1116_;
  assign new_n1118_ = pcount_2_ & new_n1110_;
  assign new_n1119_1_ = ~new_n1116_ & ~new_n1118_;
  assign new_n1120_ = ~new_n1117_ & ~new_n1119_1_;
  assign new_n1121_ = ~new_n1107_ & ~new_n1120_;
  assign new_n1122_ = new_n1103_ & ~new_n1121_;
  assign new_n1123_ = new_n1114_1_ & new_n1122_;
  assign pdata_ready_0_ = new_n1113_ | new_n1123_;
  assign new_n1125_ = ~pencrypt_0_ & new_n1108_;
  assign new_n1126_ = new_n1105_ & new_n1114_1_;
  assign new_n1127_ = ~pcount_2_ & new_n1114_1_;
  assign new_n1128_ = pcount_2_ & ~pencrypt_0_;
  assign new_n1129_1_ = ~new_n1127_ & ~new_n1128_;
  assign new_n1130_ = ~new_n1103_ & new_n1114_1_;
  assign new_n1131_ = ~pcount_1_ & ~pcount_0_;
  assign new_n1132_ = ~pencrypt_0_ & ~new_n1131_;
  assign new_n1133_ = ~new_n1130_ & ~new_n1132_;
  assign new_n1134_1_ = new_n1129_1_ & new_n1133_;
  assign new_n1135_ = pcount_3_ & ~new_n1134_1_;
  assign new_n1136_ = pstart_0_ & ~pencrypt_0_;
  assign new_n1137_ = ~new_n1125_ & ~new_n1126_;
  assign new_n1138_ = ~new_n1135_ & ~new_n1136_;
  assign pnew_count_3_ = ~new_n1137_ | ~new_n1138_;
  assign new_n1140_ = ~pcount_0_ & ~pstart_0_;
  assign pnew_count_0_ = new_n1136_ | new_n1140_;
  assign new_n1142_ = ~pcount_2_ & ~pstart_0_;
  assign new_n1143_ = pencrypt_0_ & new_n1103_;
  assign new_n1144_1_ = new_n1142_ & new_n1143_;
  assign new_n1145_ = pcount_2_ & ~new_n1133_;
  assign new_n1146_ = ~pencrypt_0_ & new_n1107_;
  assign new_n1147_ = ~new_n1144_1_ & ~new_n1145_;
  assign new_n1148_ = ~new_n1136_ & ~new_n1146_;
  assign pnew_count_2_ = ~new_n1147_ | ~new_n1148_;
  assign new_n1150_ = ~new_n1103_ & ~new_n1131_;
  assign new_n1151_ = new_n1114_1_ & new_n1150_;
  assign new_n1152_ = ~pencrypt_0_ & ~new_n1150_;
  assign new_n1153_ = ~new_n1151_ & ~new_n1152_;
  assign new_n1154_1_ = ~pnew_count_0_ & new_n1153_;
  assign new_n1155_ = ~pstart_0_ & new_n1153_;
  assign pnew_count_1_ = ~new_n1154_1_ & ~new_n1155_;
  assign new_n1157_ = new_n1110_ & new_n1114_1_;
  assign new_n1158_ = n_n94 & new_n1157_;
  assign new_n1159_1_ = pkey_0_ & new_n1136_;
  assign new_n1160_ = ~pencrypt_0_ & new_n1121_;
  assign new_n1161_ = ~pstart_0_ & new_n1160_;
  assign new_n1162_ = n_n97 & new_n1161_;
  assign new_n1163_ = ~pencrypt_0_ & ~new_n1121_;
  assign new_n1164_1_ = ~pstart_0_ & new_n1163_;
  assign new_n1165_ = n_n96 & new_n1164_1_;
  assign new_n1166_ = ~new_n1162_ & ~new_n1165_;
  assign new_n1167_ = ~pstart_0_ & ~new_n1110_;
  assign new_n1168_ = pencrypt_0_ & new_n1167_;
  assign new_n1169_1_ = n_n2384 & new_n1168_;
  assign new_n1170_ = pstart_0_ & pencrypt_0_;
  assign new_n1171_ = pkey_57_ & new_n1170_;
  assign new_n1172_ = ~new_n1169_1_ & ~new_n1171_;
  assign new_n1173_ = ~new_n1158_ & ~new_n1159_1_;
  assign new_n1174_1_ = new_n1166_ & new_n1172_;
  assign n854 = ~new_n1173_ | ~new_n1174_1_;
  assign new_n1176_ = n_n104 & new_n1157_;
  assign new_n1177_ = pkey_219_ & new_n1136_;
  assign new_n1178_ = n_n107 & new_n1161_;
  assign new_n1179_1_ = n_n106 & new_n1164_1_;
  assign new_n1180_ = ~new_n1178_ & ~new_n1179_1_;
  assign new_n1181_ = n_n2396 & new_n1168_;
  assign new_n1182_ = pkey_211_ & new_n1170_;
  assign new_n1183_ = ~new_n1181_ & ~new_n1182_;
  assign new_n1184_1_ = ~new_n1176_ & ~new_n1177_;
  assign new_n1185_ = new_n1180_ & new_n1183_;
  assign n859 = ~new_n1184_1_ | ~new_n1185_;
  assign new_n1187_ = n_n114 & new_n1157_;
  assign new_n1188_ = pkey_213_ & new_n1136_;
  assign new_n1189_1_ = n_n115 & new_n1161_;
  assign new_n1190_ = n_n2412 & new_n1164_1_;
  assign new_n1191_ = ~new_n1189_1_ & ~new_n1190_;
  assign new_n1192_ = n_n2408 & new_n1168_;
  assign new_n1193_ = pkey_205_ & new_n1170_;
  assign new_n1194_1_ = ~new_n1192_ & ~new_n1193_;
  assign new_n1195_ = ~new_n1187_ & ~new_n1188_;
  assign new_n1196_ = new_n1191_ & new_n1194_1_;
  assign n864 = ~new_n1195_ | ~new_n1196_;
  assign new_n1198_ = n_n120 & new_n1157_;
  assign new_n1199_1_ = pkey_238_ & new_n1136_;
  assign new_n1200_ = n_n124 & new_n1161_;
  assign new_n1201_ = n_n123 & new_n1164_1_;
  assign new_n1202_ = ~new_n1200_ & ~new_n1201_;
  assign new_n1203_ = n_n121 & new_n1168_;
  assign new_n1204_1_ = pkey_230_ & new_n1170_;
  assign new_n1205_ = ~new_n1203_ & ~new_n1204_1_;
  assign new_n1206_ = ~new_n1198_ & ~new_n1199_1_;
  assign new_n1207_ = new_n1202_ & new_n1205_;
  assign n869 = ~new_n1206_ | ~new_n1207_;
  assign new_n1209_1_ = n_n130 & new_n1157_;
  assign new_n1210_ = pkey_164_ & new_n1136_;
  assign new_n1211_ = n_n134 & new_n1161_;
  assign new_n1212_ = n_n133 & new_n1164_1_;
  assign new_n1213_ = ~new_n1211_ & ~new_n1212_;
  assign new_n1214_1_ = n_n131 & new_n1168_;
  assign new_n1215_ = pkey_156_ & new_n1170_;
  assign new_n1216_ = ~new_n1214_1_ & ~new_n1215_;
  assign new_n1217_ = ~new_n1209_1_ & ~new_n1210_;
  assign new_n1218_ = new_n1213_ & new_n1216_;
  assign n874 = ~new_n1217_ | ~new_n1218_;
  assign new_n1220_ = n_n140 & new_n1157_;
  assign new_n1221_ = pkey_189_ & new_n1136_;
  assign new_n1222_ = n_n2452 & new_n1161_;
  assign new_n1223_ = n_n142 & new_n1164_1_;
  assign new_n1224_1_ = ~new_n1222_ & ~new_n1223_;
  assign new_n1225_ = n_n2448 & new_n1168_;
  assign new_n1226_ = pkey_181_ & new_n1170_;
  assign new_n1227_ = ~new_n1225_ & ~new_n1226_;
  assign new_n1228_ = ~new_n1220_ & ~new_n1221_;
  assign new_n1229_1_ = new_n1224_1_ & new_n1227_;
  assign n879 = ~new_n1228_ | ~new_n1229_1_;
  assign new_n1231_ = n_n176 & new_n1157_;
  assign new_n1232_ = pkey_28_ & new_n1136_;
  assign new_n1233_ = n_n180 & new_n1161_;
  assign new_n1234_1_ = n_n179 & new_n1164_1_;
  assign new_n1235_ = ~new_n1233_ & ~new_n1234_1_;
  assign new_n1236_ = n_n177 & new_n1168_;
  assign new_n1237_ = pkey_20_ & new_n1170_;
  assign new_n1238_ = ~new_n1236_ & ~new_n1237_;
  assign new_n1239_1_ = ~new_n1231_ & ~new_n1232_;
  assign new_n1240_ = new_n1235_ & new_n1238_;
  assign n884 = ~new_n1239_1_ | ~new_n1240_;
  assign new_n1242_ = n_n186 & new_n1157_;
  assign new_n1243_ = pkey_53_ & new_n1136_;
  assign new_n1244_1_ = n_n189 & new_n1161_;
  assign new_n1245_ = n_n188 & new_n1164_1_;
  assign new_n1246_ = ~new_n1244_1_ & ~new_n1245_;
  assign new_n1247_ = n_n187 & new_n1168_;
  assign new_n1248_ = pkey_45_ & new_n1170_;
  assign new_n1249_1_ = ~new_n1247_ & ~new_n1248_;
  assign new_n1250_ = ~new_n1242_ & ~new_n1243_;
  assign new_n1251_ = new_n1246_ & new_n1249_1_;
  assign n889 = ~new_n1250_ | ~new_n1251_;
  assign new_n1253_ = n_n2384 & new_n1157_;
  assign new_n1254_1_ = pkey_8_ & new_n1136_;
  assign new_n1255_ = n_n98 & new_n1161_;
  assign new_n1256_ = n_n97 & new_n1164_1_;
  assign new_n1257_ = ~new_n1255_ & ~new_n1256_;
  assign new_n1258_ = n_n95 & new_n1168_;
  assign new_n1259_1_ = pkey_0_ & new_n1170_;
  assign new_n1260_ = ~new_n1258_ & ~new_n1259_1_;
  assign new_n1261_ = ~new_n1253_ & ~new_n1254_1_;
  assign new_n1262_ = new_n1257_ & new_n1260_;
  assign n894 = ~new_n1261_ | ~new_n1262_;
  assign new_n1264_1_ = n_n103 & new_n1157_;
  assign new_n1265_ = pkey_211_ & new_n1136_;
  assign new_n1266_ = n_n106 & new_n1161_;
  assign new_n1267_ = n_n105 & new_n1164_1_;
  assign new_n1268_ = ~new_n1266_ & ~new_n1267_;
  assign new_n1269_1_ = n_n104 & new_n1168_;
  assign new_n1270_ = pkey_203_ & new_n1170_;
  assign new_n1271_ = ~new_n1269_1_ & ~new_n1270_;
  assign new_n1272_ = ~new_n1264_1_ & ~new_n1265_;
  assign new_n1273_ = new_n1268_ & new_n1271_;
  assign n899 = ~new_n1272_ | ~new_n1273_;
  assign new_n1275_ = n_n2408 & new_n1157_;
  assign new_n1276_ = pkey_221_ & new_n1136_;
  assign new_n1277_ = n_n116 & new_n1161_;
  assign new_n1278_ = n_n115 & new_n1164_1_;
  assign new_n1279_1_ = ~new_n1277_ & ~new_n1278_;
  assign new_n1280_ = n_n2410 & new_n1168_;
  assign new_n1281_ = pkey_213_ & new_n1170_;
  assign new_n1282_ = ~new_n1280_ & ~new_n1281_;
  assign new_n1283_ = ~new_n1275_ & ~new_n1276_;
  assign new_n1284_1_ = new_n1279_1_ & new_n1282_;
  assign n904 = ~new_n1283_ | ~new_n1284_1_;
  assign new_n1286_ = n_n119 & new_n1157_;
  assign new_n1287_ = pkey_230_ & new_n1136_;
  assign new_n1288_ = n_n123 & new_n1161_;
  assign new_n1289_1_ = n_n122 & new_n1164_1_;
  assign new_n1290_ = ~new_n1288_ & ~new_n1289_1_;
  assign new_n1291_ = n_n120 & new_n1168_;
  assign new_n1292_ = pkey_222_ & new_n1170_;
  assign new_n1293_ = ~new_n1291_ & ~new_n1292_;
  assign new_n1294_1_ = ~new_n1286_ & ~new_n1287_;
  assign new_n1295_ = new_n1290_ & new_n1293_;
  assign n909 = ~new_n1294_1_ | ~new_n1295_;
  assign new_n1297_ = n_n131 & new_n1157_;
  assign new_n1298_ = pkey_172_ & new_n1136_;
  assign new_n1299_1_ = n_n2440 & new_n1161_;
  assign new_n1300_ = n_n134 & new_n1164_1_;
  assign new_n1301_ = ~new_n1299_1_ & ~new_n1300_;
  assign new_n1302_ = n_n132 & new_n1168_;
  assign new_n1303_ = pkey_164_ & new_n1170_;
  assign new_n1304_1_ = ~new_n1302_ & ~new_n1303_;
  assign new_n1305_ = ~new_n1297_ & ~new_n1298_;
  assign new_n1306_ = new_n1301_ & new_n1304_1_;
  assign n914 = ~new_n1305_ | ~new_n1306_;
  assign new_n1308_ = n_n139 & new_n1157_;
  assign new_n1309_1_ = pkey_181_ & new_n1136_;
  assign new_n1310_ = n_n142 & new_n1161_;
  assign new_n1311_ = n_n141 & new_n1164_1_;
  assign new_n1312_ = ~new_n1310_ & ~new_n1311_;
  assign new_n1313_ = n_n140 & new_n1168_;
  assign new_n1314_1_ = pkey_173_ & new_n1170_;
  assign new_n1315_ = ~new_n1313_ & ~new_n1314_1_;
  assign new_n1316_ = ~new_n1308_ & ~new_n1309_1_;
  assign new_n1317_ = new_n1312_ & new_n1315_;
  assign n919 = ~new_n1316_ | ~new_n1317_;
  assign new_n1319_1_ = n_n177 & new_n1157_;
  assign new_n1320_ = pkey_36_ & new_n1136_;
  assign new_n1321_ = n_n181 & new_n1161_;
  assign new_n1322_ = n_n180 & new_n1164_1_;
  assign new_n1323_ = ~new_n1321_ & ~new_n1322_;
  assign new_n1324_1_ = n_n178 & new_n1168_;
  assign new_n1325_ = pkey_28_ & new_n1170_;
  assign new_n1326_ = ~new_n1324_1_ & ~new_n1325_;
  assign new_n1327_ = ~new_n1319_1_ & ~new_n1320_;
  assign new_n1328_ = new_n1323_ & new_n1326_;
  assign n924 = ~new_n1327_ | ~new_n1328_;
  assign new_n1330_ = n_n185 & new_n1157_;
  assign new_n1331_ = pkey_45_ & new_n1136_;
  assign new_n1332_ = n_n188 & new_n1161_;
  assign new_n1333_ = n_n2513 & new_n1164_1_;
  assign new_n1334_1_ = ~new_n1332_ & ~new_n1333_;
  assign new_n1335_ = n_n186 & new_n1168_;
  assign new_n1336_ = pkey_37_ & new_n1170_;
  assign new_n1337_ = ~new_n1335_ & ~new_n1336_;
  assign new_n1338_ = ~new_n1330_ & ~new_n1331_;
  assign new_n1339_1_ = new_n1334_1_ & new_n1337_;
  assign n929 = ~new_n1338_ | ~new_n1339_1_;
  assign new_n1341_ = n_n95 & new_n1157_;
  assign new_n1342_ = pkey_16_ & new_n1136_;
  assign new_n1343_ = n_n99 & new_n1161_;
  assign new_n1344_1_ = n_n98 & new_n1164_1_;
  assign new_n1345_ = ~new_n1343_ & ~new_n1344_1_;
  assign new_n1346_ = n_n96 & new_n1168_;
  assign new_n1347_ = pkey_8_ & new_n1170_;
  assign new_n1348_ = ~new_n1346_ & ~new_n1347_;
  assign new_n1349_1_ = ~new_n1341_ & ~new_n1342_;
  assign new_n1350_ = new_n1345_ & new_n1348_;
  assign n934 = ~new_n1349_1_ | ~new_n1350_;
  assign new_n1352_ = n_n105 & new_n1157_;
  assign new_n1353_ = pkey_204_ & new_n1136_;
  assign new_n1354_1_ = n_n109 & new_n1161_;
  assign new_n1355_ = n_n108 & new_n1164_1_;
  assign new_n1356_ = ~new_n1354_1_ & ~new_n1355_;
  assign new_n1357_ = n_n106 & new_n1168_;
  assign new_n1358_ = pkey_196_ & new_n1170_;
  assign new_n1359_1_ = ~new_n1357_ & ~new_n1358_;
  assign new_n1360_ = ~new_n1352_ & ~new_n1353_;
  assign new_n1361_ = new_n1356_ & new_n1359_1_;
  assign n939 = ~new_n1360_ | ~new_n1361_;
  assign new_n1363_ = n_n112 & new_n1157_;
  assign new_n1364_1_ = pkey_197_ & new_n1136_;
  assign new_n1365_ = n_n2410 & new_n1161_;
  assign new_n1366_ = n_n2408 & new_n1164_1_;
  assign new_n1367_ = ~new_n1365_ & ~new_n1366_;
  assign new_n1368_ = n_n113 & new_n1168_;
  assign new_n1369_1_ = pkey_252_ & new_n1170_;
  assign new_n1370_ = ~new_n1368_ & ~new_n1369_1_;
  assign new_n1371_ = ~new_n1363_ & ~new_n1364_1_;
  assign new_n1372_ = new_n1367_ & new_n1370_;
  assign n944 = ~new_n1371_ | ~new_n1372_;
  assign new_n1374_1_ = n_n2420 & new_n1157_;
  assign new_n1375_ = pkey_222_ & new_n1136_;
  assign new_n1376_ = n_n122 & new_n1161_;
  assign new_n1377_ = n_n121 & new_n1164_1_;
  assign new_n1378_ = ~new_n1376_ & ~new_n1377_;
  assign new_n1379_1_ = n_n119 & new_n1168_;
  assign new_n1380_ = pkey_214_ & new_n1170_;
  assign new_n1381_ = ~new_n1379_1_ & ~new_n1380_;
  assign new_n1382_ = ~new_n1374_1_ & ~new_n1375_;
  assign new_n1383_ = new_n1378_ & new_n1381_;
  assign n949 = ~new_n1382_ | ~new_n1383_;
  assign new_n1385_ = n_n147 & new_n1157_;
  assign new_n1386_ = pkey_67_ & new_n1136_;
  assign new_n1387_ = n_n2462 & new_n1161_;
  assign new_n1388_ = n_n150 & new_n1164_1_;
  assign new_n1389_1_ = ~new_n1387_ & ~new_n1388_;
  assign new_n1390_ = n_n148 & new_n1168_;
  assign new_n1391_ = pkey_190_ & new_n1170_;
  assign new_n1392_ = ~new_n1390_ & ~new_n1391_;
  assign new_n1393_ = ~new_n1385_ & ~new_n1386_;
  assign new_n1394_1_ = new_n1389_1_ & new_n1392_;
  assign n954 = ~new_n1393_ | ~new_n1394_1_;
  assign new_n1396_ = n_n157 & new_n1157_;
  assign new_n1397_ = pkey_124_ & new_n1136_;
  assign new_n1398_ = n_n2474 & new_n1161_;
  assign new_n1399_1_ = n_n160 & new_n1164_1_;
  assign new_n1400_ = ~new_n1398_ & ~new_n1399_1_;
  assign new_n1401_ = n_n158 & new_n1168_;
  assign new_n1402_ = pkey_116_ & new_n1170_;
  assign new_n1403_ = ~new_n1401_ & ~new_n1402_;
  assign new_n1404_1_ = ~new_n1396_ & ~new_n1397_;
  assign new_n1405_ = new_n1400_ & new_n1403_;
  assign n959 = ~new_n1404_1_ | ~new_n1405_;
  assign new_n1407_ = n_n178 & new_n1157_;
  assign new_n1408_ = pkey_44_ & new_n1136_;
  assign new_n1409_1_ = n_n182 & new_n1161_;
  assign new_n1410_ = n_n181 & new_n1164_1_;
  assign new_n1411_ = ~new_n1409_1_ & ~new_n1410_;
  assign new_n1412_ = n_n179 & new_n1168_;
  assign new_n1413_ = pkey_36_ & new_n1170_;
  assign new_n1414_1_ = ~new_n1412_ & ~new_n1413_;
  assign new_n1415_ = ~new_n1407_ & ~new_n1408_;
  assign new_n1416_ = new_n1411_ & new_n1414_1_;
  assign n964 = ~new_n1415_ | ~new_n1416_;
  assign new_n1418_ = n_n2513 & new_n1157_;
  assign new_n1419_1_ = pkey_6_ & new_n1136_;
  assign new_n1420_ = n_n190 & new_n1161_;
  assign new_n1421_ = n_n2517 & new_n1164_1_;
  assign new_n1422_ = ~new_n1420_ & ~new_n1421_;
  assign new_n1423_ = n_n188 & new_n1168_;
  assign new_n1424_1_ = pkey_61_ & new_n1170_;
  assign new_n1425_ = ~new_n1423_ & ~new_n1424_1_;
  assign new_n1426_ = ~new_n1418_ & ~new_n1419_1_;
  assign new_n1427_ = new_n1422_ & new_n1425_;
  assign n969 = ~new_n1426_ | ~new_n1427_;
  assign new_n1429_1_ = n_n193 & new_n1157_;
  assign new_n1430_ = pkey_62_ & new_n1136_;
  assign new_n1431_ = n_n104 & new_n1161_;
  assign new_n1432_ = n_n103 & new_n1164_1_;
  assign new_n1433_ = ~new_n1431_ & ~new_n1432_;
  assign new_n1434_1_ = n_n194 & new_n1168_;
  assign new_n1435_ = pkey_54_ & new_n1170_;
  assign new_n1436_ = ~new_n1434_1_ & ~new_n1435_;
  assign new_n1437_ = ~new_n1429_1_ & ~new_n1430_;
  assign new_n1438_ = new_n1433_ & new_n1436_;
  assign n974 = ~new_n1437_ | ~new_n1438_;
  assign new_n1440_ = n_n96 & new_n1157_;
  assign new_n1441_ = pkey_24_ & new_n1136_;
  assign new_n1442_ = n_n100 & new_n1161_;
  assign new_n1443_ = n_n99 & new_n1164_1_;
  assign new_n1444_1_ = ~new_n1442_ & ~new_n1443_;
  assign new_n1445_ = n_n97 & new_n1168_;
  assign new_n1446_ = pkey_16_ & new_n1170_;
  assign new_n1447_ = ~new_n1445_ & ~new_n1446_;
  assign new_n1448_ = ~new_n1440_ & ~new_n1441_;
  assign new_n1449_1_ = new_n1444_1_ & new_n1447_;
  assign n979 = ~new_n1448_ | ~new_n1449_1_;
  assign new_n1451_ = n_n2396 & new_n1157_;
  assign new_n1452_ = pkey_196_ & new_n1136_;
  assign new_n1453_ = n_n108 & new_n1161_;
  assign new_n1454_1_ = n_n107 & new_n1164_1_;
  assign new_n1455_ = ~new_n1453_ & ~new_n1454_1_;
  assign new_n1456_ = n_n105 & new_n1168_;
  assign new_n1457_ = pkey_219_ & new_n1170_;
  assign new_n1458_ = ~new_n1456_ & ~new_n1457_;
  assign new_n1459_1_ = ~new_n1451_ & ~new_n1452_;
  assign new_n1460_ = new_n1455_ & new_n1458_;
  assign n984 = ~new_n1459_1_ | ~new_n1460_;
  assign new_n1462_ = n_n113 & new_n1157_;
  assign new_n1463_ = pkey_205_ & new_n1136_;
  assign new_n1464_1_ = n_n2412 & new_n1161_;
  assign new_n1465_ = n_n2410 & new_n1164_1_;
  assign new_n1466_ = ~new_n1464_1_ & ~new_n1465_;
  assign new_n1467_ = n_n114 & new_n1168_;
  assign new_n1468_ = pkey_197_ & new_n1170_;
  assign new_n1469_1_ = ~new_n1467_ & ~new_n1468_;
  assign new_n1470_ = ~new_n1462_ & ~new_n1463_;
  assign new_n1471_ = new_n1466_ & new_n1469_1_;
  assign n989 = ~new_n1470_ | ~new_n1471_;
  assign new_n1473_ = n_n118 & new_n1157_;
  assign new_n1474_1_ = pkey_214_ & new_n1136_;
  assign new_n1475_ = n_n121 & new_n1161_;
  assign new_n1476_ = n_n120 & new_n1164_1_;
  assign new_n1477_ = ~new_n1475_ & ~new_n1476_;
  assign new_n1478_ = n_n2420 & new_n1168_;
  assign new_n1479_1_ = pkey_206_ & new_n1170_;
  assign new_n1480_ = ~new_n1478_ & ~new_n1479_1_;
  assign new_n1481_ = ~new_n1473_ & ~new_n1474_1_;
  assign new_n1482_ = new_n1477_ & new_n1480_;
  assign n994 = ~new_n1481_ | ~new_n1482_;
  assign new_n1484_1_ = n_n148 & new_n1157_;
  assign new_n1485_ = pkey_75_ & new_n1136_;
  assign new_n1486_ = n_n151 & new_n1161_;
  assign new_n1487_ = n_n2462 & new_n1164_1_;
  assign new_n1488_ = ~new_n1486_ & ~new_n1487_;
  assign new_n1489_1_ = n_n149 & new_n1168_;
  assign new_n1490_ = pkey_67_ & new_n1170_;
  assign new_n1491_ = ~new_n1489_1_ & ~new_n1490_;
  assign new_n1492_ = ~new_n1484_1_ & ~new_n1485_;
  assign new_n1493_ = new_n1488_ & new_n1491_;
  assign n999 = ~new_n1492_ | ~new_n1493_;
  assign new_n1495_ = n_n156 & new_n1157_;
  assign new_n1496_ = pkey_116_ & new_n1136_;
  assign new_n1497_ = n_n160 & new_n1161_;
  assign new_n1498_ = n_n159 & new_n1164_1_;
  assign new_n1499_1_ = ~new_n1497_ & ~new_n1498_;
  assign new_n1500_ = n_n157 & new_n1168_;
  assign new_n1501_ = pkey_44_ & new_n1170_;
  assign new_n1502_ = ~new_n1500_ & ~new_n1501_;
  assign new_n1503_ = ~new_n1495_ & ~new_n1496_;
  assign new_n1504_1_ = new_n1499_1_ & new_n1502_;
  assign n1004 = ~new_n1503_ | ~new_n1504_1_;
  assign new_n1506_ = n_n179 & new_n1157_;
  assign new_n1507_ = pkey_52_ & new_n1136_;
  assign new_n1508_ = n_n183 & new_n1161_;
  assign new_n1509_1_ = n_n182 & new_n1164_1_;
  assign new_n1510_ = ~new_n1508_ & ~new_n1509_1_;
  assign new_n1511_ = n_n180 & new_n1168_;
  assign new_n1512_ = ~new_n1501_ & ~new_n1511_;
  assign new_n1513_ = ~new_n1506_ & ~new_n1507_;
  assign new_n1514_1_ = new_n1510_ & new_n1512_;
  assign n1009 = ~new_n1513_ | ~new_n1514_1_;
  assign new_n1516_ = n_n187 & new_n1157_;
  assign new_n1517_ = pkey_61_ & new_n1136_;
  assign new_n1518_ = n_n2517 & new_n1161_;
  assign new_n1519_1_ = n_n189 & new_n1164_1_;
  assign new_n1520_ = ~new_n1518_ & ~new_n1519_1_;
  assign new_n1521_ = n_n2513 & new_n1168_;
  assign new_n1522_ = pkey_53_ & new_n1170_;
  assign new_n1523_ = ~new_n1521_ & ~new_n1522_;
  assign new_n1524_1_ = ~new_n1516_ & ~new_n1517_;
  assign new_n1525_ = new_n1520_ & new_n1523_;
  assign n1014 = ~new_n1524_1_ | ~new_n1525_;
  assign new_n1527_ = n_n13 & new_n1157_;
  assign new_n1528_ = pkey_234_ & new_n1136_;
  assign new_n1529_1_ = n_n16 & new_n1161_;
  assign new_n1530_ = n_n2277 & new_n1164_1_;
  assign new_n1531_ = ~new_n1529_1_ & ~new_n1530_;
  assign new_n1532_ = n_n14 & new_n1168_;
  assign new_n1533_ = pkey_226_ & new_n1170_;
  assign new_n1534_1_ = ~new_n1532_ & ~new_n1533_;
  assign new_n1535_ = ~new_n1527_ & ~new_n1528_;
  assign new_n1536_ = new_n1531_ & new_n1534_1_;
  assign n1019 = ~new_n1535_ | ~new_n1536_;
  assign new_n1538_ = n_n90 & new_n1157_;
  assign new_n1539_1_ = pkey_33_ & new_n1136_;
  assign new_n1540_ = n_n94 & new_n1161_;
  assign new_n1541_ = n_n93 & new_n1164_1_;
  assign new_n1542_ = ~new_n1540_ & ~new_n1541_;
  assign new_n1543_ = n_n91 & new_n1168_;
  assign new_n1544_1_ = pkey_25_ & new_n1170_;
  assign new_n1545_ = ~new_n1543_ & ~new_n1544_1_;
  assign new_n1546_ = ~new_n1538_ & ~new_n1539_1_;
  assign new_n1547_ = new_n1542_ & new_n1545_;
  assign n1024 = ~new_n1546_ | ~new_n1547_;
  assign new_n1549_1_ = n_n100 & new_n1157_;
  assign new_n1550_ = pkey_56_ & new_n1136_;
  assign new_n1551_ = n_n9 & new_n1161_;
  assign new_n1552_ = n_n8 & new_n1164_1_;
  assign new_n1553_ = ~new_n1551_ & ~new_n1552_;
  assign new_n1554_1_ = n_n101 & new_n1168_;
  assign new_n1555_ = pkey_48_ & new_n1170_;
  assign new_n1556_ = ~new_n1554_1_ & ~new_n1555_;
  assign new_n1557_ = ~new_n1549_1_ & ~new_n1550_;
  assign new_n1558_ = new_n1553_ & new_n1556_;
  assign n1029 = ~new_n1557_ | ~new_n1558_;
  assign new_n1560_ = n_n110 & new_n1157_;
  assign new_n1561_ = pkey_244_ & new_n1136_;
  assign new_n1562_ = n_n114 & new_n1161_;
  assign new_n1563_ = n_n113 & new_n1164_1_;
  assign new_n1564_1_ = ~new_n1562_ & ~new_n1563_;
  assign new_n1565_ = n_n111 & new_n1168_;
  assign new_n1566_ = pkey_172_ & new_n1170_;
  assign new_n1567_ = ~new_n1565_ & ~new_n1566_;
  assign new_n1568_ = ~new_n1560_ & ~new_n1561_;
  assign new_n1569_1_ = new_n1564_1_ & new_n1567_;
  assign n1034 = ~new_n1568_ | ~new_n1569_1_;
  assign new_n1571_ = n_n117 & new_n1157_;
  assign new_n1572_ = pkey_206_ & new_n1136_;
  assign new_n1573_ = n_n120 & new_n1161_;
  assign new_n1574_1_ = n_n119 & new_n1164_1_;
  assign new_n1575_ = ~new_n1573_ & ~new_n1574_1_;
  assign new_n1576_ = n_n118 & new_n1168_;
  assign new_n1577_ = pkey_198_ & new_n1170_;
  assign new_n1578_ = ~new_n1576_ & ~new_n1577_;
  assign new_n1579_1_ = ~new_n1571_ & ~new_n1572_;
  assign new_n1580_ = new_n1575_ & new_n1578_;
  assign n1039 = ~new_n1579_1_ | ~new_n1580_;
  assign new_n1582_ = n_n2481 & new_n1157_;
  assign new_n1583_ = pkey_70_ & new_n1136_;
  assign new_n1584_1_ = n_n166 & new_n1161_;
  assign new_n1585_ = n_n2485 & new_n1164_1_;
  assign new_n1586_ = ~new_n1584_1_ & ~new_n1585_;
  assign new_n1587_ = n_n164 & new_n1168_;
  assign new_n1588_ = pkey_125_ & new_n1170_;
  assign new_n1589_1_ = ~new_n1587_ & ~new_n1588_;
  assign new_n1590_ = ~new_n1582_ & ~new_n1583_;
  assign new_n1591_ = new_n1586_ & new_n1589_1_;
  assign n1044 = ~new_n1590_ | ~new_n1591_;
  assign new_n1593_ = n_n173 & new_n1157_;
  assign new_n1594_1_ = pkey_27_ & new_n1136_;
  assign new_n1595_ = n_n176 & new_n1161_;
  assign new_n1596_ = n_n175 & new_n1164_1_;
  assign new_n1597_ = ~new_n1595_ & ~new_n1596_;
  assign new_n1598_ = n_n2495 & new_n1168_;
  assign new_n1599_1_ = pkey_19_ & new_n1170_;
  assign new_n1600_ = ~new_n1598_ & ~new_n1599_1_;
  assign new_n1601_ = ~new_n1593_ & ~new_n1594_1_;
  assign new_n1602_ = new_n1597_ & new_n1600_;
  assign n1049 = ~new_n1601_ | ~new_n1602_;
  assign new_n1604_1_ = n_n183 & new_n1157_;
  assign new_n1605_ = pkey_21_ & new_n1136_;
  assign new_n1606_ = n_n186 & new_n1161_;
  assign new_n1607_ = n_n185 & new_n1164_1_;
  assign new_n1608_ = ~new_n1606_ & ~new_n1607_;
  assign new_n1609_1_ = n_n2507 & new_n1168_;
  assign new_n1610_ = pkey_13_ & new_n1170_;
  assign new_n1611_ = ~new_n1609_1_ & ~new_n1610_;
  assign new_n1612_ = ~new_n1604_1_ & ~new_n1605_;
  assign new_n1613_ = new_n1608_ & new_n1611_;
  assign n1054 = ~new_n1612_ | ~new_n1613_;
  assign new_n1615_ = n_n191 & new_n1157_;
  assign new_n1616_ = pkey_46_ & new_n1136_;
  assign new_n1617_ = n_n195 & new_n1161_;
  assign new_n1618_ = n_n194 & new_n1164_1_;
  assign new_n1619_1_ = ~new_n1617_ & ~new_n1618_;
  assign new_n1620_ = n_n192 & new_n1168_;
  assign new_n1621_ = pkey_38_ & new_n1170_;
  assign new_n1622_ = ~new_n1620_ & ~new_n1621_;
  assign new_n1623_ = ~new_n1615_ & ~new_n1616_;
  assign new_n1624_1_ = new_n1619_1_ & new_n1622_;
  assign n1059 = ~new_n1623_ | ~new_n1624_1_;
  assign new_n1626_ = n_n91 & new_n1157_;
  assign new_n1627_ = pkey_41_ & new_n1136_;
  assign new_n1628_ = n_n2384 & new_n1161_;
  assign new_n1629_1_ = n_n94 & new_n1164_1_;
  assign new_n1630_ = ~new_n1628_ & ~new_n1629_1_;
  assign new_n1631_ = n_n92 & new_n1168_;
  assign new_n1632_ = pkey_33_ & new_n1170_;
  assign new_n1633_ = ~new_n1631_ & ~new_n1632_;
  assign new_n1634_1_ = ~new_n1626_ & ~new_n1627_;
  assign new_n1635_ = new_n1630_ & new_n1633_;
  assign n1064 = ~new_n1634_1_ | ~new_n1635_;
  assign new_n1637_ = n_n99 & new_n1157_;
  assign new_n1638_ = pkey_48_ & new_n1136_;
  assign new_n1639_1_ = n_n8 & new_n1161_;
  assign new_n1640_ = n_n102 & new_n1164_1_;
  assign new_n1641_ = ~new_n1639_1_ & ~new_n1640_;
  assign new_n1642_ = n_n100 & new_n1168_;
  assign new_n1643_ = pkey_40_ & new_n1170_;
  assign new_n1644_1_ = ~new_n1642_ & ~new_n1643_;
  assign new_n1645_ = ~new_n1637_ & ~new_n1638_;
  assign new_n1646_ = new_n1641_ & new_n1644_1_;
  assign n1069 = ~new_n1645_ | ~new_n1646_;
  assign new_n1648_ = n_n111 & new_n1157_;
  assign new_n1649_1_ = pkey_252_ & new_n1136_;
  assign new_n1650_ = n_n2408 & new_n1161_;
  assign new_n1651_ = n_n114 & new_n1164_1_;
  assign new_n1652_ = ~new_n1650_ & ~new_n1651_;
  assign new_n1653_ = n_n112 & new_n1168_;
  assign new_n1654_1_ = pkey_244_ & new_n1170_;
  assign new_n1655_ = ~new_n1653_ & ~new_n1654_1_;
  assign new_n1656_ = ~new_n1648_ & ~new_n1649_1_;
  assign new_n1657_ = new_n1652_ & new_n1655_;
  assign n1074 = ~new_n1656_ | ~new_n1657_;
  assign new_n1659_1_ = n_n2416 & new_n1157_;
  assign new_n1660_ = pkey_198_ & new_n1136_;
  assign new_n1661_ = n_n119 & new_n1161_;
  assign new_n1662_ = n_n2420 & new_n1164_1_;
  assign new_n1663_ = ~new_n1661_ & ~new_n1662_;
  assign new_n1664_1_ = n_n117 & new_n1168_;
  assign new_n1665_ = pkey_253_ & new_n1170_;
  assign new_n1666_ = ~new_n1664_1_ & ~new_n1665_;
  assign new_n1667_ = ~new_n1659_1_ & ~new_n1660_;
  assign new_n1668_ = new_n1663_ & new_n1666_;
  assign n1079 = ~new_n1667_ | ~new_n1668_;
  assign new_n1670_ = n_n164 & new_n1157_;
  assign new_n1671_ = pkey_78_ & new_n1136_;
  assign new_n1672_ = n_n167 & new_n1161_;
  assign new_n1673_ = n_n166 & new_n1164_1_;
  assign new_n1674_1_ = ~new_n1672_ & ~new_n1673_;
  assign new_n1675_ = n_n165 & new_n1168_;
  assign new_n1676_ = pkey_70_ & new_n1170_;
  assign new_n1677_ = ~new_n1675_ & ~new_n1676_;
  assign new_n1678_ = ~new_n1670_ & ~new_n1671_;
  assign new_n1679_1_ = new_n1674_1_ & new_n1677_;
  assign n1084 = ~new_n1678_ | ~new_n1679_1_;
  assign new_n1681_ = n_n172 & new_n1157_;
  assign new_n1682_ = pkey_19_ & new_n1136_;
  assign new_n1683_ = n_n175 & new_n1161_;
  assign new_n1684_1_ = n_n174 & new_n1164_1_;
  assign new_n1685_ = ~new_n1683_ & ~new_n1684_1_;
  assign new_n1686_ = n_n173 & new_n1168_;
  assign new_n1687_ = pkey_11_ & new_n1170_;
  assign new_n1688_ = ~new_n1686_ & ~new_n1687_;
  assign new_n1689_1_ = ~new_n1681_ & ~new_n1682_;
  assign new_n1690_ = new_n1685_ & new_n1688_;
  assign n1089 = ~new_n1689_1_ | ~new_n1690_;
  assign new_n1692_ = n_n2495 & new_n1157_;
  assign new_n1693_ = pkey_4_ & new_n1136_;
  assign new_n1694_1_ = n_n177 & new_n1161_;
  assign new_n1695_ = n_n176 & new_n1164_1_;
  assign new_n1696_ = ~new_n1694_1_ & ~new_n1695_;
  assign new_n1697_ = n_n174 & new_n1168_;
  assign new_n1698_ = pkey_27_ & new_n1170_;
  assign new_n1699_1_ = ~new_n1697_ & ~new_n1698_;
  assign new_n1700_ = ~new_n1692_ & ~new_n1693_;
  assign new_n1701_ = new_n1696_ & new_n1699_1_;
  assign n1094 = ~new_n1700_ | ~new_n1701_;
  assign new_n1703_ = n_n192 & new_n1157_;
  assign new_n1704_1_ = pkey_54_ & new_n1136_;
  assign new_n1705_ = n_n103 & new_n1161_;
  assign new_n1706_ = n_n195 & new_n1164_1_;
  assign new_n1707_ = ~new_n1705_ & ~new_n1706_;
  assign new_n1708_ = n_n193 & new_n1168_;
  assign new_n1709_1_ = pkey_46_ & new_n1170_;
  assign new_n1710_ = ~new_n1708_ & ~new_n1709_1_;
  assign new_n1711_ = ~new_n1703_ & ~new_n1704_1_;
  assign new_n1712_ = new_n1707_ & new_n1710_;
  assign n1099 = ~new_n1711_ | ~new_n1712_;
  assign new_n1714_1_ = n_n92 & new_n1157_;
  assign new_n1715_ = pkey_49_ & new_n1136_;
  assign new_n1716_ = n_n95 & new_n1161_;
  assign new_n1717_ = n_n2384 & new_n1164_1_;
  assign new_n1718_ = ~new_n1716_ & ~new_n1717_;
  assign new_n1719_1_ = n_n93 & new_n1168_;
  assign new_n1720_ = pkey_41_ & new_n1170_;
  assign new_n1721_ = ~new_n1719_1_ & ~new_n1720_;
  assign new_n1722_ = ~new_n1714_1_ & ~new_n1715_;
  assign new_n1723_ = new_n1718_ & new_n1721_;
  assign n1104 = ~new_n1722_ | ~new_n1723_;
  assign new_n1725_ = n_n195 & new_n1157_;
  assign new_n1726_ = pkey_203_ & new_n1136_;
  assign new_n1727_ = n_n105 & new_n1161_;
  assign new_n1728_ = n_n2396 & new_n1164_1_;
  assign new_n1729_1_ = ~new_n1727_ & ~new_n1728_;
  assign new_n1730_ = n_n103 & new_n1168_;
  assign new_n1731_ = pkey_195_ & new_n1170_;
  assign new_n1732_ = ~new_n1730_ & ~new_n1731_;
  assign new_n1733_ = ~new_n1725_ & ~new_n1726_;
  assign new_n1734_1_ = new_n1729_1_ & new_n1732_;
  assign n1109 = ~new_n1733_ | ~new_n1734_1_;
  assign new_n1736_ = n_n108 & new_n1157_;
  assign new_n1737_ = pkey_228_ & new_n1136_;
  assign new_n1738_ = n_n112 & new_n1161_;
  assign new_n1739_1_ = n_n111 & new_n1164_1_;
  assign new_n1740_ = ~new_n1738_ & ~new_n1739_1_;
  assign new_n1741_ = n_n109 & new_n1168_;
  assign new_n1742_ = pkey_220_ & new_n1170_;
  assign new_n1743_ = ~new_n1741_ & ~new_n1742_;
  assign new_n1744_1_ = ~new_n1736_ & ~new_n1737_;
  assign new_n1745_ = new_n1740_ & new_n1743_;
  assign n1114 = ~new_n1744_1_ | ~new_n1745_;
  assign new_n1747_ = n_n116 & new_n1157_;
  assign new_n1748_ = pkey_253_ & new_n1136_;
  assign new_n1749_1_ = n_n2420 & new_n1161_;
  assign new_n1750_ = n_n118 & new_n1164_1_;
  assign new_n1751_ = ~new_n1749_1_ & ~new_n1750_;
  assign new_n1752_ = n_n2416 & new_n1168_;
  assign new_n1753_ = pkey_245_ & new_n1170_;
  assign new_n1754_1_ = ~new_n1752_ & ~new_n1753_;
  assign new_n1755_ = ~new_n1747_ & ~new_n1748_;
  assign new_n1756_ = new_n1751_ & new_n1754_1_;
  assign n1119 = ~new_n1755_ | ~new_n1756_;
  assign new_n1758_ = n_n174 & new_n1157_;
  assign new_n1759_1_ = pkey_12_ & new_n1136_;
  assign new_n1760_ = n_n178 & new_n1161_;
  assign new_n1761_ = n_n177 & new_n1164_1_;
  assign new_n1762_ = ~new_n1760_ & ~new_n1761_;
  assign new_n1763_ = n_n175 & new_n1168_;
  assign new_n1764_1_ = pkey_4_ & new_n1170_;
  assign new_n1765_ = ~new_n1763_ & ~new_n1764_1_;
  assign new_n1766_ = ~new_n1758_ & ~new_n1759_1_;
  assign new_n1767_ = new_n1762_ & new_n1765_;
  assign n1124 = ~new_n1766_ | ~new_n1767_;
  assign new_n1769_1_ = n_n184 & new_n1157_;
  assign new_n1770_ = pkey_37_ & new_n1136_;
  assign new_n1771_ = n_n2513 & new_n1161_;
  assign new_n1772_ = n_n187 & new_n1164_1_;
  assign new_n1773_ = ~new_n1771_ & ~new_n1772_;
  assign new_n1774_1_ = n_n185 & new_n1168_;
  assign new_n1775_ = pkey_29_ & new_n1170_;
  assign new_n1776_ = ~new_n1774_1_ & ~new_n1775_;
  assign new_n1777_ = ~new_n1769_1_ & ~new_n1770_;
  assign new_n1778_ = new_n1773_ & new_n1776_;
  assign n1129 = ~new_n1777_ | ~new_n1778_;
  assign new_n1780_ = n_n93 & new_n1157_;
  assign new_n1781_ = pkey_57_ & new_n1136_;
  assign new_n1782_ = n_n96 & new_n1161_;
  assign new_n1783_ = n_n95 & new_n1164_1_;
  assign new_n1784_1_ = ~new_n1782_ & ~new_n1783_;
  assign new_n1785_ = n_n94 & new_n1168_;
  assign new_n1786_ = pkey_49_ & new_n1170_;
  assign new_n1787_ = ~new_n1785_ & ~new_n1786_;
  assign new_n1788_ = ~new_n1780_ & ~new_n1781_;
  assign new_n1789_1_ = new_n1784_1_ & new_n1787_;
  assign n1134 = ~new_n1788_ | ~new_n1789_1_;
  assign new_n1791_ = n_n194 & new_n1157_;
  assign new_n1792_ = pkey_195_ & new_n1136_;
  assign new_n1793_ = n_n2396 & new_n1161_;
  assign new_n1794_1_ = n_n104 & new_n1164_1_;
  assign new_n1795_ = ~new_n1793_ & ~new_n1794_1_;
  assign new_n1796_ = n_n195 & new_n1168_;
  assign new_n1797_ = pkey_62_ & new_n1170_;
  assign new_n1798_ = ~new_n1796_ & ~new_n1797_;
  assign new_n1799_1_ = ~new_n1791_ & ~new_n1792_;
  assign new_n1800_ = new_n1795_ & new_n1798_;
  assign n1139 = ~new_n1799_1_ | ~new_n1800_;
  assign new_n1802_ = n_n109 & new_n1157_;
  assign new_n1803_ = n_n113 & new_n1161_;
  assign new_n1804_1_ = n_n112 & new_n1164_1_;
  assign new_n1805_ = ~new_n1803_ & ~new_n1804_1_;
  assign new_n1806_ = n_n110 & new_n1168_;
  assign new_n1807_ = pkey_228_ & new_n1170_;
  assign new_n1808_ = ~new_n1806_ & ~new_n1807_;
  assign new_n1809_1_ = ~new_n1298_ & ~new_n1802_;
  assign new_n1810_ = new_n1805_ & new_n1808_;
  assign n1144 = ~new_n1809_1_ | ~new_n1810_;
  assign new_n1812_ = n_n115 & new_n1157_;
  assign new_n1813_ = pkey_245_ & new_n1136_;
  assign new_n1814_1_ = n_n118 & new_n1161_;
  assign new_n1815_ = n_n117 & new_n1164_1_;
  assign new_n1816_ = ~new_n1814_1_ & ~new_n1815_;
  assign new_n1817_ = n_n116 & new_n1168_;
  assign new_n1818_ = pkey_237_ & new_n1170_;
  assign new_n1819_1_ = ~new_n1817_ & ~new_n1818_;
  assign new_n1820_ = ~new_n1812_ & ~new_n1813_;
  assign new_n1821_ = new_n1816_ & new_n1819_1_;
  assign n1149 = ~new_n1820_ | ~new_n1821_;
  assign new_n1823_ = n_n175 & new_n1157_;
  assign new_n1824_1_ = pkey_20_ & new_n1136_;
  assign new_n1825_ = n_n179 & new_n1161_;
  assign new_n1826_ = n_n178 & new_n1164_1_;
  assign new_n1827_ = ~new_n1825_ & ~new_n1826_;
  assign new_n1828_ = n_n176 & new_n1168_;
  assign new_n1829_1_ = pkey_12_ & new_n1170_;
  assign new_n1830_ = ~new_n1828_ & ~new_n1829_1_;
  assign new_n1831_ = ~new_n1823_ & ~new_n1824_1_;
  assign new_n1832_ = new_n1827_ & new_n1830_;
  assign n1154 = ~new_n1831_ | ~new_n1832_;
  assign new_n1834_1_ = n_n2507 & new_n1157_;
  assign new_n1835_ = pkey_29_ & new_n1136_;
  assign new_n1836_ = n_n187 & new_n1161_;
  assign new_n1837_ = n_n186 & new_n1164_1_;
  assign new_n1838_ = ~new_n1836_ & ~new_n1837_;
  assign new_n1839_1_ = n_n184 & new_n1168_;
  assign new_n1840_ = pkey_21_ & new_n1170_;
  assign new_n1841_ = ~new_n1839_1_ & ~new_n1840_;
  assign new_n1842_ = ~new_n1834_1_ & ~new_n1835_;
  assign new_n1843_ = new_n1838_ & new_n1841_;
  assign n1159 = ~new_n1842_ | ~new_n1843_;
  assign new_n1845_ = n_n190 & new_n1157_;
  assign new_n1846_ = pkey_38_ & new_n1136_;
  assign new_n1847_ = n_n194 & new_n1161_;
  assign new_n1848_ = n_n193 & new_n1164_1_;
  assign new_n1849_1_ = ~new_n1847_ & ~new_n1848_;
  assign new_n1850_ = n_n191 & new_n1168_;
  assign new_n1851_ = pkey_30_ & new_n1170_;
  assign new_n1852_ = ~new_n1850_ & ~new_n1851_;
  assign new_n1853_ = ~new_n1845_ & ~new_n1846_;
  assign new_n1854_1_ = new_n1849_1_ & new_n1852_;
  assign n1164 = ~new_n1853_ | ~new_n1854_1_;
  assign new_n1856_ = n_n2268 & new_n1157_;
  assign new_n1857_ = pkey_202_ & new_n1136_;
  assign new_n1858_ = n_n13 & new_n1161_;
  assign new_n1859_1_ = n_n2272 & new_n1164_1_;
  assign new_n1860_ = ~new_n1858_ & ~new_n1859_1_;
  assign new_n1861_ = n_n11 & new_n1168_;
  assign new_n1862_ = pkey_194_ & new_n1170_;
  assign new_n1863_ = ~new_n1861_ & ~new_n1862_;
  assign new_n1864_1_ = ~new_n1856_ & ~new_n1857_;
  assign new_n1865_ = new_n1860_ & new_n1863_;
  assign n1169 = ~new_n1864_1_ | ~new_n1865_;
  assign new_n1867_ = n_n123 & new_n1157_;
  assign new_n1868_ = pkey_131_ & new_n1136_;
  assign new_n1869_1_ = n_n2430 & new_n1161_;
  assign new_n1870_ = n_n126 & new_n1164_1_;
  assign new_n1871_ = ~new_n1869_1_ & ~new_n1870_;
  assign new_n1872_ = n_n124 & new_n1168_;
  assign new_n1873_ = pkey_254_ & new_n1170_;
  assign new_n1874_1_ = ~new_n1872_ & ~new_n1873_;
  assign new_n1875_ = ~new_n1867_ & ~new_n1868_;
  assign new_n1876_ = new_n1871_ & new_n1874_1_;
  assign n1174 = ~new_n1875_ | ~new_n1876_;
  assign new_n1878_ = n_n133 & new_n1157_;
  assign new_n1879_1_ = pkey_188_ & new_n1136_;
  assign new_n1880_ = n_n136 & new_n1161_;
  assign new_n1881_ = n_n135 & new_n1164_1_;
  assign new_n1882_ = ~new_n1880_ & ~new_n1881_;
  assign new_n1883_ = n_n134 & new_n1168_;
  assign new_n1884_1_ = pkey_180_ & new_n1170_;
  assign new_n1885_ = ~new_n1883_ & ~new_n1884_1_;
  assign new_n1886_ = ~new_n1878_ & ~new_n1879_1_;
  assign new_n1887_ = new_n1882_ & new_n1885_;
  assign n1179 = ~new_n1886_ | ~new_n1887_;
  assign new_n1889_1_ = n_n142 & new_n1157_;
  assign new_n1890_ = pkey_150_ & new_n1136_;
  assign new_n1891_ = n_n145 & new_n1161_;
  assign new_n1892_ = n_n144 & new_n1164_1_;
  assign new_n1893_ = ~new_n1891_ & ~new_n1892_;
  assign new_n1894_1_ = n_n2452 & new_n1168_;
  assign new_n1895_ = pkey_142_ & new_n1170_;
  assign new_n1896_ = ~new_n1894_1_ & ~new_n1895_;
  assign new_n1897_ = ~new_n1889_1_ & ~new_n1890_;
  assign new_n1898_ = new_n1893_ & new_n1896_;
  assign n1184 = ~new_n1897_ | ~new_n1898_;
  assign new_n1900_ = n_n151 & new_n1157_;
  assign new_n1901_ = pkey_76_ & new_n1136_;
  assign new_n1902_ = n_n155 & new_n1161_;
  assign new_n1903_ = n_n154 & new_n1164_1_;
  assign new_n1904_1_ = ~new_n1902_ & ~new_n1903_;
  assign new_n1905_ = n_n152 & new_n1168_;
  assign new_n1906_ = pkey_68_ & new_n1170_;
  assign new_n1907_ = ~new_n1905_ & ~new_n1906_;
  assign new_n1908_ = ~new_n1900_ & ~new_n1901_;
  assign new_n1909_1_ = new_n1904_1_ & new_n1907_;
  assign n1189 = ~new_n1908_ | ~new_n1909_1_;
  assign new_n1911_ = n_n2476 & new_n1157_;
  assign new_n1912_ = pkey_101_ & new_n1136_;
  assign new_n1913_ = n_n2481 & new_n1161_;
  assign new_n1914_1_ = n_n163 & new_n1164_1_;
  assign new_n1915_ = ~new_n1913_ & ~new_n1914_1_;
  assign new_n1916_ = n_n161 & new_n1168_;
  assign new_n1917_ = pkey_93_ & new_n1170_;
  assign new_n1918_ = ~new_n1916_ & ~new_n1917_;
  assign new_n1919_1_ = ~new_n1911_ & ~new_n1912_;
  assign new_n1920_ = new_n1915_ & new_n1918_;
  assign n1194 = ~new_n1919_1_ | ~new_n1920_;
  assign new_n1922_ = n_n169 & new_n1157_;
  assign new_n1923_ = pkey_126_ & new_n1136_;
  assign new_n1924_1_ = n_n173 & new_n1161_;
  assign new_n1925_ = n_n172 & new_n1164_1_;
  assign new_n1926_ = ~new_n1924_1_ & ~new_n1925_;
  assign new_n1927_ = n_n170 & new_n1168_;
  assign new_n1928_ = pkey_118_ & new_n1170_;
  assign new_n1929_1_ = ~new_n1927_ & ~new_n1928_;
  assign new_n1930_ = ~new_n1922_ & ~new_n1923_;
  assign new_n1931_ = new_n1926_ & new_n1929_1_;
  assign n1199 = ~new_n1930_ | ~new_n1931_;
  assign new_n1933_ = n_n11 & new_n1157_;
  assign new_n1934_1_ = pkey_210_ & new_n1136_;
  assign new_n1935_ = n_n14 & new_n1161_;
  assign new_n1936_ = n_n13 & new_n1164_1_;
  assign new_n1937_ = ~new_n1935_ & ~new_n1936_;
  assign new_n1938_ = n_n12 & new_n1168_;
  assign new_n1939_1_ = pkey_202_ & new_n1170_;
  assign new_n1940_ = ~new_n1938_ & ~new_n1939_1_;
  assign new_n1941_ = ~new_n1933_ & ~new_n1934_1_;
  assign new_n1942_ = new_n1937_ & new_n1940_;
  assign n1204 = ~new_n1941_ | ~new_n1942_;
  assign new_n1944_1_ = n_n124 & new_n1157_;
  assign new_n1945_ = pkey_139_ & new_n1136_;
  assign new_n1946_ = n_n127 & new_n1161_;
  assign new_n1947_ = n_n2430 & new_n1164_1_;
  assign new_n1948_ = ~new_n1946_ & ~new_n1947_;
  assign new_n1949_1_ = n_n125 & new_n1168_;
  assign new_n1950_ = pkey_131_ & new_n1170_;
  assign new_n1951_ = ~new_n1949_1_ & ~new_n1950_;
  assign new_n1952_ = ~new_n1944_1_ & ~new_n1945_;
  assign new_n1953_ = new_n1948_ & new_n1951_;
  assign n1209 = ~new_n1952_ | ~new_n1953_;
  assign new_n1955_ = n_n132 & new_n1157_;
  assign new_n1956_ = pkey_180_ & new_n1136_;
  assign new_n1957_ = n_n135 & new_n1161_;
  assign new_n1958_ = n_n2440 & new_n1164_1_;
  assign new_n1959_1_ = ~new_n1957_ & ~new_n1958_;
  assign new_n1960_ = n_n133 & new_n1168_;
  assign new_n1961_ = ~new_n1566_ & ~new_n1960_;
  assign new_n1962_ = ~new_n1955_ & ~new_n1956_;
  assign new_n1963_ = new_n1959_1_ & new_n1961_;
  assign n1214 = ~new_n1962_ | ~new_n1963_;
  assign new_n1965_ = n_n2452 & new_n1157_;
  assign new_n1966_ = pkey_158_ & new_n1136_;
  assign new_n1967_ = n_n146 & new_n1161_;
  assign new_n1968_ = n_n145 & new_n1164_1_;
  assign new_n1969_1_ = ~new_n1967_ & ~new_n1968_;
  assign new_n1970_ = n_n143 & new_n1168_;
  assign new_n1971_ = pkey_150_ & new_n1170_;
  assign new_n1972_ = ~new_n1970_ & ~new_n1971_;
  assign new_n1973_ = ~new_n1965_ & ~new_n1966_;
  assign new_n1974_ = new_n1969_1_ & new_n1972_;
  assign n1219 = ~new_n1973_ | ~new_n1974_;
  assign new_n1976_ = n_n2462 & new_n1157_;
  assign new_n1977_ = pkey_68_ & new_n1136_;
  assign new_n1978_ = n_n154 & new_n1161_;
  assign new_n1979_ = n_n153 & new_n1164_1_;
  assign new_n1980_ = ~new_n1978_ & ~new_n1979_;
  assign new_n1981_ = n_n151 & new_n1168_;
  assign new_n1982_ = pkey_91_ & new_n1170_;
  assign new_n1983_ = ~new_n1981_ & ~new_n1982_;
  assign new_n1984_ = ~new_n1976_ & ~new_n1977_;
  assign new_n1985_ = new_n1980_ & new_n1983_;
  assign n1224 = ~new_n1984_ | ~new_n1985_;
  assign new_n1987_ = n_n161 & new_n1157_;
  assign new_n1988_ = pkey_109_ & new_n1136_;
  assign new_n1989_ = n_n164 & new_n1161_;
  assign new_n1990_ = n_n2481 & new_n1164_1_;
  assign new_n1991_ = ~new_n1989_ & ~new_n1990_;
  assign new_n1992_ = n_n162 & new_n1168_;
  assign new_n1993_ = pkey_101_ & new_n1170_;
  assign new_n1994_ = ~new_n1992_ & ~new_n1993_;
  assign new_n1995_ = ~new_n1987_ & ~new_n1988_;
  assign new_n1996_ = new_n1991_ & new_n1994_;
  assign n1229 = ~new_n1995_ | ~new_n1996_;
  assign new_n1998_ = n_n168 & new_n1157_;
  assign new_n1999_ = pkey_118_ & new_n1136_;
  assign new_n2000_ = n_n172 & new_n1161_;
  assign new_n2001_ = n_n171 & new_n1164_1_;
  assign new_n2002_ = ~new_n2000_ & ~new_n2001_;
  assign new_n2003_ = n_n169 & new_n1168_;
  assign new_n2004_ = pkey_110_ & new_n1170_;
  assign new_n2005_ = ~new_n2003_ & ~new_n2004_;
  assign new_n2006_ = ~new_n1998_ & ~new_n1999_;
  assign new_n2007_ = new_n2002_ & new_n2005_;
  assign n1234 = ~new_n2006_ | ~new_n2007_;
  assign new_n2009_ = n_n12 & new_n1157_;
  assign new_n2010_ = pkey_218_ & new_n1136_;
  assign new_n2011_ = n_n15 & new_n1161_;
  assign new_n2012_ = n_n14 & new_n1164_1_;
  assign new_n2013_ = ~new_n2011_ & ~new_n2012_;
  assign new_n2014_ = n_n2272 & new_n1168_;
  assign new_n2015_ = pkey_210_ & new_n1170_;
  assign new_n2016_ = ~new_n2014_ & ~new_n2015_;
  assign new_n2017_ = ~new_n2009_ & ~new_n2010_;
  assign new_n2018_ = new_n2013_ & new_n2016_;
  assign n1239 = ~new_n2017_ | ~new_n2018_;
  assign new_n2020_ = n_n125 & new_n1157_;
  assign new_n2021_ = pkey_147_ & new_n1136_;
  assign new_n2022_ = n_n128 & new_n1161_;
  assign new_n2023_ = n_n127 & new_n1164_1_;
  assign new_n2024_ = ~new_n2022_ & ~new_n2023_;
  assign new_n2025_ = n_n126 & new_n1168_;
  assign new_n2026_ = pkey_139_ & new_n1170_;
  assign new_n2027_ = ~new_n2025_ & ~new_n2026_;
  assign new_n2028_ = ~new_n2020_ & ~new_n2021_;
  assign new_n2029_ = new_n2024_ & new_n2027_;
  assign n1244 = ~new_n2028_ | ~new_n2029_;
  assign new_n2031_ = n_n2440 & new_n1157_;
  assign new_n2032_ = pkey_141_ & new_n1136_;
  assign new_n2033_ = n_n138 & new_n1161_;
  assign new_n2034_ = n_n137 & new_n1164_1_;
  assign new_n2035_ = ~new_n2033_ & ~new_n2034_;
  assign new_n2036_ = n_n135 & new_n1168_;
  assign new_n2037_ = pkey_133_ & new_n1170_;
  assign new_n2038_ = ~new_n2036_ & ~new_n2037_;
  assign new_n2039_ = ~new_n2031_ & ~new_n2032_;
  assign new_n2040_ = new_n2035_ & new_n2038_;
  assign n1249 = ~new_n2039_ | ~new_n2040_;
  assign new_n2042_ = n_n2448 & new_n1157_;
  assign new_n2043_ = pkey_134_ & new_n1136_;
  assign new_n2044_ = n_n143 & new_n1161_;
  assign new_n2045_ = n_n2452 & new_n1164_1_;
  assign new_n2046_ = ~new_n2044_ & ~new_n2045_;
  assign new_n2047_ = n_n141 & new_n1168_;
  assign new_n2048_ = pkey_189_ & new_n1170_;
  assign new_n2049_ = ~new_n2047_ & ~new_n2048_;
  assign new_n2050_ = ~new_n2042_ & ~new_n2043_;
  assign new_n2051_ = new_n2046_ & new_n2049_;
  assign n1254 = ~new_n2050_ | ~new_n2051_;
  assign new_n2053_ = n_n150 & new_n1157_;
  assign new_n2054_ = pkey_91_ & new_n1136_;
  assign new_n2055_ = n_n153 & new_n1161_;
  assign new_n2056_ = n_n152 & new_n1164_1_;
  assign new_n2057_ = ~new_n2055_ & ~new_n2056_;
  assign new_n2058_ = n_n2462 & new_n1168_;
  assign new_n2059_ = pkey_83_ & new_n1170_;
  assign new_n2060_ = ~new_n2058_ & ~new_n2059_;
  assign new_n2061_ = ~new_n2053_ & ~new_n2054_;
  assign new_n2062_ = new_n2057_ & new_n2060_;
  assign n1259 = ~new_n2061_ | ~new_n2062_;
  assign new_n2064_ = n_n162 & new_n1157_;
  assign new_n2065_ = pkey_117_ & new_n1136_;
  assign new_n2066_ = n_n165 & new_n1161_;
  assign new_n2067_ = n_n164 & new_n1164_1_;
  assign new_n2068_ = ~new_n2066_ & ~new_n2067_;
  assign new_n2069_ = n_n163 & new_n1168_;
  assign new_n2070_ = pkey_109_ & new_n1170_;
  assign new_n2071_ = ~new_n2069_ & ~new_n2070_;
  assign new_n2072_ = ~new_n2064_ & ~new_n2065_;
  assign new_n2073_ = new_n2068_ & new_n2071_;
  assign n1264 = ~new_n2072_ | ~new_n2073_;
  assign new_n2075_ = n_n171 & new_n1157_;
  assign new_n2076_ = pkey_11_ & new_n1136_;
  assign new_n2077_ = n_n174 & new_n1161_;
  assign new_n2078_ = n_n2495 & new_n1164_1_;
  assign new_n2079_ = ~new_n2077_ & ~new_n2078_;
  assign new_n2080_ = n_n172 & new_n1168_;
  assign new_n2081_ = pkey_3_ & new_n1170_;
  assign new_n2082_ = ~new_n2080_ & ~new_n2081_;
  assign new_n2083_ = ~new_n2075_ & ~new_n2076_;
  assign new_n2084_ = new_n2079_ & new_n2082_;
  assign n1269 = ~new_n2083_ | ~new_n2084_;
  assign new_n2086_ = n_n2272 & new_n1157_;
  assign new_n2087_ = pkey_226_ & new_n1136_;
  assign new_n2088_ = n_n2277 & new_n1161_;
  assign new_n2089_ = n_n15 & new_n1164_1_;
  assign new_n2090_ = ~new_n2088_ & ~new_n2089_;
  assign new_n2091_ = n_n13 & new_n1168_;
  assign new_n2092_ = pkey_218_ & new_n1170_;
  assign new_n2093_ = ~new_n2091_ & ~new_n2092_;
  assign new_n2094_ = ~new_n2086_ & ~new_n2087_;
  assign new_n2095_ = new_n2090_ & new_n2093_;
  assign n1274 = ~new_n2094_ | ~new_n2095_;
  assign new_n2097_ = n_n126 & new_n1157_;
  assign new_n2098_ = pkey_155_ & new_n1136_;
  assign new_n2099_ = n_n129 & new_n1161_;
  assign new_n2100_ = n_n128 & new_n1164_1_;
  assign new_n2101_ = ~new_n2099_ & ~new_n2100_;
  assign new_n2102_ = n_n2430 & new_n1168_;
  assign new_n2103_ = pkey_147_ & new_n1170_;
  assign new_n2104_ = ~new_n2102_ & ~new_n2103_;
  assign new_n2105_ = ~new_n2097_ & ~new_n2098_;
  assign new_n2106_ = new_n2101_ & new_n2104_;
  assign n1279 = ~new_n2105_ | ~new_n2106_;
  assign new_n2108_ = n_n134 & new_n1157_;
  assign new_n2109_ = pkey_133_ & new_n1136_;
  assign new_n2110_ = n_n137 & new_n1161_;
  assign new_n2111_ = n_n136 & new_n1164_1_;
  assign new_n2112_ = ~new_n2110_ & ~new_n2111_;
  assign new_n2113_ = n_n2440 & new_n1168_;
  assign new_n2114_ = pkey_188_ & new_n1170_;
  assign new_n2115_ = ~new_n2113_ & ~new_n2114_;
  assign new_n2116_ = ~new_n2108_ & ~new_n2109_;
  assign new_n2117_ = new_n2112_ & new_n2115_;
  assign n1284 = ~new_n2116_ | ~new_n2117_;
  assign new_n2119_ = n_n141 & new_n1157_;
  assign new_n2120_ = pkey_142_ & new_n1136_;
  assign new_n2121_ = n_n144 & new_n1161_;
  assign new_n2122_ = n_n143 & new_n1164_1_;
  assign new_n2123_ = ~new_n2121_ & ~new_n2122_;
  assign new_n2124_ = n_n142 & new_n1168_;
  assign new_n2125_ = pkey_134_ & new_n1170_;
  assign new_n2126_ = ~new_n2124_ & ~new_n2125_;
  assign new_n2127_ = ~new_n2119_ & ~new_n2120_;
  assign new_n2128_ = new_n2123_ & new_n2126_;
  assign n1289 = ~new_n2127_ | ~new_n2128_;
  assign new_n2130_ = n_n149 & new_n1157_;
  assign new_n2131_ = pkey_83_ & new_n1136_;
  assign new_n2132_ = n_n152 & new_n1161_;
  assign new_n2133_ = n_n151 & new_n1164_1_;
  assign new_n2134_ = ~new_n2132_ & ~new_n2133_;
  assign new_n2135_ = n_n150 & new_n1168_;
  assign new_n2136_ = pkey_75_ & new_n1170_;
  assign new_n2137_ = ~new_n2135_ & ~new_n2136_;
  assign new_n2138_ = ~new_n2130_ & ~new_n2131_;
  assign new_n2139_ = new_n2134_ & new_n2137_;
  assign n1294 = ~new_n2138_ | ~new_n2139_;
  assign new_n2141_ = n_n163 & new_n1157_;
  assign new_n2142_ = pkey_125_ & new_n1136_;
  assign new_n2143_ = n_n2485 & new_n1161_;
  assign new_n2144_ = n_n165 & new_n1164_1_;
  assign new_n2145_ = ~new_n2143_ & ~new_n2144_;
  assign new_n2146_ = n_n2481 & new_n1168_;
  assign new_n2147_ = pkey_117_ & new_n1170_;
  assign new_n2148_ = ~new_n2146_ & ~new_n2147_;
  assign new_n2149_ = ~new_n2141_ & ~new_n2142_;
  assign new_n2150_ = new_n2145_ & new_n2148_;
  assign n1299 = ~new_n2149_ | ~new_n2150_;
  assign new_n2152_ = n_n170 & new_n1157_;
  assign new_n2153_ = pkey_3_ & new_n1136_;
  assign new_n2154_ = n_n2495 & new_n1161_;
  assign new_n2155_ = n_n173 & new_n1164_1_;
  assign new_n2156_ = ~new_n2154_ & ~new_n2155_;
  assign new_n2157_ = n_n171 & new_n1168_;
  assign new_n2158_ = pkey_126_ & new_n1170_;
  assign new_n2159_ = ~new_n2157_ & ~new_n2158_;
  assign new_n2160_ = ~new_n2152_ & ~new_n2153_;
  assign new_n2161_ = new_n2156_ & new_n2159_;
  assign n1304 = ~new_n2160_ | ~new_n2161_;
  assign new_n2163_ = n_n102 & new_n1157_;
  assign new_n2164_ = pkey_235_ & new_n1136_;
  assign new_n2165_ = n_n2268 & new_n1161_;
  assign new_n2166_ = n_n10 & new_n1164_1_;
  assign new_n2167_ = ~new_n2165_ & ~new_n2166_;
  assign new_n2168_ = n_n8 & new_n1168_;
  assign new_n2169_ = pkey_227_ & new_n1170_;
  assign new_n2170_ = ~new_n2168_ & ~new_n2169_;
  assign new_n2171_ = ~new_n2163_ & ~new_n2164_;
  assign new_n2172_ = new_n2167_ & new_n2170_;
  assign n1309 = ~new_n2171_ | ~new_n2172_;
  assign new_n2174_ = n_n97 & new_n1157_;
  assign new_n2175_ = pkey_32_ & new_n1136_;
  assign new_n2176_ = n_n101 & new_n1161_;
  assign new_n2177_ = n_n100 & new_n1164_1_;
  assign new_n2178_ = ~new_n2176_ & ~new_n2177_;
  assign new_n2179_ = n_n98 & new_n1168_;
  assign new_n2180_ = pkey_24_ & new_n1170_;
  assign new_n2181_ = ~new_n2179_ & ~new_n2180_;
  assign new_n2182_ = ~new_n2174_ & ~new_n2175_;
  assign new_n2183_ = new_n2178_ & new_n2181_;
  assign n1314 = ~new_n2182_ | ~new_n2183_;
  assign new_n2185_ = n_n107 & new_n1157_;
  assign new_n2186_ = pkey_220_ & new_n1136_;
  assign new_n2187_ = n_n111 & new_n1161_;
  assign new_n2188_ = n_n110 & new_n1164_1_;
  assign new_n2189_ = ~new_n2187_ & ~new_n2188_;
  assign new_n2190_ = n_n108 & new_n1168_;
  assign new_n2191_ = pkey_212_ & new_n1170_;
  assign new_n2192_ = ~new_n2190_ & ~new_n2191_;
  assign new_n2193_ = ~new_n2185_ & ~new_n2186_;
  assign new_n2194_ = new_n2189_ & new_n2192_;
  assign n1319 = ~new_n2193_ | ~new_n2194_;
  assign new_n2196_ = n_n2430 & new_n1157_;
  assign new_n2197_ = pkey_132_ & new_n1136_;
  assign new_n2198_ = n_n130 & new_n1161_;
  assign new_n2199_ = n_n129 & new_n1164_1_;
  assign new_n2200_ = ~new_n2198_ & ~new_n2199_;
  assign new_n2201_ = n_n127 & new_n1168_;
  assign new_n2202_ = pkey_155_ & new_n1170_;
  assign new_n2203_ = ~new_n2201_ & ~new_n2202_;
  assign new_n2204_ = ~new_n2196_ & ~new_n2197_;
  assign new_n2205_ = new_n2200_ & new_n2203_;
  assign n1324 = ~new_n2204_ | ~new_n2205_;
  assign new_n2207_ = n_n136 & new_n1157_;
  assign new_n2208_ = pkey_157_ & new_n1136_;
  assign new_n2209_ = n_n140 & new_n1161_;
  assign new_n2210_ = n_n139 & new_n1164_1_;
  assign new_n2211_ = ~new_n2209_ & ~new_n2210_;
  assign new_n2212_ = n_n137 & new_n1168_;
  assign new_n2213_ = pkey_149_ & new_n1170_;
  assign new_n2214_ = ~new_n2212_ & ~new_n2213_;
  assign new_n2215_ = ~new_n2207_ & ~new_n2208_;
  assign new_n2216_ = new_n2211_ & new_n2214_;
  assign n1329 = ~new_n2215_ | ~new_n2216_;
  assign new_n2218_ = n_n145 & new_n1157_;
  assign new_n2219_ = pkey_182_ & new_n1136_;
  assign new_n2220_ = n_n149 & new_n1161_;
  assign new_n2221_ = n_n148 & new_n1164_1_;
  assign new_n2222_ = ~new_n2220_ & ~new_n2221_;
  assign new_n2223_ = n_n146 & new_n1168_;
  assign new_n2224_ = pkey_174_ & new_n1170_;
  assign new_n2225_ = ~new_n2223_ & ~new_n2224_;
  assign new_n2226_ = ~new_n2218_ & ~new_n2219_;
  assign new_n2227_ = new_n2222_ & new_n2225_;
  assign n1334 = ~new_n2226_ | ~new_n2227_;
  assign new_n2229_ = n_n155 & new_n1157_;
  assign new_n2230_ = n_n159 & new_n1161_;
  assign new_n2231_ = n_n158 & new_n1164_1_;
  assign new_n2232_ = ~new_n2230_ & ~new_n2231_;
  assign new_n2233_ = n_n156 & new_n1168_;
  assign new_n2234_ = pkey_100_ & new_n1170_;
  assign new_n2235_ = ~new_n2233_ & ~new_n2234_;
  assign new_n2236_ = ~new_n1408_ & ~new_n2229_;
  assign new_n2237_ = new_n2232_ & new_n2235_;
  assign n1339 = ~new_n2236_ | ~new_n2237_;
  assign new_n2239_ = n_n158 & new_n1157_;
  assign new_n2240_ = pkey_69_ & new_n1136_;
  assign new_n2241_ = n_n2476 & new_n1161_;
  assign new_n2242_ = n_n2474 & new_n1164_1_;
  assign new_n2243_ = ~new_n2241_ & ~new_n2242_;
  assign new_n2244_ = n_n159 & new_n1168_;
  assign new_n2245_ = pkey_124_ & new_n1170_;
  assign new_n2246_ = ~new_n2244_ & ~new_n2245_;
  assign new_n2247_ = ~new_n2239_ & ~new_n2240_;
  assign new_n2248_ = new_n2243_ & new_n2246_;
  assign n1344 = ~new_n2247_ | ~new_n2248_;
  assign new_n2250_ = n_n2485 & new_n1157_;
  assign new_n2251_ = pkey_94_ & new_n1136_;
  assign new_n2252_ = n_n169 & new_n1161_;
  assign new_n2253_ = n_n168 & new_n1164_1_;
  assign new_n2254_ = ~new_n2252_ & ~new_n2253_;
  assign new_n2255_ = n_n166 & new_n1168_;
  assign new_n2256_ = pkey_86_ & new_n1170_;
  assign new_n2257_ = ~new_n2255_ & ~new_n2256_;
  assign new_n2258_ = ~new_n2250_ & ~new_n2251_;
  assign new_n2259_ = new_n2254_ & new_n2257_;
  assign n1349 = ~new_n2258_ | ~new_n2259_;
  assign new_n2261_ = n_n180 & new_n1157_;
  assign new_n2262_ = pkey_60_ & new_n1136_;
  assign new_n2263_ = n_n2507 & new_n1161_;
  assign new_n2264_ = n_n183 & new_n1164_1_;
  assign new_n2265_ = ~new_n2263_ & ~new_n2264_;
  assign new_n2266_ = n_n181 & new_n1168_;
  assign new_n2267_ = pkey_52_ & new_n1170_;
  assign new_n2268_ = ~new_n2266_ & ~new_n2267_;
  assign new_n2269_ = ~new_n2261_ & ~new_n2262_;
  assign new_n2270_ = new_n2265_ & new_n2268_;
  assign n1354 = ~new_n2269_ | ~new_n2270_;
  assign new_n2272_ = n_n189 & new_n1157_;
  assign new_n2273_ = pkey_22_ & new_n1136_;
  assign new_n2274_ = n_n192 & new_n1161_;
  assign new_n2275_ = n_n191 & new_n1164_1_;
  assign new_n2276_ = ~new_n2274_ & ~new_n2275_;
  assign new_n2277_ = n_n2517 & new_n1168_;
  assign new_n2278_ = pkey_14_ & new_n1170_;
  assign new_n2279_ = ~new_n2277_ & ~new_n2278_;
  assign new_n2280_ = ~new_n2272_ & ~new_n2273_;
  assign new_n2281_ = new_n2276_ & new_n2279_;
  assign n1359 = ~new_n2280_ | ~new_n2281_;
  assign new_n2283_ = n_n8 & new_n1157_;
  assign new_n2284_ = pkey_243_ & new_n1136_;
  assign new_n2285_ = n_n11 & new_n1161_;
  assign new_n2286_ = n_n2268 & new_n1164_1_;
  assign new_n2287_ = ~new_n2285_ & ~new_n2286_;
  assign new_n2288_ = n_n9 & new_n1168_;
  assign new_n2289_ = pkey_235_ & new_n1170_;
  assign new_n2290_ = ~new_n2288_ & ~new_n2289_;
  assign new_n2291_ = ~new_n2283_ & ~new_n2284_;
  assign new_n2292_ = new_n2287_ & new_n2290_;
  assign n1364 = ~new_n2291_ | ~new_n2292_;
  assign new_n2294_ = n_n98 & new_n1157_;
  assign new_n2295_ = pkey_40_ & new_n1136_;
  assign new_n2296_ = n_n102 & new_n1161_;
  assign new_n2297_ = n_n101 & new_n1164_1_;
  assign new_n2298_ = ~new_n2296_ & ~new_n2297_;
  assign new_n2299_ = n_n99 & new_n1168_;
  assign new_n2300_ = pkey_32_ & new_n1170_;
  assign new_n2301_ = ~new_n2299_ & ~new_n2300_;
  assign new_n2302_ = ~new_n2294_ & ~new_n2295_;
  assign new_n2303_ = new_n2298_ & new_n2301_;
  assign n1369 = ~new_n2302_ | ~new_n2303_;
  assign new_n2305_ = n_n106 & new_n1157_;
  assign new_n2306_ = pkey_212_ & new_n1136_;
  assign new_n2307_ = n_n110 & new_n1161_;
  assign new_n2308_ = n_n109 & new_n1164_1_;
  assign new_n2309_ = ~new_n2307_ & ~new_n2308_;
  assign new_n2310_ = n_n107 & new_n1168_;
  assign new_n2311_ = pkey_204_ & new_n1170_;
  assign new_n2312_ = ~new_n2310_ & ~new_n2311_;
  assign new_n2313_ = ~new_n2305_ & ~new_n2306_;
  assign new_n2314_ = new_n2309_ & new_n2312_;
  assign n1374 = ~new_n2313_ | ~new_n2314_;
  assign new_n2316_ = n_n127 & new_n1157_;
  assign new_n2317_ = pkey_140_ & new_n1136_;
  assign new_n2318_ = n_n131 & new_n1161_;
  assign new_n2319_ = n_n130 & new_n1164_1_;
  assign new_n2320_ = ~new_n2318_ & ~new_n2319_;
  assign new_n2321_ = n_n128 & new_n1168_;
  assign new_n2322_ = pkey_132_ & new_n1170_;
  assign new_n2323_ = ~new_n2321_ & ~new_n2322_;
  assign new_n2324_ = ~new_n2316_ & ~new_n2317_;
  assign new_n2325_ = new_n2320_ & new_n2323_;
  assign n1379 = ~new_n2324_ | ~new_n2325_;
  assign new_n2327_ = n_n135 & new_n1157_;
  assign new_n2328_ = pkey_149_ & new_n1136_;
  assign new_n2329_ = n_n139 & new_n1161_;
  assign new_n2330_ = n_n138 & new_n1164_1_;
  assign new_n2331_ = ~new_n2329_ & ~new_n2330_;
  assign new_n2332_ = n_n136 & new_n1168_;
  assign new_n2333_ = pkey_141_ & new_n1170_;
  assign new_n2334_ = ~new_n2332_ & ~new_n2333_;
  assign new_n2335_ = ~new_n2327_ & ~new_n2328_;
  assign new_n2336_ = new_n2331_ & new_n2334_;
  assign n1384 = ~new_n2335_ | ~new_n2336_;
  assign new_n2338_ = n_n146 & new_n1157_;
  assign new_n2339_ = pkey_190_ & new_n1136_;
  assign new_n2340_ = n_n150 & new_n1161_;
  assign new_n2341_ = n_n149 & new_n1164_1_;
  assign new_n2342_ = ~new_n2340_ & ~new_n2341_;
  assign new_n2343_ = n_n147 & new_n1168_;
  assign new_n2344_ = pkey_182_ & new_n1170_;
  assign new_n2345_ = ~new_n2343_ & ~new_n2344_;
  assign new_n2346_ = ~new_n2338_ & ~new_n2339_;
  assign new_n2347_ = new_n2342_ & new_n2345_;
  assign n1389 = ~new_n2346_ | ~new_n2347_;
  assign new_n2349_ = n_n154 & new_n1157_;
  assign new_n2350_ = pkey_100_ & new_n1136_;
  assign new_n2351_ = n_n158 & new_n1161_;
  assign new_n2352_ = n_n157 & new_n1164_1_;
  assign new_n2353_ = ~new_n2351_ & ~new_n2352_;
  assign new_n2354_ = n_n155 & new_n1168_;
  assign new_n2355_ = pkey_92_ & new_n1170_;
  assign new_n2356_ = ~new_n2354_ & ~new_n2355_;
  assign new_n2357_ = ~new_n2349_ & ~new_n2350_;
  assign new_n2358_ = new_n2353_ & new_n2356_;
  assign n1394 = ~new_n2357_ | ~new_n2358_;
  assign new_n2360_ = n_n159 & new_n1157_;
  assign new_n2361_ = pkey_77_ & new_n1136_;
  assign new_n2362_ = n_n161 & new_n1161_;
  assign new_n2363_ = n_n2476 & new_n1164_1_;
  assign new_n2364_ = ~new_n2362_ & ~new_n2363_;
  assign new_n2365_ = n_n160 & new_n1168_;
  assign new_n2366_ = pkey_69_ & new_n1170_;
  assign new_n2367_ = ~new_n2365_ & ~new_n2366_;
  assign new_n2368_ = ~new_n2360_ & ~new_n2361_;
  assign new_n2369_ = new_n2364_ & new_n2367_;
  assign n1399 = ~new_n2368_ | ~new_n2369_;
  assign new_n2371_ = n_n165 & new_n1157_;
  assign new_n2372_ = pkey_86_ & new_n1136_;
  assign new_n2373_ = n_n168 & new_n1161_;
  assign new_n2374_ = n_n167 & new_n1164_1_;
  assign new_n2375_ = ~new_n2373_ & ~new_n2374_;
  assign new_n2376_ = n_n2485 & new_n1168_;
  assign new_n2377_ = pkey_78_ & new_n1170_;
  assign new_n2378_ = ~new_n2376_ & ~new_n2377_;
  assign new_n2379_ = ~new_n2371_ & ~new_n2372_;
  assign new_n2380_ = new_n2375_ & new_n2378_;
  assign n1404 = ~new_n2379_ | ~new_n2380_;
  assign new_n2382_ = n_n181 & new_n1157_;
  assign new_n2383_ = pkey_5_ & new_n1136_;
  assign new_n2384_ = n_n184 & new_n1161_;
  assign new_n2385_ = n_n2507 & new_n1164_1_;
  assign new_n2386_ = ~new_n2384_ & ~new_n2385_;
  assign new_n2387_ = n_n182 & new_n1168_;
  assign new_n2388_ = pkey_60_ & new_n1170_;
  assign new_n2389_ = ~new_n2387_ & ~new_n2388_;
  assign new_n2390_ = ~new_n2382_ & ~new_n2383_;
  assign new_n2391_ = new_n2386_ & new_n2389_;
  assign n1409 = ~new_n2390_ | ~new_n2391_;
  assign new_n2393_ = n_n188 & new_n1157_;
  assign new_n2394_ = pkey_14_ & new_n1136_;
  assign new_n2395_ = n_n191 & new_n1161_;
  assign new_n2396_ = n_n190 & new_n1164_1_;
  assign new_n2397_ = ~new_n2395_ & ~new_n2396_;
  assign new_n2398_ = n_n189 & new_n1168_;
  assign new_n2399_ = pkey_6_ & new_n1170_;
  assign new_n2400_ = ~new_n2398_ & ~new_n2399_;
  assign new_n2401_ = ~new_n2393_ & ~new_n2394_;
  assign new_n2402_ = new_n2397_ & new_n2400_;
  assign n1414 = ~new_n2401_ | ~new_n2402_;
  assign new_n2404_ = n_n9 & new_n1157_;
  assign new_n2405_ = pkey_251_ & new_n1136_;
  assign new_n2406_ = n_n12 & new_n1161_;
  assign new_n2407_ = n_n11 & new_n1164_1_;
  assign new_n2408_ = ~new_n2406_ & ~new_n2407_;
  assign new_n2409_ = n_n10 & new_n1168_;
  assign new_n2410_ = pkey_243_ & new_n1170_;
  assign new_n2411_ = ~new_n2409_ & ~new_n2410_;
  assign new_n2412_ = ~new_n2404_ & ~new_n2405_;
  assign new_n2413_ = new_n2408_ & new_n2411_;
  assign n1419 = ~new_n2412_ | ~new_n2413_;
  assign new_n2415_ = n_n2410 & new_n1157_;
  assign new_n2416_ = pkey_229_ & new_n1136_;
  assign new_n2417_ = n_n2416 & new_n1161_;
  assign new_n2418_ = n_n116 & new_n1164_1_;
  assign new_n2419_ = ~new_n2417_ & ~new_n2418_;
  assign new_n2420_ = n_n2412 & new_n1168_;
  assign new_n2421_ = pkey_221_ & new_n1170_;
  assign new_n2422_ = ~new_n2420_ & ~new_n2421_;
  assign new_n2423_ = ~new_n2415_ & ~new_n2416_;
  assign new_n2424_ = new_n2419_ & new_n2422_;
  assign n1424 = ~new_n2423_ | ~new_n2424_;
  assign new_n2426_ = n_n122 & new_n1157_;
  assign new_n2427_ = pkey_254_ & new_n1136_;
  assign new_n2428_ = n_n126 & new_n1161_;
  assign new_n2429_ = n_n125 & new_n1164_1_;
  assign new_n2430_ = ~new_n2428_ & ~new_n2429_;
  assign new_n2431_ = n_n123 & new_n1168_;
  assign new_n2432_ = pkey_246_ & new_n1170_;
  assign new_n2433_ = ~new_n2431_ & ~new_n2432_;
  assign new_n2434_ = ~new_n2426_ & ~new_n2427_;
  assign new_n2435_ = new_n2430_ & new_n2433_;
  assign n1429 = ~new_n2434_ | ~new_n2435_;
  assign new_n2437_ = n_n128 & new_n1157_;
  assign new_n2438_ = pkey_148_ & new_n1136_;
  assign new_n2439_ = n_n132 & new_n1161_;
  assign new_n2440_ = n_n131 & new_n1164_1_;
  assign new_n2441_ = ~new_n2439_ & ~new_n2440_;
  assign new_n2442_ = n_n129 & new_n1168_;
  assign new_n2443_ = pkey_140_ & new_n1170_;
  assign new_n2444_ = ~new_n2442_ & ~new_n2443_;
  assign new_n2445_ = ~new_n2437_ & ~new_n2438_;
  assign new_n2446_ = new_n2441_ & new_n2444_;
  assign n1434 = ~new_n2445_ | ~new_n2446_;
  assign new_n2448_ = n_n138 & new_n1157_;
  assign new_n2449_ = pkey_173_ & new_n1136_;
  assign new_n2450_ = n_n141 & new_n1161_;
  assign new_n2451_ = n_n2448 & new_n1164_1_;
  assign new_n2452_ = ~new_n2450_ & ~new_n2451_;
  assign new_n2453_ = n_n139 & new_n1168_;
  assign new_n2454_ = pkey_165_ & new_n1170_;
  assign new_n2455_ = ~new_n2453_ & ~new_n2454_;
  assign new_n2456_ = ~new_n2448_ & ~new_n2449_;
  assign new_n2457_ = new_n2452_ & new_n2455_;
  assign n1439 = ~new_n2456_ | ~new_n2457_;
  assign new_n2459_ = n_n143 & new_n1157_;
  assign new_n2460_ = pkey_166_ & new_n1136_;
  assign new_n2461_ = n_n147 & new_n1161_;
  assign new_n2462_ = n_n146 & new_n1164_1_;
  assign new_n2463_ = ~new_n2461_ & ~new_n2462_;
  assign new_n2464_ = n_n144 & new_n1168_;
  assign new_n2465_ = pkey_158_ & new_n1170_;
  assign new_n2466_ = ~new_n2464_ & ~new_n2465_;
  assign new_n2467_ = ~new_n2459_ & ~new_n2460_;
  assign new_n2468_ = new_n2463_ & new_n2466_;
  assign n1444 = ~new_n2467_ | ~new_n2468_;
  assign new_n2470_ = n_n153 & new_n1157_;
  assign new_n2471_ = pkey_92_ & new_n1136_;
  assign new_n2472_ = n_n157 & new_n1161_;
  assign new_n2473_ = n_n156 & new_n1164_1_;
  assign new_n2474_ = ~new_n2472_ & ~new_n2473_;
  assign new_n2475_ = n_n154 & new_n1168_;
  assign new_n2476_ = pkey_84_ & new_n1170_;
  assign new_n2477_ = ~new_n2475_ & ~new_n2476_;
  assign new_n2478_ = ~new_n2470_ & ~new_n2471_;
  assign new_n2479_ = new_n2474_ & new_n2477_;
  assign n1449 = ~new_n2478_ | ~new_n2479_;
  assign new_n2481_ = n_n160 & new_n1157_;
  assign new_n2482_ = pkey_85_ & new_n1136_;
  assign new_n2483_ = n_n162 & new_n1161_;
  assign new_n2484_ = n_n161 & new_n1164_1_;
  assign new_n2485_ = ~new_n2483_ & ~new_n2484_;
  assign new_n2486_ = n_n2474 & new_n1168_;
  assign new_n2487_ = pkey_77_ & new_n1170_;
  assign new_n2488_ = ~new_n2486_ & ~new_n2487_;
  assign new_n2489_ = ~new_n2481_ & ~new_n2482_;
  assign new_n2490_ = new_n2485_ & new_n2488_;
  assign n1454 = ~new_n2489_ | ~new_n2490_;
  assign new_n2492_ = n_n167 & new_n1157_;
  assign new_n2493_ = pkey_110_ & new_n1136_;
  assign new_n2494_ = n_n171 & new_n1161_;
  assign new_n2495_ = n_n170 & new_n1164_1_;
  assign new_n2496_ = ~new_n2494_ & ~new_n2495_;
  assign new_n2497_ = n_n168 & new_n1168_;
  assign new_n2498_ = pkey_102_ & new_n1170_;
  assign new_n2499_ = ~new_n2497_ & ~new_n2498_;
  assign new_n2500_ = ~new_n2492_ & ~new_n2493_;
  assign new_n2501_ = new_n2496_ & new_n2499_;
  assign n1459 = ~new_n2500_ | ~new_n2501_;
  assign new_n2503_ = n_n182 & new_n1157_;
  assign new_n2504_ = pkey_13_ & new_n1136_;
  assign new_n2505_ = n_n185 & new_n1161_;
  assign new_n2506_ = n_n184 & new_n1164_1_;
  assign new_n2507_ = ~new_n2505_ & ~new_n2506_;
  assign new_n2508_ = n_n183 & new_n1168_;
  assign new_n2509_ = pkey_5_ & new_n1170_;
  assign new_n2510_ = ~new_n2508_ & ~new_n2509_;
  assign new_n2511_ = ~new_n2503_ & ~new_n2504_;
  assign new_n2512_ = new_n2507_ & new_n2510_;
  assign n1464 = ~new_n2511_ | ~new_n2512_;
  assign new_n2514_ = n_n10 & new_n1157_;
  assign new_n2515_ = pkey_194_ & new_n1136_;
  assign new_n2516_ = n_n2272 & new_n1161_;
  assign new_n2517_ = n_n12 & new_n1164_1_;
  assign new_n2518_ = ~new_n2516_ & ~new_n2517_;
  assign new_n2519_ = n_n2268 & new_n1168_;
  assign new_n2520_ = pkey_251_ & new_n1170_;
  assign new_n2521_ = ~new_n2519_ & ~new_n2520_;
  assign new_n2522_ = ~new_n2514_ & ~new_n2515_;
  assign new_n2523_ = new_n2518_ & new_n2521_;
  assign n1469 = ~new_n2522_ | ~new_n2523_;
  assign new_n2525_ = n_n2412 & new_n1157_;
  assign new_n2526_ = pkey_237_ & new_n1136_;
  assign new_n2527_ = n_n117 & new_n1161_;
  assign new_n2528_ = n_n2416 & new_n1164_1_;
  assign new_n2529_ = ~new_n2527_ & ~new_n2528_;
  assign new_n2530_ = n_n115 & new_n1168_;
  assign new_n2531_ = pkey_229_ & new_n1170_;
  assign new_n2532_ = ~new_n2530_ & ~new_n2531_;
  assign new_n2533_ = ~new_n2525_ & ~new_n2526_;
  assign new_n2534_ = new_n2529_ & new_n2532_;
  assign n1474 = ~new_n2533_ | ~new_n2534_;
  assign new_n2536_ = n_n121 & new_n1157_;
  assign new_n2537_ = pkey_246_ & new_n1136_;
  assign new_n2538_ = n_n125 & new_n1161_;
  assign new_n2539_ = n_n124 & new_n1164_1_;
  assign new_n2540_ = ~new_n2538_ & ~new_n2539_;
  assign new_n2541_ = n_n122 & new_n1168_;
  assign new_n2542_ = pkey_238_ & new_n1170_;
  assign new_n2543_ = ~new_n2541_ & ~new_n2542_;
  assign new_n2544_ = ~new_n2536_ & ~new_n2537_;
  assign new_n2545_ = new_n2540_ & new_n2543_;
  assign n1479 = ~new_n2544_ | ~new_n2545_;
  assign new_n2547_ = n_n129 & new_n1157_;
  assign new_n2548_ = pkey_156_ & new_n1136_;
  assign new_n2549_ = n_n133 & new_n1161_;
  assign new_n2550_ = n_n132 & new_n1164_1_;
  assign new_n2551_ = ~new_n2549_ & ~new_n2550_;
  assign new_n2552_ = n_n130 & new_n1168_;
  assign new_n2553_ = pkey_148_ & new_n1170_;
  assign new_n2554_ = ~new_n2552_ & ~new_n2553_;
  assign new_n2555_ = ~new_n2547_ & ~new_n2548_;
  assign new_n2556_ = new_n2551_ & new_n2554_;
  assign n1484 = ~new_n2555_ | ~new_n2556_;
  assign new_n2558_ = n_n137 & new_n1157_;
  assign new_n2559_ = pkey_165_ & new_n1136_;
  assign new_n2560_ = n_n2448 & new_n1161_;
  assign new_n2561_ = n_n140 & new_n1164_1_;
  assign new_n2562_ = ~new_n2560_ & ~new_n2561_;
  assign new_n2563_ = n_n138 & new_n1168_;
  assign new_n2564_ = pkey_157_ & new_n1170_;
  assign new_n2565_ = ~new_n2563_ & ~new_n2564_;
  assign new_n2566_ = ~new_n2558_ & ~new_n2559_;
  assign new_n2567_ = new_n2562_ & new_n2565_;
  assign n1489 = ~new_n2566_ | ~new_n2567_;
  assign new_n2569_ = n_n144 & new_n1157_;
  assign new_n2570_ = pkey_174_ & new_n1136_;
  assign new_n2571_ = n_n148 & new_n1161_;
  assign new_n2572_ = n_n147 & new_n1164_1_;
  assign new_n2573_ = ~new_n2571_ & ~new_n2572_;
  assign new_n2574_ = n_n145 & new_n1168_;
  assign new_n2575_ = pkey_166_ & new_n1170_;
  assign new_n2576_ = ~new_n2574_ & ~new_n2575_;
  assign new_n2577_ = ~new_n2569_ & ~new_n2570_;
  assign new_n2578_ = new_n2573_ & new_n2576_;
  assign n1494 = ~new_n2577_ | ~new_n2578_;
  assign new_n2580_ = n_n152 & new_n1157_;
  assign new_n2581_ = pkey_84_ & new_n1136_;
  assign new_n2582_ = n_n156 & new_n1161_;
  assign new_n2583_ = n_n155 & new_n1164_1_;
  assign new_n2584_ = ~new_n2582_ & ~new_n2583_;
  assign new_n2585_ = n_n153 & new_n1168_;
  assign new_n2586_ = pkey_76_ & new_n1170_;
  assign new_n2587_ = ~new_n2585_ & ~new_n2586_;
  assign new_n2588_ = ~new_n2580_ & ~new_n2581_;
  assign new_n2589_ = new_n2584_ & new_n2587_;
  assign n1499 = ~new_n2588_ | ~new_n2589_;
  assign new_n2591_ = n_n2474 & new_n1157_;
  assign new_n2592_ = pkey_93_ & new_n1136_;
  assign new_n2593_ = n_n163 & new_n1161_;
  assign new_n2594_ = n_n162 & new_n1164_1_;
  assign new_n2595_ = ~new_n2593_ & ~new_n2594_;
  assign new_n2596_ = n_n2476 & new_n1168_;
  assign new_n2597_ = pkey_85_ & new_n1170_;
  assign new_n2598_ = ~new_n2596_ & ~new_n2597_;
  assign new_n2599_ = ~new_n2591_ & ~new_n2592_;
  assign new_n2600_ = new_n2595_ & new_n2598_;
  assign n1504 = ~new_n2599_ | ~new_n2600_;
  assign new_n2602_ = n_n166 & new_n1157_;
  assign new_n2603_ = pkey_102_ & new_n1136_;
  assign new_n2604_ = n_n170 & new_n1161_;
  assign new_n2605_ = n_n169 & new_n1164_1_;
  assign new_n2606_ = ~new_n2604_ & ~new_n2605_;
  assign new_n2607_ = n_n167 & new_n1168_;
  assign new_n2608_ = pkey_94_ & new_n1170_;
  assign new_n2609_ = ~new_n2607_ & ~new_n2608_;
  assign new_n2610_ = ~new_n2602_ & ~new_n2603_;
  assign new_n2611_ = new_n2606_ & new_n2609_;
  assign n1509 = ~new_n2610_ | ~new_n2611_;
  assign new_n2613_ = n_n2517 & new_n1157_;
  assign new_n2614_ = pkey_30_ & new_n1136_;
  assign new_n2615_ = n_n193 & new_n1161_;
  assign new_n2616_ = n_n192 & new_n1164_1_;
  assign new_n2617_ = ~new_n2615_ & ~new_n2616_;
  assign new_n2618_ = n_n190 & new_n1168_;
  assign new_n2619_ = pkey_22_ & new_n1170_;
  assign new_n2620_ = ~new_n2618_ & ~new_n2619_;
  assign new_n2621_ = ~new_n2613_ & ~new_n2614_;
  assign new_n2622_ = new_n2617_ & new_n2620_;
  assign n1514 = ~new_n2621_ | ~new_n2622_;
  assign new_n2624_ = n_n47 & new_n1157_;
  assign new_n2625_ = pkey_144_ & new_n1136_;
  assign new_n2626_ = n_n51 & new_n1161_;
  assign new_n2627_ = n_n50 & new_n1164_1_;
  assign new_n2628_ = ~new_n2626_ & ~new_n2627_;
  assign new_n2629_ = n_n48 & new_n1168_;
  assign new_n2630_ = pkey_136_ & new_n1170_;
  assign new_n2631_ = ~new_n2629_ & ~new_n2630_;
  assign new_n2632_ = ~new_n2624_ & ~new_n2625_;
  assign new_n2633_ = new_n2628_ & new_n2631_;
  assign n1519 = ~new_n2632_ | ~new_n2633_;
  assign new_n2635_ = n_n2333 & new_n1157_;
  assign new_n2636_ = pkey_74_ & new_n1136_;
  assign new_n2637_ = n_n60 & new_n1161_;
  assign new_n2638_ = n_n2337 & new_n1164_1_;
  assign new_n2639_ = ~new_n2637_ & ~new_n2638_;
  assign new_n2640_ = n_n58 & new_n1168_;
  assign new_n2641_ = pkey_66_ & new_n1170_;
  assign new_n2642_ = ~new_n2640_ & ~new_n2641_;
  assign new_n2643_ = ~new_n2635_ & ~new_n2636_;
  assign new_n2644_ = new_n2639_ & new_n2642_;
  assign n1524 = ~new_n2643_ | ~new_n2644_;
  assign new_n2646_ = n_n66 & new_n1157_;
  assign new_n2647_ = pkey_97_ & new_n1136_;
  assign new_n2648_ = n_n70 & new_n1161_;
  assign new_n2649_ = n_n69 & new_n1164_1_;
  assign new_n2650_ = ~new_n2648_ & ~new_n2649_;
  assign new_n2651_ = n_n67 & new_n1168_;
  assign new_n2652_ = pkey_89_ & new_n1170_;
  assign new_n2653_ = ~new_n2651_ & ~new_n2652_;
  assign new_n2654_ = ~new_n2646_ & ~new_n2647_;
  assign new_n2655_ = new_n2650_ & new_n2653_;
  assign n1529 = ~new_n2654_ | ~new_n2655_;
  assign new_n2657_ = n_n76 & new_n1157_;
  assign new_n2658_ = pkey_120_ & new_n1136_;
  assign new_n2659_ = n_n80 & new_n1161_;
  assign new_n2660_ = n_n79 & new_n1164_1_;
  assign new_n2661_ = ~new_n2659_ & ~new_n2660_;
  assign new_n2662_ = n_n77 & new_n1168_;
  assign new_n2663_ = pkey_112_ & new_n1170_;
  assign new_n2664_ = ~new_n2662_ & ~new_n2663_;
  assign new_n2665_ = ~new_n2657_ & ~new_n2658_;
  assign new_n2666_ = new_n2661_ & new_n2664_;
  assign n1534 = ~new_n2665_ | ~new_n2666_;
  assign new_n2668_ = n_n85 & new_n1157_;
  assign new_n2669_ = pkey_50_ & new_n1136_;
  assign new_n2670_ = n_n88 & new_n1161_;
  assign new_n2671_ = n_n87 & new_n1164_1_;
  assign new_n2672_ = ~new_n2670_ & ~new_n2671_;
  assign new_n2673_ = n_n86 & new_n1168_;
  assign new_n2674_ = pkey_42_ & new_n1170_;
  assign new_n2675_ = ~new_n2673_ & ~new_n2674_;
  assign new_n2676_ = ~new_n2668_ & ~new_n2669_;
  assign new_n2677_ = new_n2672_ & new_n2675_;
  assign n1539 = ~new_n2676_ | ~new_n2677_;
  assign new_n2679_ = n_n48 & new_n1157_;
  assign new_n2680_ = pkey_152_ & new_n1136_;
  assign new_n2681_ = n_n52 & new_n1161_;
  assign new_n2682_ = n_n51 & new_n1164_1_;
  assign new_n2683_ = ~new_n2681_ & ~new_n2682_;
  assign new_n2684_ = n_n49 & new_n1168_;
  assign new_n2685_ = pkey_144_ & new_n1170_;
  assign new_n2686_ = ~new_n2684_ & ~new_n2685_;
  assign new_n2687_ = ~new_n2679_ & ~new_n2680_;
  assign new_n2688_ = new_n2683_ & new_n2686_;
  assign n1544 = ~new_n2687_ | ~new_n2688_;
  assign new_n2690_ = n_n57 & new_n1157_;
  assign new_n2691_ = pkey_66_ & new_n1136_;
  assign new_n2692_ = n_n2337 & new_n1161_;
  assign new_n2693_ = n_n59 & new_n1164_1_;
  assign new_n2694_ = ~new_n2692_ & ~new_n2693_;
  assign new_n2695_ = n_n2333 & new_n1168_;
  assign new_n2696_ = pkey_123_ & new_n1170_;
  assign new_n2697_ = ~new_n2695_ & ~new_n2696_;
  assign new_n2698_ = ~new_n2690_ & ~new_n2691_;
  assign new_n2699_ = new_n2694_ & new_n2697_;
  assign n1549 = ~new_n2698_ | ~new_n2699_;
  assign new_n2701_ = n_n67 & new_n1157_;
  assign new_n2702_ = pkey_105_ & new_n1136_;
  assign new_n2703_ = n_n2352 & new_n1161_;
  assign new_n2704_ = n_n70 & new_n1164_1_;
  assign new_n2705_ = ~new_n2703_ & ~new_n2704_;
  assign new_n2706_ = n_n68 & new_n1168_;
  assign new_n2707_ = pkey_97_ & new_n1170_;
  assign new_n2708_ = ~new_n2706_ & ~new_n2707_;
  assign new_n2709_ = ~new_n2701_ & ~new_n2702_;
  assign new_n2710_ = new_n2705_ & new_n2708_;
  assign n1554 = ~new_n2709_ | ~new_n2710_;
  assign new_n2712_ = n_n75 & new_n1157_;
  assign new_n2713_ = pkey_112_ & new_n1136_;
  assign new_n2714_ = n_n79 & new_n1161_;
  assign new_n2715_ = n_n78 & new_n1164_1_;
  assign new_n2716_ = ~new_n2714_ & ~new_n2715_;
  assign new_n2717_ = n_n76 & new_n1168_;
  assign new_n2718_ = pkey_104_ & new_n1170_;
  assign new_n2719_ = ~new_n2717_ & ~new_n2718_;
  assign new_n2720_ = ~new_n2712_ & ~new_n2713_;
  assign new_n2721_ = new_n2716_ & new_n2719_;
  assign n1559 = ~new_n2720_ | ~new_n2721_;
  assign new_n2723_ = n_n86 & new_n1157_;
  assign new_n2724_ = pkey_58_ & new_n1136_;
  assign new_n2725_ = n_n89 & new_n1161_;
  assign new_n2726_ = n_n88 & new_n1164_1_;
  assign new_n2727_ = ~new_n2725_ & ~new_n2726_;
  assign new_n2728_ = n_n2374 & new_n1168_;
  assign new_n2729_ = pkey_50_ & new_n1170_;
  assign new_n2730_ = ~new_n2728_ & ~new_n2729_;
  assign new_n2731_ = ~new_n2723_ & ~new_n2724_;
  assign new_n2732_ = new_n2727_ & new_n2730_;
  assign n1564 = ~new_n2731_ | ~new_n2732_;
  assign new_n2734_ = n_n49 & new_n1157_;
  assign new_n2735_ = pkey_160_ & new_n1136_;
  assign new_n2736_ = n_n53 & new_n1161_;
  assign new_n2737_ = n_n52 & new_n1164_1_;
  assign new_n2738_ = ~new_n2736_ & ~new_n2737_;
  assign new_n2739_ = n_n50 & new_n1168_;
  assign new_n2740_ = pkey_152_ & new_n1170_;
  assign new_n2741_ = ~new_n2739_ & ~new_n2740_;
  assign new_n2742_ = ~new_n2734_ & ~new_n2735_;
  assign new_n2743_ = new_n2738_ & new_n2741_;
  assign n1569 = ~new_n2742_ | ~new_n2743_;
  assign new_n2745_ = n_n59 & new_n1157_;
  assign new_n2746_ = pkey_90_ & new_n1136_;
  assign new_n2747_ = n_n62 & new_n1161_;
  assign new_n2748_ = n_n61 & new_n1164_1_;
  assign new_n2749_ = ~new_n2747_ & ~new_n2748_;
  assign new_n2750_ = n_n2337 & new_n1168_;
  assign new_n2751_ = pkey_82_ & new_n1170_;
  assign new_n2752_ = ~new_n2750_ & ~new_n2751_;
  assign new_n2753_ = ~new_n2745_ & ~new_n2746_;
  assign new_n2754_ = new_n2749_ & new_n2752_;
  assign n1574 = ~new_n2753_ | ~new_n2754_;
  assign new_n2756_ = n_n64 & new_n1157_;
  assign new_n2757_ = pkey_81_ & new_n1136_;
  assign new_n2758_ = n_n68 & new_n1161_;
  assign new_n2759_ = n_n67 & new_n1164_1_;
  assign new_n2760_ = ~new_n2758_ & ~new_n2759_;
  assign new_n2761_ = n_n65 & new_n1168_;
  assign new_n2762_ = pkey_73_ & new_n1170_;
  assign new_n2763_ = ~new_n2761_ & ~new_n2762_;
  assign new_n2764_ = ~new_n2756_ & ~new_n2757_;
  assign new_n2765_ = new_n2760_ & new_n2763_;
  assign n1579 = ~new_n2764_ | ~new_n2765_;
  assign new_n2767_ = n_n74 & new_n1157_;
  assign new_n2768_ = pkey_104_ & new_n1136_;
  assign new_n2769_ = n_n78 & new_n1161_;
  assign new_n2770_ = n_n77 & new_n1164_1_;
  assign new_n2771_ = ~new_n2769_ & ~new_n2770_;
  assign new_n2772_ = n_n75 & new_n1168_;
  assign new_n2773_ = pkey_96_ & new_n1170_;
  assign new_n2774_ = ~new_n2772_ & ~new_n2773_;
  assign new_n2775_ = ~new_n2767_ & ~new_n2768_;
  assign new_n2776_ = new_n2771_ & new_n2774_;
  assign n1584 = ~new_n2775_ | ~new_n2776_;
  assign new_n2778_ = n_n2374 & new_n1157_;
  assign new_n2779_ = pkey_1_ & new_n1136_;
  assign new_n2780_ = n_n90 & new_n1161_;
  assign new_n2781_ = n_n89 & new_n1164_1_;
  assign new_n2782_ = ~new_n2780_ & ~new_n2781_;
  assign new_n2783_ = n_n87 & new_n1168_;
  assign new_n2784_ = pkey_58_ & new_n1170_;
  assign new_n2785_ = ~new_n2783_ & ~new_n2784_;
  assign new_n2786_ = ~new_n2778_ & ~new_n2779_;
  assign new_n2787_ = new_n2782_ & new_n2785_;
  assign n1589 = ~new_n2786_ | ~new_n2787_;
  assign new_n2789_ = n_n101 & new_n1157_;
  assign new_n2790_ = pkey_227_ & new_n1136_;
  assign new_n2791_ = n_n10 & new_n1161_;
  assign new_n2792_ = n_n9 & new_n1164_1_;
  assign new_n2793_ = ~new_n2791_ & ~new_n2792_;
  assign new_n2794_ = n_n102 & new_n1168_;
  assign new_n2795_ = pkey_56_ & new_n1170_;
  assign new_n2796_ = ~new_n2794_ & ~new_n2795_;
  assign new_n2797_ = ~new_n2789_ & ~new_n2790_;
  assign new_n2798_ = new_n2793_ & new_n2796_;
  assign n1594 = ~new_n2797_ | ~new_n2798_;
  assign new_n2800_ = n_n50 & new_n1157_;
  assign new_n2801_ = pkey_168_ & new_n1136_;
  assign new_n2802_ = n_n54 & new_n1161_;
  assign new_n2803_ = n_n53 & new_n1164_1_;
  assign new_n2804_ = ~new_n2802_ & ~new_n2803_;
  assign new_n2805_ = n_n51 & new_n1168_;
  assign new_n2806_ = pkey_160_ & new_n1170_;
  assign new_n2807_ = ~new_n2805_ & ~new_n2806_;
  assign new_n2808_ = ~new_n2800_ & ~new_n2801_;
  assign new_n2809_ = new_n2804_ & new_n2807_;
  assign n1599 = ~new_n2808_ | ~new_n2809_;
  assign new_n2811_ = n_n58 & new_n1157_;
  assign new_n2812_ = pkey_82_ & new_n1136_;
  assign new_n2813_ = n_n61 & new_n1161_;
  assign new_n2814_ = n_n60 & new_n1164_1_;
  assign new_n2815_ = ~new_n2813_ & ~new_n2814_;
  assign new_n2816_ = n_n59 & new_n1168_;
  assign new_n2817_ = pkey_74_ & new_n1170_;
  assign new_n2818_ = ~new_n2816_ & ~new_n2817_;
  assign new_n2819_ = ~new_n2811_ & ~new_n2812_;
  assign new_n2820_ = new_n2815_ & new_n2818_;
  assign n1604 = ~new_n2819_ | ~new_n2820_;
  assign new_n2822_ = n_n65 & new_n1157_;
  assign new_n2823_ = pkey_89_ & new_n1136_;
  assign new_n2824_ = n_n69 & new_n1161_;
  assign new_n2825_ = n_n68 & new_n1164_1_;
  assign new_n2826_ = ~new_n2824_ & ~new_n2825_;
  assign new_n2827_ = n_n66 & new_n1168_;
  assign new_n2828_ = pkey_81_ & new_n1170_;
  assign new_n2829_ = ~new_n2827_ & ~new_n2828_;
  assign new_n2830_ = ~new_n2822_ & ~new_n2823_;
  assign new_n2831_ = new_n2826_ & new_n2829_;
  assign n1609 = ~new_n2830_ | ~new_n2831_;
  assign new_n2833_ = n_n73 & new_n1157_;
  assign new_n2834_ = pkey_96_ & new_n1136_;
  assign new_n2835_ = n_n77 & new_n1161_;
  assign new_n2836_ = n_n76 & new_n1164_1_;
  assign new_n2837_ = ~new_n2835_ & ~new_n2836_;
  assign new_n2838_ = n_n74 & new_n1168_;
  assign new_n2839_ = pkey_88_ & new_n1170_;
  assign new_n2840_ = ~new_n2838_ & ~new_n2839_;
  assign new_n2841_ = ~new_n2833_ & ~new_n2834_;
  assign new_n2842_ = new_n2837_ & new_n2840_;
  assign n1614 = ~new_n2841_ | ~new_n2842_;
  assign new_n2844_ = n_n87 & new_n1157_;
  assign new_n2845_ = pkey_9_ & new_n1136_;
  assign new_n2846_ = n_n91 & new_n1161_;
  assign new_n2847_ = n_n90 & new_n1164_1_;
  assign new_n2848_ = ~new_n2846_ & ~new_n2847_;
  assign new_n2849_ = n_n88 & new_n1168_;
  assign new_n2850_ = pkey_1_ & new_n1170_;
  assign new_n2851_ = ~new_n2849_ & ~new_n2850_;
  assign new_n2852_ = ~new_n2844_ & ~new_n2845_;
  assign new_n2853_ = new_n2848_ & new_n2851_;
  assign n1619 = ~new_n2852_ | ~new_n2853_;
  assign new_n2855_ = n_n14 & new_n1157_;
  assign new_n2856_ = pkey_242_ & new_n1136_;
  assign new_n2857_ = n_n2280 & new_n1161_;
  assign new_n2858_ = n_n16 & new_n1164_1_;
  assign new_n2859_ = ~new_n2857_ & ~new_n2858_;
  assign new_n2860_ = n_n15 & new_n1168_;
  assign new_n2861_ = pkey_234_ & new_n1170_;
  assign new_n2862_ = ~new_n2860_ & ~new_n2861_;
  assign new_n2863_ = ~new_n2855_ & ~new_n2856_;
  assign new_n2864_ = new_n2859_ & new_n2862_;
  assign n1624 = ~new_n2863_ | ~new_n2864_;
  assign new_n2866_ = n_n2288 & new_n1157_;
  assign new_n2867_ = pkey_200_ & new_n1136_;
  assign new_n2868_ = n_n26 & new_n1161_;
  assign new_n2869_ = n_n25 & new_n1164_1_;
  assign new_n2870_ = ~new_n2868_ & ~new_n2869_;
  assign new_n2871_ = n_n23 & new_n1168_;
  assign new_n2872_ = pkey_192_ & new_n1170_;
  assign new_n2873_ = ~new_n2871_ & ~new_n2872_;
  assign new_n2874_ = ~new_n2866_ & ~new_n2867_;
  assign new_n2875_ = new_n2870_ & new_n2873_;
  assign n1629 = ~new_n2874_ | ~new_n2875_;
  assign new_n2877_ = n_n33 & new_n1157_;
  assign new_n2878_ = pkey_130_ & new_n1136_;
  assign new_n2879_ = n_n2305 & new_n1161_;
  assign new_n2880_ = n_n35 & new_n1164_1_;
  assign new_n2881_ = ~new_n2879_ & ~new_n2880_;
  assign new_n2882_ = n_n2301 & new_n1168_;
  assign new_n2883_ = pkey_187_ & new_n1170_;
  assign new_n2884_ = ~new_n2882_ & ~new_n2883_;
  assign new_n2885_ = ~new_n2877_ & ~new_n2878_;
  assign new_n2886_ = new_n2881_ & new_n2884_;
  assign n1634 = ~new_n2885_ | ~new_n2886_;
  assign new_n2888_ = n_n41 & new_n1157_;
  assign new_n2889_ = pkey_153_ & new_n1136_;
  assign new_n2890_ = n_n45 & new_n1161_;
  assign new_n2891_ = n_n44 & new_n1164_1_;
  assign new_n2892_ = ~new_n2890_ & ~new_n2891_;
  assign new_n2893_ = n_n42 & new_n1168_;
  assign new_n2894_ = pkey_145_ & new_n1170_;
  assign new_n2895_ = ~new_n2893_ & ~new_n2894_;
  assign new_n2896_ = ~new_n2888_ & ~new_n2889_;
  assign new_n2897_ = new_n2892_ & new_n2895_;
  assign n1639 = ~new_n2896_ | ~new_n2897_;
  assign new_n2899_ = n_n88 & new_n1157_;
  assign new_n2900_ = pkey_17_ & new_n1136_;
  assign new_n2901_ = n_n92 & new_n1161_;
  assign new_n2902_ = n_n91 & new_n1164_1_;
  assign new_n2903_ = ~new_n2901_ & ~new_n2902_;
  assign new_n2904_ = n_n89 & new_n1168_;
  assign new_n2905_ = pkey_9_ & new_n1170_;
  assign new_n2906_ = ~new_n2904_ & ~new_n2905_;
  assign new_n2907_ = ~new_n2899_ & ~new_n2900_;
  assign new_n2908_ = new_n2903_ & new_n2906_;
  assign n1644 = ~new_n2907_ | ~new_n2908_;
  assign new_n2910_ = n_n15 & new_n1157_;
  assign new_n2911_ = pkey_250_ & new_n1136_;
  assign new_n2912_ = n_n17 & new_n1161_;
  assign new_n2913_ = n_n2280 & new_n1164_1_;
  assign new_n2914_ = ~new_n2912_ & ~new_n2913_;
  assign new_n2915_ = n_n2277 & new_n1168_;
  assign new_n2916_ = pkey_242_ & new_n1170_;
  assign new_n2917_ = ~new_n2915_ & ~new_n2916_;
  assign new_n2918_ = ~new_n2910_ & ~new_n2911_;
  assign new_n2919_ = new_n2914_ & new_n2917_;
  assign n1649 = ~new_n2918_ | ~new_n2919_;
  assign new_n2921_ = n_n22 & new_n1157_;
  assign new_n2922_ = pkey_192_ & new_n1136_;
  assign new_n2923_ = n_n25 & new_n1161_;
  assign new_n2924_ = n_n24 & new_n1164_1_;
  assign new_n2925_ = ~new_n2923_ & ~new_n2924_;
  assign new_n2926_ = n_n2288 & new_n1168_;
  assign new_n2927_ = pkey_249_ & new_n1170_;
  assign new_n2928_ = ~new_n2926_ & ~new_n2927_;
  assign new_n2929_ = ~new_n2921_ & ~new_n2922_;
  assign new_n2930_ = new_n2925_ & new_n2928_;
  assign n1654 = ~new_n2929_ | ~new_n2930_;
  assign new_n2932_ = n_n2301 & new_n1157_;
  assign new_n2933_ = pkey_138_ & new_n1136_;
  assign new_n2934_ = n_n36 & new_n1161_;
  assign new_n2935_ = n_n2305 & new_n1164_1_;
  assign new_n2936_ = ~new_n2934_ & ~new_n2935_;
  assign new_n2937_ = n_n34 & new_n1168_;
  assign new_n2938_ = pkey_130_ & new_n1170_;
  assign new_n2939_ = ~new_n2937_ & ~new_n2938_;
  assign new_n2940_ = ~new_n2932_ & ~new_n2933_;
  assign new_n2941_ = new_n2936_ & new_n2939_;
  assign n1659 = ~new_n2940_ | ~new_n2941_;
  assign new_n2943_ = n_n40 & new_n1157_;
  assign new_n2944_ = pkey_145_ & new_n1136_;
  assign new_n2945_ = n_n44 & new_n1161_;
  assign new_n2946_ = n_n43 & new_n1164_1_;
  assign new_n2947_ = ~new_n2945_ & ~new_n2946_;
  assign new_n2948_ = n_n41 & new_n1168_;
  assign new_n2949_ = pkey_137_ & new_n1170_;
  assign new_n2950_ = ~new_n2948_ & ~new_n2949_;
  assign new_n2951_ = ~new_n2943_ & ~new_n2944_;
  assign new_n2952_ = new_n2947_ & new_n2950_;
  assign n1664 = ~new_n2951_ | ~new_n2952_;
  assign new_n2954_ = n_n89 & new_n1157_;
  assign new_n2955_ = pkey_25_ & new_n1136_;
  assign new_n2956_ = n_n93 & new_n1161_;
  assign new_n2957_ = n_n92 & new_n1164_1_;
  assign new_n2958_ = ~new_n2956_ & ~new_n2957_;
  assign new_n2959_ = n_n90 & new_n1168_;
  assign new_n2960_ = pkey_17_ & new_n1170_;
  assign new_n2961_ = ~new_n2959_ & ~new_n2960_;
  assign new_n2962_ = ~new_n2954_ & ~new_n2955_;
  assign new_n2963_ = new_n2958_ & new_n2961_;
  assign n1669 = ~new_n2962_ | ~new_n2963_;
  assign new_n2965_ = n_n2277 & new_n1157_;
  assign new_n2966_ = pkey_193_ & new_n1136_;
  assign new_n2967_ = n_n18 & new_n1161_;
  assign new_n2968_ = n_n17 & new_n1164_1_;
  assign new_n2969_ = ~new_n2967_ & ~new_n2968_;
  assign new_n2970_ = n_n16 & new_n1168_;
  assign new_n2971_ = pkey_250_ & new_n1170_;
  assign new_n2972_ = ~new_n2970_ & ~new_n2971_;
  assign new_n2973_ = ~new_n2965_ & ~new_n2966_;
  assign new_n2974_ = new_n2969_ & new_n2972_;
  assign n1674 = ~new_n2973_ | ~new_n2974_;
  assign new_n2976_ = n_n24 & new_n1157_;
  assign new_n2977_ = pkey_216_ & new_n1136_;
  assign new_n2978_ = n_n28 & new_n1161_;
  assign new_n2979_ = n_n27 & new_n1164_1_;
  assign new_n2980_ = ~new_n2978_ & ~new_n2979_;
  assign new_n2981_ = n_n25 & new_n1168_;
  assign new_n2982_ = pkey_208_ & new_n1170_;
  assign new_n2983_ = ~new_n2981_ & ~new_n2982_;
  assign new_n2984_ = ~new_n2976_ & ~new_n2977_;
  assign new_n2985_ = new_n2980_ & new_n2983_;
  assign n1679 = ~new_n2984_ | ~new_n2985_;
  assign new_n2987_ = n_n31 & new_n1157_;
  assign new_n2988_ = pkey_179_ & new_n1136_;
  assign new_n2989_ = n_n34 & new_n1161_;
  assign new_n2990_ = n_n2301 & new_n1164_1_;
  assign new_n2991_ = ~new_n2989_ & ~new_n2990_;
  assign new_n2992_ = n_n32 & new_n1168_;
  assign new_n2993_ = pkey_171_ & new_n1170_;
  assign new_n2994_ = ~new_n2992_ & ~new_n2993_;
  assign new_n2995_ = ~new_n2987_ & ~new_n2988_;
  assign new_n2996_ = new_n2991_ & new_n2994_;
  assign n1684 = ~new_n2995_ | ~new_n2996_;
  assign new_n2998_ = n_n39 & new_n1157_;
  assign new_n2999_ = pkey_137_ & new_n1136_;
  assign new_n3000_ = n_n43 & new_n1161_;
  assign new_n3001_ = n_n42 & new_n1164_1_;
  assign new_n3002_ = ~new_n3000_ & ~new_n3001_;
  assign new_n3003_ = n_n40 & new_n1168_;
  assign new_n3004_ = pkey_129_ & new_n1170_;
  assign new_n3005_ = ~new_n3003_ & ~new_n3004_;
  assign new_n3006_ = ~new_n2998_ & ~new_n2999_;
  assign new_n3007_ = new_n3002_ & new_n3005_;
  assign n1689 = ~new_n3006_ | ~new_n3007_;
  assign new_n3009_ = n_n16 & new_n1157_;
  assign new_n3010_ = pkey_201_ & new_n1136_;
  assign new_n3011_ = n_n19 & new_n1161_;
  assign new_n3012_ = n_n18 & new_n1164_1_;
  assign new_n3013_ = ~new_n3011_ & ~new_n3012_;
  assign new_n3014_ = n_n2280 & new_n1168_;
  assign new_n3015_ = pkey_193_ & new_n1170_;
  assign new_n3016_ = ~new_n3014_ & ~new_n3015_;
  assign new_n3017_ = ~new_n3009_ & ~new_n3010_;
  assign new_n3018_ = new_n3013_ & new_n3016_;
  assign n1694 = ~new_n3017_ | ~new_n3018_;
  assign new_n3020_ = n_n23 & new_n1157_;
  assign new_n3021_ = pkey_208_ & new_n1136_;
  assign new_n3022_ = n_n27 & new_n1161_;
  assign new_n3023_ = n_n26 & new_n1164_1_;
  assign new_n3024_ = ~new_n3022_ & ~new_n3023_;
  assign new_n3025_ = n_n24 & new_n1168_;
  assign new_n3026_ = pkey_200_ & new_n1170_;
  assign new_n3027_ = ~new_n3025_ & ~new_n3026_;
  assign new_n3028_ = ~new_n3020_ & ~new_n3021_;
  assign new_n3029_ = new_n3024_ & new_n3027_;
  assign n1699 = ~new_n3028_ | ~new_n3029_;
  assign new_n3031_ = n_n32 & new_n1157_;
  assign new_n3032_ = pkey_187_ & new_n1136_;
  assign new_n3033_ = n_n35 & new_n1161_;
  assign new_n3034_ = n_n34 & new_n1164_1_;
  assign new_n3035_ = ~new_n3033_ & ~new_n3034_;
  assign new_n3036_ = n_n33 & new_n1168_;
  assign new_n3037_ = pkey_179_ & new_n1170_;
  assign new_n3038_ = ~new_n3036_ & ~new_n3037_;
  assign new_n3039_ = ~new_n3031_ & ~new_n3032_;
  assign new_n3040_ = new_n3035_ & new_n3038_;
  assign n1704 = ~new_n3039_ | ~new_n3040_;
  assign new_n3042_ = n_n2310 & new_n1157_;
  assign new_n3043_ = pkey_129_ & new_n1136_;
  assign new_n3044_ = n_n42 & new_n1161_;
  assign new_n3045_ = n_n41 & new_n1164_1_;
  assign new_n3046_ = ~new_n3044_ & ~new_n3045_;
  assign new_n3047_ = n_n39 & new_n1168_;
  assign new_n3048_ = pkey_186_ & new_n1170_;
  assign new_n3049_ = ~new_n3047_ & ~new_n3048_;
  assign new_n3050_ = ~new_n3042_ & ~new_n3043_;
  assign new_n3051_ = new_n3046_ & new_n3049_;
  assign n1709 = ~new_n3050_ | ~new_n3051_;
  assign new_n3053_ = n_n2280 & new_n1157_;
  assign new_n3054_ = pkey_209_ & new_n1136_;
  assign new_n3055_ = n_n20 & new_n1161_;
  assign new_n3056_ = n_n19 & new_n1164_1_;
  assign new_n3057_ = ~new_n3055_ & ~new_n3056_;
  assign new_n3058_ = n_n17 & new_n1168_;
  assign new_n3059_ = pkey_201_ & new_n1170_;
  assign new_n3060_ = ~new_n3058_ & ~new_n3059_;
  assign new_n3061_ = ~new_n3053_ & ~new_n3054_;
  assign new_n3062_ = new_n3057_ & new_n3060_;
  assign n1714 = ~new_n3061_ | ~new_n3062_;
  assign new_n3064_ = n_n26 & new_n1157_;
  assign new_n3065_ = pkey_232_ & new_n1136_;
  assign new_n3066_ = n_n30 & new_n1161_;
  assign new_n3067_ = n_n29 & new_n1164_1_;
  assign new_n3068_ = ~new_n3066_ & ~new_n3067_;
  assign new_n3069_ = n_n27 & new_n1168_;
  assign new_n3070_ = pkey_224_ & new_n1170_;
  assign new_n3071_ = ~new_n3069_ & ~new_n3070_;
  assign new_n3072_ = ~new_n3064_ & ~new_n3065_;
  assign new_n3073_ = new_n3068_ & new_n3071_;
  assign n1719 = ~new_n3072_ | ~new_n3073_;
  assign new_n3075_ = n_n2305 & new_n1157_;
  assign new_n3076_ = pkey_162_ & new_n1136_;
  assign new_n3077_ = n_n2310 & new_n1161_;
  assign new_n3078_ = n_n38 & new_n1164_1_;
  assign new_n3079_ = ~new_n3077_ & ~new_n3078_;
  assign new_n3080_ = n_n36 & new_n1168_;
  assign new_n3081_ = pkey_154_ & new_n1170_;
  assign new_n3082_ = ~new_n3080_ & ~new_n3081_;
  assign new_n3083_ = ~new_n3075_ & ~new_n3076_;
  assign new_n3084_ = new_n3079_ & new_n3082_;
  assign n1724 = ~new_n3083_ | ~new_n3084_;
  assign new_n3086_ = n_n45 & new_n1157_;
  assign new_n3087_ = pkey_185_ & new_n1136_;
  assign new_n3088_ = n_n48 & new_n1161_;
  assign new_n3089_ = n_n47 & new_n1164_1_;
  assign new_n3090_ = ~new_n3088_ & ~new_n3089_;
  assign new_n3091_ = n_n46 & new_n1168_;
  assign new_n3092_ = pkey_177_ & new_n1170_;
  assign new_n3093_ = ~new_n3091_ & ~new_n3092_;
  assign new_n3094_ = ~new_n3086_ & ~new_n3087_;
  assign new_n3095_ = new_n3090_ & new_n3093_;
  assign n1729 = ~new_n3094_ | ~new_n3095_;
  assign new_n3097_ = n_n55 & new_n1157_;
  assign new_n3098_ = pkey_115_ & new_n1136_;
  assign new_n3099_ = n_n58 & new_n1161_;
  assign new_n3100_ = n_n2333 & new_n1164_1_;
  assign new_n3101_ = ~new_n3099_ & ~new_n3100_;
  assign new_n3102_ = n_n56 & new_n1168_;
  assign new_n3103_ = pkey_107_ & new_n1170_;
  assign new_n3104_ = ~new_n3102_ & ~new_n3103_;
  assign new_n3105_ = ~new_n3097_ & ~new_n3098_;
  assign new_n3106_ = new_n3101_ & new_n3104_;
  assign n1734 = ~new_n3105_ | ~new_n3106_;
  assign new_n3108_ = n_n63 & new_n1157_;
  assign new_n3109_ = pkey_73_ & new_n1136_;
  assign new_n3110_ = n_n67 & new_n1161_;
  assign new_n3111_ = n_n66 & new_n1164_1_;
  assign new_n3112_ = ~new_n3110_ & ~new_n3111_;
  assign new_n3113_ = n_n64 & new_n1168_;
  assign new_n3114_ = pkey_65_ & new_n1170_;
  assign new_n3115_ = ~new_n3113_ & ~new_n3114_;
  assign new_n3116_ = ~new_n3108_ & ~new_n3109_;
  assign new_n3117_ = new_n3112_ & new_n3115_;
  assign n1739 = ~new_n3116_ | ~new_n3117_;
  assign new_n3119_ = n_n17 & new_n1157_;
  assign new_n3120_ = pkey_217_ & new_n1136_;
  assign new_n3121_ = n_n21 & new_n1161_;
  assign new_n3122_ = n_n20 & new_n1164_1_;
  assign new_n3123_ = ~new_n3121_ & ~new_n3122_;
  assign new_n3124_ = n_n18 & new_n1168_;
  assign new_n3125_ = pkey_209_ & new_n1170_;
  assign new_n3126_ = ~new_n3124_ & ~new_n3125_;
  assign new_n3127_ = ~new_n3119_ & ~new_n3120_;
  assign new_n3128_ = new_n3123_ & new_n3126_;
  assign n1744 = ~new_n3127_ | ~new_n3128_;
  assign new_n3130_ = n_n25 & new_n1157_;
  assign new_n3131_ = pkey_224_ & new_n1136_;
  assign new_n3132_ = n_n29 & new_n1161_;
  assign new_n3133_ = n_n28 & new_n1164_1_;
  assign new_n3134_ = ~new_n3132_ & ~new_n3133_;
  assign new_n3135_ = n_n26 & new_n1168_;
  assign new_n3136_ = pkey_216_ & new_n1170_;
  assign new_n3137_ = ~new_n3135_ & ~new_n3136_;
  assign new_n3138_ = ~new_n3130_ & ~new_n3131_;
  assign new_n3139_ = new_n3134_ & new_n3137_;
  assign n1749 = ~new_n3138_ | ~new_n3139_;
  assign new_n3141_ = n_n36 & new_n1157_;
  assign new_n3142_ = pkey_170_ & new_n1136_;
  assign new_n3143_ = n_n39 & new_n1161_;
  assign new_n3144_ = n_n2310 & new_n1164_1_;
  assign new_n3145_ = ~new_n3143_ & ~new_n3144_;
  assign new_n3146_ = n_n37 & new_n1168_;
  assign new_n3147_ = pkey_162_ & new_n1170_;
  assign new_n3148_ = ~new_n3146_ & ~new_n3147_;
  assign new_n3149_ = ~new_n3141_ & ~new_n3142_;
  assign new_n3150_ = new_n3145_ & new_n3148_;
  assign n1754 = ~new_n3149_ | ~new_n3150_;
  assign new_n3152_ = n_n44 & new_n1157_;
  assign new_n3153_ = pkey_177_ & new_n1136_;
  assign new_n3154_ = n_n47 & new_n1161_;
  assign new_n3155_ = n_n2320 & new_n1164_1_;
  assign new_n3156_ = ~new_n3154_ & ~new_n3155_;
  assign new_n3157_ = n_n45 & new_n1168_;
  assign new_n3158_ = pkey_169_ & new_n1170_;
  assign new_n3159_ = ~new_n3157_ & ~new_n3158_;
  assign new_n3160_ = ~new_n3152_ & ~new_n3153_;
  assign new_n3161_ = new_n3156_ & new_n3159_;
  assign n1759 = ~new_n3160_ | ~new_n3161_;
  assign new_n3163_ = n_n56 & new_n1157_;
  assign new_n3164_ = pkey_123_ & new_n1136_;
  assign new_n3165_ = n_n59 & new_n1161_;
  assign new_n3166_ = n_n58 & new_n1164_1_;
  assign new_n3167_ = ~new_n3165_ & ~new_n3166_;
  assign new_n3168_ = n_n57 & new_n1168_;
  assign new_n3169_ = pkey_115_ & new_n1170_;
  assign new_n3170_ = ~new_n3168_ & ~new_n3169_;
  assign new_n3171_ = ~new_n3163_ & ~new_n3164_;
  assign new_n3172_ = new_n3167_ & new_n3170_;
  assign n1764 = ~new_n3171_ | ~new_n3172_;
  assign new_n3174_ = n_n2342 & new_n1157_;
  assign new_n3175_ = pkey_65_ & new_n1136_;
  assign new_n3176_ = n_n66 & new_n1161_;
  assign new_n3177_ = n_n65 & new_n1164_1_;
  assign new_n3178_ = ~new_n3176_ & ~new_n3177_;
  assign new_n3179_ = n_n63 & new_n1168_;
  assign new_n3180_ = pkey_122_ & new_n1170_;
  assign new_n3181_ = ~new_n3179_ & ~new_n3180_;
  assign new_n3182_ = ~new_n3174_ & ~new_n3175_;
  assign new_n3183_ = new_n3178_ & new_n3181_;
  assign n1769 = ~new_n3182_ | ~new_n3183_;
  assign new_n3185_ = n_n18 & new_n1157_;
  assign new_n3186_ = pkey_225_ & new_n1136_;
  assign new_n3187_ = n_n22 & new_n1161_;
  assign new_n3188_ = n_n21 & new_n1164_1_;
  assign new_n3189_ = ~new_n3187_ & ~new_n3188_;
  assign new_n3190_ = n_n19 & new_n1168_;
  assign new_n3191_ = pkey_217_ & new_n1170_;
  assign new_n3192_ = ~new_n3190_ & ~new_n3191_;
  assign new_n3193_ = ~new_n3185_ & ~new_n3186_;
  assign new_n3194_ = new_n3189_ & new_n3192_;
  assign n1774 = ~new_n3193_ | ~new_n3194_;
  assign new_n3196_ = n_n28 & new_n1157_;
  assign new_n3197_ = pkey_248_ & new_n1136_;
  assign new_n3198_ = n_n32 & new_n1161_;
  assign new_n3199_ = n_n31 & new_n1164_1_;
  assign new_n3200_ = ~new_n3198_ & ~new_n3199_;
  assign new_n3201_ = n_n29 & new_n1168_;
  assign new_n3202_ = pkey_240_ & new_n1170_;
  assign new_n3203_ = ~new_n3201_ & ~new_n3202_;
  assign new_n3204_ = ~new_n3196_ & ~new_n3197_;
  assign new_n3205_ = new_n3200_ & new_n3203_;
  assign n1779 = ~new_n3204_ | ~new_n3205_;
  assign new_n3207_ = n_n34 & new_n1157_;
  assign new_n3208_ = pkey_146_ & new_n1136_;
  assign new_n3209_ = n_n37 & new_n1161_;
  assign new_n3210_ = n_n36 & new_n1164_1_;
  assign new_n3211_ = ~new_n3209_ & ~new_n3210_;
  assign new_n3212_ = n_n35 & new_n1168_;
  assign new_n3213_ = pkey_138_ & new_n1170_;
  assign new_n3214_ = ~new_n3212_ & ~new_n3213_;
  assign new_n3215_ = ~new_n3207_ & ~new_n3208_;
  assign new_n3216_ = new_n3211_ & new_n3214_;
  assign n1784 = ~new_n3215_ | ~new_n3216_;
  assign new_n3218_ = n_n43 & new_n1157_;
  assign new_n3219_ = pkey_169_ & new_n1136_;
  assign new_n3220_ = n_n2320 & new_n1161_;
  assign new_n3221_ = n_n46 & new_n1164_1_;
  assign new_n3222_ = ~new_n3220_ & ~new_n3221_;
  assign new_n3223_ = n_n44 & new_n1168_;
  assign new_n3224_ = pkey_161_ & new_n1170_;
  assign new_n3225_ = ~new_n3223_ & ~new_n3224_;
  assign new_n3226_ = ~new_n3218_ & ~new_n3219_;
  assign new_n3227_ = new_n3222_ & new_n3225_;
  assign n1789 = ~new_n3226_ | ~new_n3227_;
  assign new_n3229_ = n_n71 & new_n1157_;
  assign new_n3230_ = pkey_80_ & new_n1136_;
  assign new_n3231_ = n_n75 & new_n1161_;
  assign new_n3232_ = n_n74 & new_n1164_1_;
  assign new_n3233_ = ~new_n3231_ & ~new_n3232_;
  assign new_n3234_ = n_n72 & new_n1168_;
  assign new_n3235_ = pkey_72_ & new_n1170_;
  assign new_n3236_ = ~new_n3234_ & ~new_n3235_;
  assign new_n3237_ = ~new_n3229_ & ~new_n3230_;
  assign new_n3238_ = new_n3233_ & new_n3236_;
  assign n1794 = ~new_n3237_ | ~new_n3238_;
  assign new_n3240_ = n_n2365 & new_n1157_;
  assign new_n3241_ = pkey_10_ & new_n1136_;
  assign new_n3242_ = n_n84 & new_n1161_;
  assign new_n3243_ = n_n2369 & new_n1164_1_;
  assign new_n3244_ = ~new_n3242_ & ~new_n3243_;
  assign new_n3245_ = n_n82 & new_n1168_;
  assign new_n3246_ = pkey_2_ & new_n1170_;
  assign new_n3247_ = ~new_n3245_ & ~new_n3246_;
  assign new_n3248_ = ~new_n3240_ & ~new_n3241_;
  assign new_n3249_ = new_n3244_ & new_n3247_;
  assign n1799 = ~new_n3248_ | ~new_n3249_;
  assign new_n3251_ = n_n19 & new_n1157_;
  assign new_n3252_ = pkey_233_ & new_n1136_;
  assign new_n3253_ = n_n2288 & new_n1161_;
  assign new_n3254_ = n_n22 & new_n1164_1_;
  assign new_n3255_ = ~new_n3253_ & ~new_n3254_;
  assign new_n3256_ = n_n20 & new_n1168_;
  assign new_n3257_ = pkey_225_ & new_n1170_;
  assign new_n3258_ = ~new_n3256_ & ~new_n3257_;
  assign new_n3259_ = ~new_n3251_ & ~new_n3252_;
  assign new_n3260_ = new_n3255_ & new_n3258_;
  assign n1804 = ~new_n3259_ | ~new_n3260_;
  assign new_n3262_ = n_n27 & new_n1157_;
  assign new_n3263_ = pkey_240_ & new_n1136_;
  assign new_n3264_ = n_n31 & new_n1161_;
  assign new_n3265_ = n_n30 & new_n1164_1_;
  assign new_n3266_ = ~new_n3264_ & ~new_n3265_;
  assign new_n3267_ = n_n28 & new_n1168_;
  assign new_n3268_ = pkey_232_ & new_n1170_;
  assign new_n3269_ = ~new_n3267_ & ~new_n3268_;
  assign new_n3270_ = ~new_n3262_ & ~new_n3263_;
  assign new_n3271_ = new_n3266_ & new_n3269_;
  assign n1809 = ~new_n3270_ | ~new_n3271_;
  assign new_n3273_ = n_n35 & new_n1157_;
  assign new_n3274_ = pkey_154_ & new_n1136_;
  assign new_n3275_ = n_n38 & new_n1161_;
  assign new_n3276_ = n_n37 & new_n1164_1_;
  assign new_n3277_ = ~new_n3275_ & ~new_n3276_;
  assign new_n3278_ = n_n2305 & new_n1168_;
  assign new_n3279_ = pkey_146_ & new_n1170_;
  assign new_n3280_ = ~new_n3278_ & ~new_n3279_;
  assign new_n3281_ = ~new_n3273_ & ~new_n3274_;
  assign new_n3282_ = new_n3277_ & new_n3280_;
  assign n1814 = ~new_n3281_ | ~new_n3282_;
  assign new_n3284_ = n_n42 & new_n1157_;
  assign new_n3285_ = pkey_161_ & new_n1136_;
  assign new_n3286_ = n_n46 & new_n1161_;
  assign new_n3287_ = n_n45 & new_n1164_1_;
  assign new_n3288_ = ~new_n3286_ & ~new_n3287_;
  assign new_n3289_ = n_n43 & new_n1168_;
  assign new_n3290_ = pkey_153_ & new_n1170_;
  assign new_n3291_ = ~new_n3289_ & ~new_n3290_;
  assign new_n3292_ = ~new_n3284_ & ~new_n3285_;
  assign new_n3293_ = new_n3288_ & new_n3291_;
  assign n1819 = ~new_n3292_ | ~new_n3293_;
  assign new_n3295_ = n_n72 & new_n1157_;
  assign new_n3296_ = pkey_88_ & new_n1136_;
  assign new_n3297_ = n_n76 & new_n1161_;
  assign new_n3298_ = n_n75 & new_n1164_1_;
  assign new_n3299_ = ~new_n3297_ & ~new_n3298_;
  assign new_n3300_ = n_n73 & new_n1168_;
  assign new_n3301_ = pkey_80_ & new_n1170_;
  assign new_n3302_ = ~new_n3300_ & ~new_n3301_;
  assign new_n3303_ = ~new_n3295_ & ~new_n3296_;
  assign new_n3304_ = new_n3299_ & new_n3302_;
  assign n1824 = ~new_n3303_ | ~new_n3304_;
  assign new_n3306_ = n_n81 & new_n1157_;
  assign new_n3307_ = pkey_2_ & new_n1136_;
  assign new_n3308_ = n_n2369 & new_n1161_;
  assign new_n3309_ = n_n83 & new_n1164_1_;
  assign new_n3310_ = ~new_n3308_ & ~new_n3309_;
  assign new_n3311_ = n_n2365 & new_n1168_;
  assign new_n3312_ = pkey_59_ & new_n1170_;
  assign new_n3313_ = ~new_n3311_ & ~new_n3312_;
  assign new_n3314_ = ~new_n3306_ & ~new_n3307_;
  assign new_n3315_ = new_n3310_ & new_n3313_;
  assign n1829 = ~new_n3314_ | ~new_n3315_;
  assign new_n3317_ = n_n20 & new_n1157_;
  assign new_n3318_ = pkey_241_ & new_n1136_;
  assign new_n3319_ = n_n23 & new_n1161_;
  assign new_n3320_ = n_n2288 & new_n1164_1_;
  assign new_n3321_ = ~new_n3319_ & ~new_n3320_;
  assign new_n3322_ = n_n21 & new_n1168_;
  assign new_n3323_ = pkey_233_ & new_n1170_;
  assign new_n3324_ = ~new_n3322_ & ~new_n3323_;
  assign new_n3325_ = ~new_n3317_ & ~new_n3318_;
  assign new_n3326_ = new_n3321_ & new_n3324_;
  assign n1834 = ~new_n3325_ | ~new_n3326_;
  assign new_n3328_ = n_n30 & new_n1157_;
  assign new_n3329_ = pkey_171_ & new_n1136_;
  assign new_n3330_ = n_n2301 & new_n1161_;
  assign new_n3331_ = n_n33 & new_n1164_1_;
  assign new_n3332_ = ~new_n3330_ & ~new_n3331_;
  assign new_n3333_ = n_n31 & new_n1168_;
  assign new_n3334_ = pkey_163_ & new_n1170_;
  assign new_n3335_ = ~new_n3333_ & ~new_n3334_;
  assign new_n3336_ = ~new_n3328_ & ~new_n3329_;
  assign new_n3337_ = new_n3332_ & new_n3335_;
  assign n1839 = ~new_n3336_ | ~new_n3337_;
  assign new_n3339_ = n_n51 & new_n1157_;
  assign new_n3340_ = pkey_176_ & new_n1136_;
  assign new_n3341_ = n_n55 & new_n1161_;
  assign new_n3342_ = n_n54 & new_n1164_1_;
  assign new_n3343_ = ~new_n3341_ & ~new_n3342_;
  assign new_n3344_ = n_n52 & new_n1168_;
  assign new_n3345_ = pkey_168_ & new_n1170_;
  assign new_n3346_ = ~new_n3344_ & ~new_n3345_;
  assign new_n3347_ = ~new_n3339_ & ~new_n3340_;
  assign new_n3348_ = new_n3343_ & new_n3346_;
  assign n1844 = ~new_n3347_ | ~new_n3348_;
  assign new_n3350_ = n_n60 & new_n1157_;
  assign new_n3351_ = pkey_106_ & new_n1136_;
  assign new_n3352_ = n_n63 & new_n1161_;
  assign new_n3353_ = n_n2342 & new_n1164_1_;
  assign new_n3354_ = ~new_n3352_ & ~new_n3353_;
  assign new_n3355_ = n_n61 & new_n1168_;
  assign new_n3356_ = pkey_98_ & new_n1170_;
  assign new_n3357_ = ~new_n3355_ & ~new_n3356_;
  assign new_n3358_ = ~new_n3350_ & ~new_n3351_;
  assign new_n3359_ = new_n3354_ & new_n3357_;
  assign n1849 = ~new_n3358_ | ~new_n3359_;
  assign new_n3361_ = n_n70 & new_n1157_;
  assign new_n3362_ = pkey_64_ & new_n1136_;
  assign new_n3363_ = n_n73 & new_n1161_;
  assign new_n3364_ = n_n72 & new_n1164_1_;
  assign new_n3365_ = ~new_n3363_ & ~new_n3364_;
  assign new_n3366_ = n_n2352 & new_n1168_;
  assign new_n3367_ = pkey_121_ & new_n1170_;
  assign new_n3368_ = ~new_n3366_ & ~new_n3367_;
  assign new_n3369_ = ~new_n3361_ & ~new_n3362_;
  assign new_n3370_ = new_n3365_ & new_n3368_;
  assign n1854 = ~new_n3369_ | ~new_n3370_;
  assign new_n3372_ = n_n80 & new_n1157_;
  assign new_n3373_ = pkey_59_ & new_n1136_;
  assign new_n3374_ = n_n83 & new_n1161_;
  assign new_n3375_ = n_n82 & new_n1164_1_;
  assign new_n3376_ = ~new_n3374_ & ~new_n3375_;
  assign new_n3377_ = n_n81 & new_n1168_;
  assign new_n3378_ = pkey_51_ & new_n1170_;
  assign new_n3379_ = ~new_n3377_ & ~new_n3378_;
  assign new_n3380_ = ~new_n3372_ & ~new_n3373_;
  assign new_n3381_ = new_n3376_ & new_n3379_;
  assign n1859 = ~new_n3380_ | ~new_n3381_;
  assign new_n3383_ = n_n82 & new_n1157_;
  assign new_n3384_ = pkey_18_ & new_n1136_;
  assign new_n3385_ = n_n85 & new_n1161_;
  assign new_n3386_ = n_n84 & new_n1164_1_;
  assign new_n3387_ = ~new_n3385_ & ~new_n3386_;
  assign new_n3388_ = n_n83 & new_n1168_;
  assign new_n3389_ = pkey_10_ & new_n1170_;
  assign new_n3390_ = ~new_n3388_ & ~new_n3389_;
  assign new_n3391_ = ~new_n3383_ & ~new_n3384_;
  assign new_n3392_ = new_n3387_ & new_n3390_;
  assign n1864 = ~new_n3391_ | ~new_n3392_;
  assign new_n3394_ = n_n21 & new_n1157_;
  assign new_n3395_ = pkey_249_ & new_n1136_;
  assign new_n3396_ = n_n24 & new_n1161_;
  assign new_n3397_ = n_n23 & new_n1164_1_;
  assign new_n3398_ = ~new_n3396_ & ~new_n3397_;
  assign new_n3399_ = n_n22 & new_n1168_;
  assign new_n3400_ = pkey_241_ & new_n1170_;
  assign new_n3401_ = ~new_n3399_ & ~new_n3400_;
  assign new_n3402_ = ~new_n3394_ & ~new_n3395_;
  assign new_n3403_ = new_n3398_ & new_n3401_;
  assign n1869 = ~new_n3402_ | ~new_n3403_;
  assign new_n3405_ = n_n29 & new_n1157_;
  assign new_n3406_ = pkey_163_ & new_n1136_;
  assign new_n3407_ = n_n33 & new_n1161_;
  assign new_n3408_ = n_n32 & new_n1164_1_;
  assign new_n3409_ = ~new_n3407_ & ~new_n3408_;
  assign new_n3410_ = n_n30 & new_n1168_;
  assign new_n3411_ = pkey_248_ & new_n1170_;
  assign new_n3412_ = ~new_n3410_ & ~new_n3411_;
  assign new_n3413_ = ~new_n3405_ & ~new_n3406_;
  assign new_n3414_ = new_n3409_ & new_n3412_;
  assign n1874 = ~new_n3413_ | ~new_n3414_;
  assign new_n3416_ = n_n52 & new_n1157_;
  assign new_n3417_ = pkey_184_ & new_n1136_;
  assign new_n3418_ = n_n56 & new_n1161_;
  assign new_n3419_ = n_n55 & new_n1164_1_;
  assign new_n3420_ = ~new_n3418_ & ~new_n3419_;
  assign new_n3421_ = n_n53 & new_n1168_;
  assign new_n3422_ = pkey_176_ & new_n1170_;
  assign new_n3423_ = ~new_n3421_ & ~new_n3422_;
  assign new_n3424_ = ~new_n3416_ & ~new_n3417_;
  assign new_n3425_ = new_n3420_ & new_n3423_;
  assign n1879 = ~new_n3424_ | ~new_n3425_;
  assign new_n3427_ = n_n2337 & new_n1157_;
  assign new_n3428_ = pkey_98_ & new_n1136_;
  assign new_n3429_ = n_n2342 & new_n1161_;
  assign new_n3430_ = n_n62 & new_n1164_1_;
  assign new_n3431_ = ~new_n3429_ & ~new_n3430_;
  assign new_n3432_ = n_n60 & new_n1168_;
  assign new_n3433_ = pkey_90_ & new_n1170_;
  assign new_n3434_ = ~new_n3432_ & ~new_n3433_;
  assign new_n3435_ = ~new_n3427_ & ~new_n3428_;
  assign new_n3436_ = new_n3431_ & new_n3434_;
  assign n1884 = ~new_n3435_ | ~new_n3436_;
  assign new_n3438_ = n_n2352 & new_n1157_;
  assign new_n3439_ = pkey_72_ & new_n1136_;
  assign new_n3440_ = n_n74 & new_n1161_;
  assign new_n3441_ = n_n73 & new_n1164_1_;
  assign new_n3442_ = ~new_n3440_ & ~new_n3441_;
  assign new_n3443_ = n_n71 & new_n1168_;
  assign new_n3444_ = pkey_64_ & new_n1170_;
  assign new_n3445_ = ~new_n3443_ & ~new_n3444_;
  assign new_n3446_ = ~new_n3438_ & ~new_n3439_;
  assign new_n3447_ = new_n3442_ & new_n3445_;
  assign n1889 = ~new_n3446_ | ~new_n3447_;
  assign new_n3449_ = n_n79 & new_n1157_;
  assign new_n3450_ = pkey_51_ & new_n1136_;
  assign new_n3451_ = n_n82 & new_n1161_;
  assign new_n3452_ = n_n2365 & new_n1164_1_;
  assign new_n3453_ = ~new_n3451_ & ~new_n3452_;
  assign new_n3454_ = n_n80 & new_n1168_;
  assign new_n3455_ = pkey_43_ & new_n1170_;
  assign new_n3456_ = ~new_n3454_ & ~new_n3455_;
  assign new_n3457_ = ~new_n3449_ & ~new_n3450_;
  assign new_n3458_ = new_n3453_ & new_n3456_;
  assign n1894 = ~new_n3457_ | ~new_n3458_;
  assign new_n3460_ = n_n83 & new_n1157_;
  assign new_n3461_ = pkey_26_ & new_n1136_;
  assign new_n3462_ = n_n86 & new_n1161_;
  assign new_n3463_ = n_n85 & new_n1164_1_;
  assign new_n3464_ = ~new_n3462_ & ~new_n3463_;
  assign new_n3465_ = n_n2369 & new_n1168_;
  assign new_n3466_ = pkey_18_ & new_n1170_;
  assign new_n3467_ = ~new_n3465_ & ~new_n3466_;
  assign new_n3468_ = ~new_n3460_ & ~new_n3461_;
  assign new_n3469_ = new_n3464_ & new_n3467_;
  assign n1899 = ~new_n3468_ | ~new_n3469_;
  assign new_n3471_ = n_n37 & new_n1157_;
  assign new_n3472_ = pkey_178_ & new_n1136_;
  assign new_n3473_ = n_n40 & new_n1161_;
  assign new_n3474_ = n_n39 & new_n1164_1_;
  assign new_n3475_ = ~new_n3473_ & ~new_n3474_;
  assign new_n3476_ = n_n38 & new_n1168_;
  assign new_n3477_ = pkey_170_ & new_n1170_;
  assign new_n3478_ = ~new_n3476_ & ~new_n3477_;
  assign new_n3479_ = ~new_n3471_ & ~new_n3472_;
  assign new_n3480_ = new_n3475_ & new_n3478_;
  assign n1904 = ~new_n3479_ | ~new_n3480_;
  assign new_n3482_ = n_n2320 & new_n1157_;
  assign new_n3483_ = pkey_136_ & new_n1136_;
  assign new_n3484_ = n_n50 & new_n1161_;
  assign new_n3485_ = n_n49 & new_n1164_1_;
  assign new_n3486_ = ~new_n3484_ & ~new_n3485_;
  assign new_n3487_ = n_n47 & new_n1168_;
  assign new_n3488_ = pkey_128_ & new_n1170_;
  assign new_n3489_ = ~new_n3487_ & ~new_n3488_;
  assign new_n3490_ = ~new_n3482_ & ~new_n3483_;
  assign new_n3491_ = new_n3486_ & new_n3489_;
  assign n1909 = ~new_n3490_ | ~new_n3491_;
  assign new_n3493_ = n_n53 & new_n1157_;
  assign new_n3494_ = pkey_99_ & new_n1136_;
  assign new_n3495_ = n_n57 & new_n1161_;
  assign new_n3496_ = n_n56 & new_n1164_1_;
  assign new_n3497_ = ~new_n3495_ & ~new_n3496_;
  assign new_n3498_ = n_n54 & new_n1168_;
  assign new_n3499_ = pkey_184_ & new_n1170_;
  assign new_n3500_ = ~new_n3498_ & ~new_n3499_;
  assign new_n3501_ = ~new_n3493_ & ~new_n3494_;
  assign new_n3502_ = new_n3497_ & new_n3500_;
  assign n1914 = ~new_n3501_ | ~new_n3502_;
  assign new_n3504_ = n_n62 & new_n1157_;
  assign new_n3505_ = pkey_122_ & new_n1136_;
  assign new_n3506_ = n_n65 & new_n1161_;
  assign new_n3507_ = n_n64 & new_n1164_1_;
  assign new_n3508_ = ~new_n3506_ & ~new_n3507_;
  assign new_n3509_ = n_n2342 & new_n1168_;
  assign new_n3510_ = pkey_114_ & new_n1170_;
  assign new_n3511_ = ~new_n3509_ & ~new_n3510_;
  assign new_n3512_ = ~new_n3504_ & ~new_n3505_;
  assign new_n3513_ = new_n3508_ & new_n3511_;
  assign n1919 = ~new_n3512_ | ~new_n3513_;
  assign new_n3515_ = n_n68 & new_n1157_;
  assign new_n3516_ = pkey_113_ & new_n1136_;
  assign new_n3517_ = n_n71 & new_n1161_;
  assign new_n3518_ = n_n2352 & new_n1164_1_;
  assign new_n3519_ = ~new_n3517_ & ~new_n3518_;
  assign new_n3520_ = n_n69 & new_n1168_;
  assign new_n3521_ = pkey_105_ & new_n1170_;
  assign new_n3522_ = ~new_n3520_ & ~new_n3521_;
  assign new_n3523_ = ~new_n3515_ & ~new_n3516_;
  assign new_n3524_ = new_n3519_ & new_n3522_;
  assign n1924 = ~new_n3523_ | ~new_n3524_;
  assign new_n3526_ = n_n78 & new_n1157_;
  assign new_n3527_ = pkey_43_ & new_n1136_;
  assign new_n3528_ = n_n2365 & new_n1161_;
  assign new_n3529_ = n_n81 & new_n1164_1_;
  assign new_n3530_ = ~new_n3528_ & ~new_n3529_;
  assign new_n3531_ = n_n79 & new_n1168_;
  assign new_n3532_ = pkey_35_ & new_n1170_;
  assign new_n3533_ = ~new_n3531_ & ~new_n3532_;
  assign new_n3534_ = ~new_n3526_ & ~new_n3527_;
  assign new_n3535_ = new_n3530_ & new_n3533_;
  assign n1929 = ~new_n3534_ | ~new_n3535_;
  assign new_n3537_ = n_n2369 & new_n1157_;
  assign new_n3538_ = pkey_34_ & new_n1136_;
  assign new_n3539_ = n_n2374 & new_n1161_;
  assign new_n3540_ = n_n86 & new_n1164_1_;
  assign new_n3541_ = ~new_n3539_ & ~new_n3540_;
  assign new_n3542_ = n_n84 & new_n1168_;
  assign new_n3543_ = pkey_26_ & new_n1170_;
  assign new_n3544_ = ~new_n3542_ & ~new_n3543_;
  assign new_n3545_ = ~new_n3537_ & ~new_n3538_;
  assign new_n3546_ = new_n3541_ & new_n3544_;
  assign n1934 = ~new_n3545_ | ~new_n3546_;
  assign new_n3548_ = n_n38 & new_n1157_;
  assign new_n3549_ = pkey_186_ & new_n1136_;
  assign new_n3550_ = n_n41 & new_n1161_;
  assign new_n3551_ = n_n40 & new_n1164_1_;
  assign new_n3552_ = ~new_n3550_ & ~new_n3551_;
  assign new_n3553_ = n_n2310 & new_n1168_;
  assign new_n3554_ = pkey_178_ & new_n1170_;
  assign new_n3555_ = ~new_n3553_ & ~new_n3554_;
  assign new_n3556_ = ~new_n3548_ & ~new_n3549_;
  assign new_n3557_ = new_n3552_ & new_n3555_;
  assign n1939 = ~new_n3556_ | ~new_n3557_;
  assign new_n3559_ = n_n46 & new_n1157_;
  assign new_n3560_ = pkey_128_ & new_n1136_;
  assign new_n3561_ = n_n49 & new_n1161_;
  assign new_n3562_ = n_n48 & new_n1164_1_;
  assign new_n3563_ = ~new_n3561_ & ~new_n3562_;
  assign new_n3564_ = n_n2320 & new_n1168_;
  assign new_n3565_ = pkey_185_ & new_n1170_;
  assign new_n3566_ = ~new_n3564_ & ~new_n3565_;
  assign new_n3567_ = ~new_n3559_ & ~new_n3560_;
  assign new_n3568_ = new_n3563_ & new_n3566_;
  assign n1944 = ~new_n3567_ | ~new_n3568_;
  assign new_n3570_ = n_n54 & new_n1157_;
  assign new_n3571_ = pkey_107_ & new_n1136_;
  assign new_n3572_ = n_n2333 & new_n1161_;
  assign new_n3573_ = n_n57 & new_n1164_1_;
  assign new_n3574_ = ~new_n3572_ & ~new_n3573_;
  assign new_n3575_ = n_n55 & new_n1168_;
  assign new_n3576_ = pkey_99_ & new_n1170_;
  assign new_n3577_ = ~new_n3575_ & ~new_n3576_;
  assign new_n3578_ = ~new_n3570_ & ~new_n3571_;
  assign new_n3579_ = new_n3574_ & new_n3577_;
  assign n1949 = ~new_n3578_ | ~new_n3579_;
  assign new_n3581_ = n_n61 & new_n1157_;
  assign new_n3582_ = pkey_114_ & new_n1136_;
  assign new_n3583_ = n_n64 & new_n1161_;
  assign new_n3584_ = n_n63 & new_n1164_1_;
  assign new_n3585_ = ~new_n3583_ & ~new_n3584_;
  assign new_n3586_ = n_n62 & new_n1168_;
  assign new_n3587_ = pkey_106_ & new_n1170_;
  assign new_n3588_ = ~new_n3586_ & ~new_n3587_;
  assign new_n3589_ = ~new_n3581_ & ~new_n3582_;
  assign new_n3590_ = new_n3585_ & new_n3588_;
  assign n1954 = ~new_n3589_ | ~new_n3590_;
  assign new_n3592_ = n_n69 & new_n1157_;
  assign new_n3593_ = pkey_121_ & new_n1136_;
  assign new_n3594_ = n_n72 & new_n1161_;
  assign new_n3595_ = n_n71 & new_n1164_1_;
  assign new_n3596_ = ~new_n3594_ & ~new_n3595_;
  assign new_n3597_ = n_n70 & new_n1168_;
  assign new_n3598_ = pkey_113_ & new_n1170_;
  assign new_n3599_ = ~new_n3597_ & ~new_n3598_;
  assign new_n3600_ = ~new_n3592_ & ~new_n3593_;
  assign new_n3601_ = new_n3596_ & new_n3599_;
  assign n1959 = ~new_n3600_ | ~new_n3601_;
  assign new_n3603_ = n_n77 & new_n1157_;
  assign new_n3604_ = pkey_35_ & new_n1136_;
  assign new_n3605_ = n_n81 & new_n1161_;
  assign new_n3606_ = n_n80 & new_n1164_1_;
  assign new_n3607_ = ~new_n3605_ & ~new_n3606_;
  assign new_n3608_ = n_n78 & new_n1168_;
  assign new_n3609_ = pkey_120_ & new_n1170_;
  assign new_n3610_ = ~new_n3608_ & ~new_n3609_;
  assign new_n3611_ = ~new_n3603_ & ~new_n3604_;
  assign new_n3612_ = new_n3607_ & new_n3610_;
  assign n1964 = ~new_n3611_ | ~new_n3612_;
  assign new_n3614_ = n_n84 & new_n1157_;
  assign new_n3615_ = pkey_42_ & new_n1136_;
  assign new_n3616_ = n_n87 & new_n1161_;
  assign new_n3617_ = n_n2374 & new_n1164_1_;
  assign new_n3618_ = ~new_n3616_ & ~new_n3617_;
  assign new_n3619_ = n_n85 & new_n1168_;
  assign new_n3620_ = pkey_34_ & new_n1170_;
  assign new_n3621_ = ~new_n3619_ & ~new_n3620_;
  assign new_n3622_ = ~new_n3614_ & ~new_n3615_;
  assign new_n3623_ = new_n3618_ & new_n3621_;
  assign n1969 = ~new_n3622_ | ~new_n3623_;
  assign pksi_50_ = n_n45;
  assign pksi_61_ = n_n38;
  assign pksi_72_ = n_n18;
  assign pksi_83_ = n_n22;
  assign pksi_94_ = n_n19;
  assign pksi_102_ = n_n194;
  assign pksi_115_ = n_n184;
  assign pksi_128_ = n_n153;
  assign pksi_51_ = n_n34;
  assign pksi_60_ = n_n35;
  assign pksi_73_ = n_n16;
  assign pksi_82_ = n_n13;
  assign pksi_95_ = n_n29;
  assign pksi_101_ = n_n173;
  assign pksi_116_ = n_n177;
  assign pksi_127_ = n_n162;
  assign pksi_52_ = n_n54;
  assign pksi_63_ = n_n51;
  assign pksi_70_ = n_n43;
  assign pksi_81_ = n_n25;
  assign pksi_96_ = n_n185;
  assign pksi_100_ = n_n180;
  assign pksi_113_ = n_n174;
  assign pksi_53_ = n_n50;
  assign pksi_62_ = n_n44;
  assign pksi_71_ = n_n53;
  assign pksi_80_ = n_n17;
  assign pksi_97_ = n_n175;
  assign pksi_114_ = n_n181;
  assign pksi_129_ = n_n159;
  assign pksi_54_ = n_n52;
  assign pksi_65_ = n_n47;
  assign pksi_76_ = n_n30;
  assign pksi_87_ = n_n27;
  assign pksi_90_ = n_n10;
  assign pksi_119_ = n_n192;
  assign pksi_124_ = n_n157;
  assign pksi_191_ = n_n121;
  assign pksi_55_ = n_n31;
  assign pksi_64_ = n_n33;
  assign pksi_77_ = n_n26;
  assign pksi_86_ = n_n20;
  assign pksi_91_ = n_n24;
  assign pksi_123_ = n_n164;
  assign pksi_56_ = n_n41;
  assign pksi_67_ = n_n48;
  assign pksi_74_ = n_n21;
  assign pksi_85_ = n_n15;
  assign pksi_92_ = n_n9;
  assign pksi_117_ = n_n189;
  assign pksi_126_ = n_n170;
  assign pksi_57_ = n_n49;
  assign pksi_66_ = n_n40;
  assign pksi_75_ = n_n11;
  assign pksi_84_ = n_n12;
  assign pksi_93_ = n_n14;
  assign pksi_118_ = n_n195;
  assign pksi_125_ = n_n150;
  assign pksi_190_ = n_n124;
  assign pksi_14_ = n_n92;
  assign pksi_25_ = n_n63;
  assign pksi_36_ = n_n59;
  assign pksi_47_ = n_n77;
  assign pksi_120_ = n_n161;
  assign pksi_15_ = n_n99;
  assign pksi_24_ = n_n66;
  assign pksi_37_ = n_n62;
  assign pksi_46_ = n_n67;
  assign pksi_109_ = n_n178;
  assign pksi_16_ = n_n81;
  assign pksi_27_ = n_n58;
  assign pksi_34_ = n_n60;
  assign pksi_45_ = n_n61;
  assign pksi_108_ = n_n183;
  assign pksi_122_ = n_n169;
  assign pksi_17_ = n_n95;
  assign pksi_26_ = n_n69;
  assign pksi_35_ = n_n70;
  assign pksi_44_ = n_n56;
  assign pksi_107_ = n_n179;
  assign pksi_121_ = n_n152;
  assign pksi_10_ = n_n84;
  assign pksi_21_ = n_n85;
  assign pksi_32_ = n_n65;
  assign pksi_43_ = n_n72;
  assign pksi_106_ = n_n191;
  assign pksi_111_ = n_n172;
  assign pksi_11_ = n_n94;
  assign pksi_20_ = n_n80;
  assign pksi_33_ = n_n73;
  assign pksi_42_ = n_n64;
  assign pksi_105_ = n_n182;
  assign pksi_112_ = n_n190;
  assign pksi_12_ = n_n83;
  assign pksi_23_ = n_n101;
  assign pksi_30_ = n_n76;
  assign pksi_41_ = n_n71;
  assign pksi_104_ = n_n176;
  assign pksi_13_ = n_n86;
  assign pksi_22_ = n_n91;
  assign pksi_31_ = n_n55;
  assign pksi_40_ = n_n57;
  assign pksi_103_ = n_n186;
  assign pksi_110_ = n_n187;
  assign pksi_3_ = n_n82;
  assign pksi_151_ = n_n139;
  assign pksi_164_ = n_n130;
  assign pksi_177_ = n_n113;
  assign pksi_2_ = n_n93;
  assign pksi_152_ = n_n129;
  assign pksi_163_ = n_n137;
  assign pksi_178_ = n_n120;
  assign pksi_189_ = n_n118;
  assign pksi_1_ = n_n87;
  assign pksi_166_ = n_n148;
  assign pksi_179_ = n_n110;
  assign pksi_188_ = n_n108;
  assign pksi_0_ = n_n90;
  assign pksi_150_ = n_n147;
  assign pksi_165_ = n_n142;
  assign pksi_187_ = n_n121;
  assign pksi_18_ = n_n88;
  assign pksi_29_ = n_n74;
  assign pksi_142_ = n_n171;
  assign pksi_168_ = n_n109;
  assign pksi_173_ = n_n104;
  assign pksi_186_ = n_n112;
  assign pksi_19_ = n_n96;
  assign pksi_28_ = n_n78;
  assign pksi_130_ = n_n167;
  assign pksi_141_ = n_n165;
  assign pksi_167_ = n_n145;
  assign pksi_174_ = n_n123;
  assign pksi_185_ = n_n105;
  assign pksi_38_ = n_n68;
  assign pksi_49_ = n_n39;
  assign pksi_131_ = n_n156;
  assign pksi_140_ = n_n154;
  assign pksi_175_ = n_n115;
  assign pksi_184_ = n_n119;
  assign pksi_39_ = n_n75;
  assign pksi_48_ = n_n42;
  assign pksi_132_ = n_n160;
  assign pksi_169_ = n_n106;
  assign pksi_176_ = n_n107;
  assign pksi_183_ = n_n103;
  assign pksi_58_ = n_n36;
  assign pksi_69_ = n_n37;
  assign pksi_133_ = n_n155;
  assign pksi_146_ = n_n146;
  assign pksi_159_ = n_n125;
  assign pksi_182_ = n_n116;
  assign pksi_59_ = n_n46;
  assign pksi_68_ = n_n32;
  assign pksi_134_ = n_n163;
  assign pksi_145_ = n_n128;
  assign pksi_170_ = n_n122;
  assign pksi_181_ = n_n109;
  assign pksi_9_ = n_n97;
  assign pksi_78_ = n_n28;
  assign pksi_89_ = n_n23;
  assign pksi_135_ = n_n149;
  assign pksi_144_ = n_n138;
  assign pksi_157_ = n_n131;
  assign pksi_171_ = n_n117;
  assign pksi_180_ = n_n114;
  assign pksi_8_ = n_n89;
  assign pksi_79_ = n_n8;
  assign pksi_88_ = n_n10;
  assign pksi_136_ = n_n166;
  assign pksi_143_ = n_n168;
  assign pksi_158_ = n_n140;
  assign pksi_172_ = n_n111;
  assign pksi_7_ = n_n79;
  assign pksi_98_ = n_n193;
  assign pksi_137_ = n_n151;
  assign pksi_155_ = n_n132;
  assign pksi_160_ = n_n143;
  assign pksi_6_ = n_n100;
  assign pksi_99_ = n_n188;
  assign pksi_138_ = n_n158;
  assign pksi_149_ = n_n126;
  assign pksi_156_ = n_n135;
  assign pksi_5_ = n_n98;
  assign pksi_139_ = n_n168;
  assign pksi_148_ = n_n133;
  assign pksi_153_ = n_n136;
  assign pksi_162_ = n_n134;
  assign pksi_4_ = n_n102;
  assign pksi_147_ = n_n141;
  assign pksi_154_ = n_n144;
  assign pksi_161_ = n_n127;
  always @ (posedge clock) begin
    n_n95 <= n854;
    n_n105 <= n859;
    n_n2410 <= n864;
    n_n122 <= n869;
    n_n132 <= n874;
    n_n141 <= n879;
    n_n178 <= n884;
    n_n2513 <= n889;
    n_n96 <= n894;
    n_n2396 <= n899;
    n_n2412 <= n904;
    n_n121 <= n909;
    n_n133 <= n914;
    n_n2448 <= n919;
    n_n179 <= n924;
    n_n187 <= n929;
    n_n97 <= n934;
    n_n107 <= n939;
    n_n114 <= n944;
    n_n120 <= n949;
    n_n149 <= n954;
    n_n159 <= n959;
    n_n180 <= n964;
    n_n189 <= n969;
    n_n195 <= n974;
    n_n98 <= n979;
    n_n106 <= n984;
    n_n2408 <= n989;
    n_n119 <= n994;
    n_n150 <= n999;
    n_n158 <= n1004;
    n_n181 <= n1009;
    n_n188 <= n1014;
    n_n15 <= n1019;
    n_n92 <= n1024;
    n_n102 <= n1029;
    n_n112 <= n1034;
    n_n2420 <= n1039;
    n_n165 <= n1044;
    n_n174 <= n1049;
    n_n184 <= n1054;
    n_n193 <= n1059;
    n_n93 <= n1064;
    n_n101 <= n1069;
    n_n113 <= n1074;
    n_n118 <= n1079;
    n_n2485 <= n1084;
    n_n2495 <= n1089;
    n_n175 <= n1094;
    n_n194 <= n1099;
    n_n94 <= n1104;
    n_n104 <= n1109;
    n_n110 <= n1114;
    n_n117 <= n1119;
    n_n176 <= n1124;
    n_n186 <= n1129;
    n_n2384 <= n1134;
    n_n103 <= n1139;
    n_n111 <= n1144;
    n_n2416 <= n1149;
    n_n177 <= n1154;
    n_n185 <= n1159;
    n_n192 <= n1164;
    n_n12 <= n1169;
    n_n125 <= n1174;
    n_n2440 <= n1179;
    n_n143 <= n1184;
    n_n153 <= n1189;
    n_n162 <= n1194;
    n_n171 <= n1199;
    n_n2272 <= n1204;
    n_n126 <= n1209;
    n_n134 <= n1214;
    n_n144 <= n1219;
    n_n152 <= n1224;
    n_n163 <= n1229;
    n_n170 <= n1234;
    n_n13 <= n1239;
    n_n2430 <= n1244;
    n_n136 <= n1249;
    n_n142 <= n1254;
    n_n151 <= n1259;
    n_n2481 <= n1264;
    n_n173 <= n1269;
    n_n14 <= n1274;
    n_n127 <= n1279;
    n_n135 <= n1284;
    n_n2452 <= n1289;
    n_n2462 <= n1294;
    n_n164 <= n1299;
    n_n172 <= n1304;
    n_n9 <= n1309;
    n_n99 <= n1314;
    n_n109 <= n1319;
    n_n128 <= n1324;
    n_n138 <= n1329;
    n_n147 <= n1334;
    n_n157 <= n1339;
    n_n160 <= n1344;
    n_n167 <= n1349;
    n_n182 <= n1354;
    n_n190 <= n1359;
    n_n10 <= n1364;
    n_n100 <= n1369;
    n_n108 <= n1374;
    n_n129 <= n1379;
    n_n137 <= n1384;
    n_n148 <= n1389;
    n_n156 <= n1394;
    n_n2474 <= n1399;
    n_n166 <= n1404;
    n_n183 <= n1409;
    n_n2517 <= n1414;
    n_n2268 <= n1419;
    n_n115 <= n1424;
    n_n124 <= n1429;
    n_n130 <= n1434;
    n_n140 <= n1439;
    n_n145 <= n1444;
    n_n155 <= n1449;
    n_n2476 <= n1454;
    n_n169 <= n1459;
    n_n2507 <= n1464;
    n_n11 <= n1469;
    n_n116 <= n1474;
    n_n123 <= n1479;
    n_n131 <= n1484;
    n_n139 <= n1489;
    n_n146 <= n1494;
    n_n154 <= n1499;
    n_n161 <= n1504;
    n_n168 <= n1509;
    n_n191 <= n1514;
    n_n49 <= n1519;
    n_n59 <= n1524;
    n_n68 <= n1529;
    n_n78 <= n1534;
    n_n2374 <= n1539;
    n_n50 <= n1544;
    n_n58 <= n1549;
    n_n69 <= n1554;
    n_n77 <= n1559;
    n_n87 <= n1564;
    n_n51 <= n1569;
    n_n60 <= n1574;
    n_n66 <= n1579;
    n_n76 <= n1584;
    n_n88 <= n1589;
    n_n8 <= n1594;
    n_n52 <= n1599;
    n_n2337 <= n1604;
    n_n67 <= n1609;
    n_n75 <= n1614;
    n_n89 <= n1619;
    n_n2277 <= n1624;
    n_n24 <= n1629;
    n_n34 <= n1634;
    n_n43 <= n1639;
    n_n90 <= n1644;
    n_n16 <= n1649;
    n_n23 <= n1654;
    n_n35 <= n1659;
    n_n42 <= n1664;
    n_n91 <= n1669;
    n_n2280 <= n1674;
    n_n26 <= n1679;
    n_n33 <= n1684;
    n_n41 <= n1689;
    n_n17 <= n1694;
    n_n25 <= n1699;
    n_n2301 <= n1704;
    n_n40 <= n1709;
    n_n18 <= n1714;
    n_n28 <= n1719;
    n_n37 <= n1724;
    n_n2320 <= n1729;
    n_n57 <= n1734;
    n_n65 <= n1739;
    n_n19 <= n1744;
    n_n27 <= n1749;
    n_n38 <= n1754;
    n_n46 <= n1759;
    n_n2333 <= n1764;
    n_n64 <= n1769;
    n_n20 <= n1774;
    n_n30 <= n1779;
    n_n2305 <= n1784;
    n_n45 <= n1789;
    n_n73 <= n1794;
    n_n83 <= n1799;
    n_n21 <= n1804;
    n_n29 <= n1809;
    n_n36 <= n1814;
    n_n44 <= n1819;
    n_n74 <= n1824;
    n_n82 <= n1829;
    n_n22 <= n1834;
    n_n32 <= n1839;
    n_n53 <= n1844;
    n_n62 <= n1849;
    n_n71 <= n1854;
    n_n2365 <= n1859;
    n_n2369 <= n1864;
    n_n2288 <= n1869;
    n_n31 <= n1874;
    n_n54 <= n1879;
    n_n61 <= n1884;
    n_n72 <= n1889;
    n_n81 <= n1894;
    n_n84 <= n1899;
    n_n2310 <= n1904;
    n_n48 <= n1909;
    n_n55 <= n1914;
    n_n63 <= n1919;
    n_n70 <= n1924;
    n_n80 <= n1929;
    n_n85 <= n1934;
    n_n39 <= n1939;
    n_n47 <= n1944;
    n_n56 <= n1949;
    n_n2342 <= n1954;
    n_n2352 <= n1959;
    n_n79 <= n1964;
    n_n86 <= n1969;
  end
endmodule

