module top ( 
    pa1, pb2, pc3, pd4, pe5, pp, pa0, pb3, pc2, pd5, pe4, pq, pa3, pb0,
    pc1, pf4, pg5, pr, pa2, pb1, pc0, pf5, pg4, ps, pa5, pd0, pe1, pf2,
    pg3, pt, pa4, pd1, pe0, pf3, pg2, pu, pb4, pc5, pd2, pe3, pf0, pg1, pv,
    pb5, pc4, pd3, pe2, pf1, pg0, pw, ph0, pi1, pj2, pk3, pl4, pm5, ph1,
    pi0, pj3, pk2, pl5, pm4, py, ph2, pi3, pj0, pk1, pn4, po5, pz, ph3,
    pi2, pj1, pk0, pn5, po4, ph4, pi5, pl0, pm1, pn2, po3, ph5, pi4, pl1,
    pm0, pn3, po2, pj4, pk5, pl2, pm3, pn0, po1, pj5, pk4, pl3, pm2, pn1,
    po0, pp0, pq1, pr2, ps3, pt4, pa, pp1, pq0, pr3, ps2, pu4, pb, pp2,
    pq3, pr0, ps1, pv4, pc, pp3, pq2, pr1, ps0, pw4, pd, pp4, pq5, pt0,
    pu1, pv2, pw3, pe, pp5, pq4, pt1, pu0, pv3, pw2, pf, pr4, pt2, pu3,
    pv0, pw1, pg, pr5, ps4, pt3, pu2, pv1, pw0, ph, px0, py1, pz2, pi, px1,
    py0, pz3, pj, px2, py3, pz0, pk, px3, py2, pz1, pl, px4, pm, py4, pn,
    pz4, po,
    pf6, pg7, ph8, pi9, pq10, pf7, pg6, ph9, pi8, pp10, pd6, pe7, pj8, pk9,
    ps10, pd7, pe6, pj9, pk8, pr10, pb6, pc7, pl8, pm9, pu10, pb7, pc6,
    pl9, pm8, pt10, pa7, pn8, po9, pw10, pa6, pn9, po8, pv10, pa9, pn6,
    po7, py10, pa8, pn7, po6, px10, pb8, pc9, pl6, pm7, pb9, pc8, pl7, pm6,
    pd8, pe9, pj6, pk7, pd9, pe8, pj7, pk6, pf8, pg9, ph6, pi7, pf9, pg8,
    ph7, pi6, pa10, pu5, pv6, pw7, px8, py9, pt5, pv7, pw6, px9, py8, pc10,
    pt6, pu7, pw5, pz8, pb10, pt7, pu6, pv5, pz9, pe10, pr6, ps7, pd10,
    pr7, ps6, pg10, pp6, pq7, ps5, pf10, pp7, pq6, pi10, pp8, pq9, ph10,
    pp9, pq8, pk10, pr8, ps9, pj10, pr9, ps8, pm10, pt8, pu9, py5, pz6,
    pl10, pt9, pu8, px5, pz7, po10, pv8, pw9, px6, py7, pn10, pv9, pw8,
    px7, py6, pz5  );
  input  pa1, pb2, pc3, pd4, pe5, pp, pa0, pb3, pc2, pd5, pe4, pq, pa3,
    pb0, pc1, pf4, pg5, pr, pa2, pb1, pc0, pf5, pg4, ps, pa5, pd0, pe1,
    pf2, pg3, pt, pa4, pd1, pe0, pf3, pg2, pu, pb4, pc5, pd2, pe3, pf0,
    pg1, pv, pb5, pc4, pd3, pe2, pf1, pg0, pw, ph0, pi1, pj2, pk3, pl4,
    pm5, ph1, pi0, pj3, pk2, pl5, pm4, py, ph2, pi3, pj0, pk1, pn4, po5,
    pz, ph3, pi2, pj1, pk0, pn5, po4, ph4, pi5, pl0, pm1, pn2, po3, ph5,
    pi4, pl1, pm0, pn3, po2, pj4, pk5, pl2, pm3, pn0, po1, pj5, pk4, pl3,
    pm2, pn1, po0, pp0, pq1, pr2, ps3, pt4, pa, pp1, pq0, pr3, ps2, pu4,
    pb, pp2, pq3, pr0, ps1, pv4, pc, pp3, pq2, pr1, ps0, pw4, pd, pp4, pq5,
    pt0, pu1, pv2, pw3, pe, pp5, pq4, pt1, pu0, pv3, pw2, pf, pr4, pt2,
    pu3, pv0, pw1, pg, pr5, ps4, pt3, pu2, pv1, pw0, ph, px0, py1, pz2, pi,
    px1, py0, pz3, pj, px2, py3, pz0, pk, px3, py2, pz1, pl, px4, pm, py4,
    pn, pz4, po;
  output pf6, pg7, ph8, pi9, pq10, pf7, pg6, ph9, pi8, pp10, pd6, pe7, pj8,
    pk9, ps10, pd7, pe6, pj9, pk8, pr10, pb6, pc7, pl8, pm9, pu10, pb7,
    pc6, pl9, pm8, pt10, pa7, pn8, po9, pw10, pa6, pn9, po8, pv10, pa9,
    pn6, po7, py10, pa8, pn7, po6, px10, pb8, pc9, pl6, pm7, pb9, pc8, pl7,
    pm6, pd8, pe9, pj6, pk7, pd9, pe8, pj7, pk6, pf8, pg9, ph6, pi7, pf9,
    pg8, ph7, pi6, pa10, pu5, pv6, pw7, px8, py9, pt5, pv7, pw6, px9, py8,
    pc10, pt6, pu7, pw5, pz8, pb10, pt7, pu6, pv5, pz9, pe10, pr6, ps7,
    pd10, pr7, ps6, pg10, pp6, pq7, ps5, pf10, pp7, pq6, pi10, pp8, pq9,
    ph10, pp9, pq8, pk10, pr8, ps9, pj10, pr9, ps8, pm10, pt8, pu9, py5,
    pz6, pl10, pt9, pu8, px5, pz7, po10, pv8, pw9, px6, py7, pn10, pv9,
    pw8, px7, py6, pz5;
  wire new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_,
    new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_,
    new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_,
    new_n329_, new_n330_, new_n331_, new_n332_, new_n334_, new_n335_,
    new_n337_, new_n338_, new_n339_, new_n340_, new_n341_, new_n342_,
    new_n343_, new_n344_, new_n345_, new_n346_, new_n347_, new_n348_,
    new_n349_, new_n350_, new_n351_, new_n352_, new_n354_, new_n355_,
    new_n356_, new_n357_, new_n358_, new_n359_, new_n360_, new_n361_,
    new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_,
    new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n373_,
    new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_,
    new_n380_, new_n381_, new_n382_, new_n383_, new_n384_, new_n385_,
    new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_,
    new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_,
    new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_,
    new_n404_, new_n405_, new_n406_, new_n407_, new_n408_, new_n409_,
    new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_,
    new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n422_,
    new_n423_, new_n424_, new_n425_, new_n426_, new_n427_, new_n428_,
    new_n429_, new_n430_, new_n431_, new_n432_, new_n433_, new_n434_,
    new_n435_, new_n436_, new_n437_, new_n438_, new_n439_, new_n440_,
    new_n441_, new_n442_, new_n443_, new_n444_, new_n445_, new_n446_,
    new_n447_, new_n448_, new_n449_, new_n450_, new_n451_, new_n452_,
    new_n453_, new_n454_, new_n455_, new_n456_, new_n457_, new_n458_,
    new_n459_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_,
    new_n465_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_,
    new_n471_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_,
    new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_,
    new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_,
    new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_,
    new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_,
    new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_,
    new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_,
    new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_,
    new_n528_, new_n529_, new_n530_, new_n531_, new_n532_, new_n533_,
    new_n534_, new_n535_, new_n536_, new_n537_, new_n538_, new_n539_,
    new_n540_, new_n541_, new_n542_, new_n543_, new_n544_, new_n545_,
    new_n546_, new_n547_, new_n548_, new_n549_, new_n550_, new_n551_,
    new_n552_, new_n553_, new_n554_, new_n555_, new_n556_, new_n557_,
    new_n558_, new_n559_, new_n561_, new_n562_, new_n563_, new_n564_,
    new_n565_, new_n566_, new_n567_, new_n568_, new_n570_, new_n571_,
    new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_,
    new_n591_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n732_, new_n733_, new_n734_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n783_, new_n784_,
    new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n812_, new_n813_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n847_, new_n848_, new_n850_,
    new_n851_, new_n853_, new_n854_, new_n855_, new_n857_, new_n858_,
    new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_,
    new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n876_,
    new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_,
    new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n896_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_,
    new_n959_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_,
    new_n965_, new_n966_, new_n967_, new_n969_, new_n970_, new_n971_,
    new_n972_, new_n973_, new_n974_, new_n975_, new_n976_, new_n977_,
    new_n978_, new_n979_, new_n980_, new_n981_, new_n982_, new_n983_,
    new_n984_, new_n985_, new_n986_, new_n987_, new_n988_, new_n990_,
    new_n991_, new_n992_, new_n993_, new_n994_, new_n995_, new_n996_,
    new_n997_, new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_,
    new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_,
    new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1015_, new_n1016_,
    new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_,
    new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_,
    new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_,
    new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_,
    new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_,
    new_n1047_, new_n1048_, new_n1049_, new_n1051_, new_n1052_, new_n1053_,
    new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_,
    new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_,
    new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1072_,
    new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_,
    new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_,
    new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1090_, new_n1091_,
    new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_,
    new_n1099_, new_n1100_, new_n1102_, new_n1103_, new_n1104_, new_n1105_,
    new_n1106_, new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_,
    new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_,
    new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1124_, new_n1125_,
    new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1132_,
    new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_,
    new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1145_,
    new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_,
    new_n1152_, new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_,
    new_n1159_, new_n1160_, new_n1161_, new_n1163_, new_n1164_, new_n1165_,
    new_n1167_, new_n1168_, new_n1169_, new_n1170_, new_n1171_, new_n1172_,
    new_n1173_, new_n1174_, new_n1176_, new_n1177_, new_n1178_, new_n1179_,
    new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1186_,
    new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_,
    new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_,
    new_n1199_, new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_,
    new_n1206_, new_n1207_, new_n1209_, new_n1210_, new_n1212_, new_n1213_,
    new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_, new_n1219_,
    new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_, new_n1225_,
    new_n1227_, new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_,
    new_n1233_, new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1239_,
    new_n1240_, new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_,
    new_n1247_, new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_,
    new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_,
    new_n1260_, new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_,
    new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_,
    new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_,
    new_n1279_, new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_,
    new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_,
    new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_,
    new_n1300_, new_n1301_, new_n1302_, new_n1304_, new_n1305_, new_n1306_,
    new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_, new_n1312_,
    new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_, new_n1318_,
    new_n1320_, new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_,
    new_n1326_, new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_,
    new_n1332_, new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1338_,
    new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1344_, new_n1345_,
    new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_,
    new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1357_, new_n1358_,
    new_n1359_, new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_,
    new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_,
    new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1376_,
    new_n1378_, new_n1379_, new_n1380_, new_n1381_, new_n1382_, new_n1384_,
    new_n1385_, new_n1386_, new_n1387_, new_n1388_, new_n1389_, new_n1390_,
    new_n1391_, new_n1392_, new_n1393_, new_n1395_, new_n1396_, new_n1397_,
    new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_,
    new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_,
    new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_,
    new_n1417_, new_n1418_, new_n1420_, new_n1421_, new_n1422_, new_n1423_,
    new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_, new_n1429_,
    new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_, new_n1436_,
    new_n1437_, new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1442_,
    new_n1443_, new_n1444_, new_n1445_, new_n1446_, new_n1447_, new_n1448_,
    new_n1449_, new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_,
    new_n1455_, new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_,
    new_n1461_, new_n1462_, new_n1463_, new_n1464_, new_n1465_, new_n1466_,
    new_n1467_, new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_,
    new_n1473_, new_n1475_, new_n1476_, new_n1477_, new_n1478_, new_n1479_,
    new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_, new_n1485_,
    new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_, new_n1492_,
    new_n1493_, new_n1494_, new_n1495_, new_n1496_, new_n1497_, new_n1498_,
    new_n1499_, new_n1500_, new_n1502_, new_n1503_, new_n1504_, new_n1505_,
    new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_, new_n1512_,
    new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_, new_n1518_,
    new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_, new_n1524_,
    new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_, new_n1530_,
    new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_, new_n1536_,
    new_n1537_, new_n1538_, new_n1539_, new_n1541_, new_n1542_, new_n1543_,
    new_n1544_, new_n1545_, new_n1546_, new_n1547_, new_n1548_, new_n1550_,
    new_n1551_, new_n1552_, new_n1553_, new_n1554_, new_n1555_, new_n1556_,
    new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1561_, new_n1562_,
    new_n1563_, new_n1564_, new_n1565_, new_n1566_, new_n1567_, new_n1568_,
    new_n1569_, new_n1570_, new_n1571_, new_n1573_, new_n1574_, new_n1575_,
    new_n1576_, new_n1577_, new_n1578_, new_n1579_, new_n1580_, new_n1581_,
    new_n1582_, new_n1583_, new_n1585_, new_n1586_, new_n1587_, new_n1588_,
    new_n1589_, new_n1591_, new_n1592_, new_n1593_, new_n1594_, new_n1595_,
    new_n1596_, new_n1597_, new_n1598_, new_n1600_, new_n1601_, new_n1602_,
    new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_, new_n1608_,
    new_n1609_, new_n1610_, new_n1611_, new_n1613_, new_n1614_, new_n1615_,
    new_n1616_, new_n1617_, new_n1618_, new_n1619_, new_n1620_, new_n1621_,
    new_n1622_, new_n1623_, new_n1624_, new_n1625_, new_n1626_, new_n1627_,
    new_n1628_, new_n1629_, new_n1630_, new_n1631_, new_n1632_, new_n1634_,
    new_n1635_, new_n1636_, new_n1638_, new_n1639_, new_n1640_, new_n1641_,
    new_n1642_, new_n1643_, new_n1645_, new_n1646_, new_n1647_, new_n1648_,
    new_n1649_, new_n1650_, new_n1651_, new_n1652_, new_n1654_, new_n1655_,
    new_n1656_, new_n1657_, new_n1659_, new_n1660_, new_n1661_, new_n1662_,
    new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1668_, new_n1669_,
    new_n1670_, new_n1671_, new_n1672_, new_n1673_, new_n1675_, new_n1676_,
    new_n1678_, new_n1679_, new_n1680_, new_n1681_, new_n1683_, new_n1684_,
    new_n1685_, new_n1686_, new_n1687_, new_n1688_, new_n1689_, new_n1690_,
    new_n1692_, new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_,
    new_n1698_, new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_,
    new_n1704_, new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_,
    new_n1710_, new_n1711_, new_n1713_, new_n1714_, new_n1715_, new_n1716_,
    new_n1717_, new_n1719_, new_n1720_, new_n1721_, new_n1722_, new_n1723_,
    new_n1724_, new_n1725_, new_n1726_, new_n1728_, new_n1729_, new_n1730_,
    new_n1731_, new_n1733_, new_n1734_, new_n1735_, new_n1736_, new_n1737_,
    new_n1738_, new_n1739_, new_n1740_, new_n1742_, new_n1743_, new_n1744_,
    new_n1745_, new_n1746_, new_n1747_, new_n1748_, new_n1749_, new_n1751_,
    new_n1752_, new_n1754_, new_n1755_, new_n1756_, new_n1757_, new_n1758_,
    new_n1759_, new_n1760_, new_n1762_, new_n1763_, new_n1764_, new_n1765_,
    new_n1766_, new_n1768_, new_n1769_, new_n1770_, new_n1772_, new_n1773_,
    new_n1774_, new_n1775_, new_n1776_, new_n1777_, new_n1778_, new_n1779_,
    new_n1781_, new_n1782_, new_n1783_, new_n1784_, new_n1785_, new_n1786_,
    new_n1787_, new_n1788_, new_n1790_, new_n1791_, new_n1792_, new_n1793_,
    new_n1794_, new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1800_,
    new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1805_, new_n1806_,
    new_n1807_, new_n1809_, new_n1810_, new_n1811_, new_n1812_, new_n1813_,
    new_n1814_, new_n1815_, new_n1817_, new_n1818_, new_n1819_, new_n1820_,
    new_n1821_, new_n1822_, new_n1823_, new_n1824_, new_n1825_, new_n1826_,
    new_n1827_, new_n1829_, new_n1830_, new_n1831_, new_n1832_, new_n1833_,
    new_n1834_, new_n1835_, new_n1836_, new_n1838_, new_n1839_, new_n1840_,
    new_n1841_, new_n1842_, new_n1843_, new_n1844_, new_n1845_, new_n1846_,
    new_n1847_, new_n1848_, new_n1849_, new_n1850_, new_n1851_, new_n1852_,
    new_n1853_, new_n1854_, new_n1855_, new_n1856_, new_n1857_, new_n1859_,
    new_n1860_, new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_,
    new_n1866_, new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1873_,
    new_n1874_, new_n1875_, new_n1876_, new_n1877_, new_n1878_, new_n1879_,
    new_n1880_, new_n1882_, new_n1883_, new_n1884_, new_n1885_, new_n1886_,
    new_n1887_, new_n1888_, new_n1889_, new_n1890_, new_n1891_, new_n1892_,
    new_n1893_, new_n1895_, new_n1896_, new_n1897_, new_n1898_, new_n1899_,
    new_n1900_, new_n1901_, new_n1902_, new_n1903_, new_n1904_, new_n1905_,
    new_n1906_, new_n1907_, new_n1908_, new_n1909_, new_n1910_, new_n1911_,
    new_n1912_, new_n1913_, new_n1914_, new_n1916_, new_n1917_, new_n1918_,
    new_n1919_, new_n1920_, new_n1921_, new_n1922_, new_n1923_, new_n1924_,
    new_n1926_, new_n1927_, new_n1928_, new_n1929_, new_n1930_, new_n1931_,
    new_n1932_, new_n1933_, new_n1934_, new_n1935_, new_n1936_, new_n1937_,
    new_n1938_, new_n1939_, new_n1940_, new_n1942_, new_n1943_, new_n1944_,
    new_n1945_, new_n1946_, new_n1947_, new_n1948_, new_n1949_, new_n1951_,
    new_n1952_, new_n1953_, new_n1954_, new_n1955_, new_n1956_, new_n1957_,
    new_n1958_, new_n1959_, new_n1960_, new_n1961_, new_n1962_, new_n1963_,
    new_n1964_, new_n1965_, new_n1966_, new_n1968_, new_n1969_, new_n1970_,
    new_n1971_, new_n1972_, new_n1973_, new_n1974_, new_n1976_, new_n1977_,
    new_n1978_, new_n1979_, new_n1980_, new_n1981_, new_n1982_, new_n1983_,
    new_n1985_, new_n1986_, new_n1987_, new_n1988_, new_n1989_, new_n1990_,
    new_n1991_, new_n1992_, new_n1994_, new_n1995_, new_n1996_, new_n1997_,
    new_n1998_, new_n1999_, new_n2000_, new_n2001_, new_n2002_, new_n2003_,
    new_n2005_, new_n2006_, new_n2007_, new_n2009_, new_n2010_, new_n2011_,
    new_n2012_, new_n2013_, new_n2014_, new_n2015_, new_n2016_, new_n2017_,
    new_n2018_, new_n2019_, new_n2020_, new_n2021_, new_n2022_, new_n2023_,
    new_n2024_, new_n2026_, new_n2027_, new_n2028_, new_n2029_, new_n2030_,
    new_n2031_, new_n2032_, new_n2033_, new_n2034_, new_n2035_, new_n2036_,
    new_n2037_, new_n2038_, new_n2039_, new_n2040_, new_n2041_, new_n2042_,
    new_n2043_, new_n2044_, new_n2045_;
  assign new_n311_ = ~pm1 & ~pb;
  assign new_n312_ = pl1 & pn1;
  assign new_n313_ = new_n311_ & new_n312_;
  assign new_n314_ = ~pn1 & ~pb;
  assign new_n315_ = pm1 & pl1;
  assign new_n316_ = new_n314_ & new_n315_;
  assign new_n317_ = pv0 & new_n316_;
  assign new_n318_ = pr1 & new_n317_;
  assign new_n319_ = ~pj1 & ~po1;
  assign new_n320_ = ~pk1 & po1;
  assign new_n321_ = ~new_n319_ & ~new_n320_;
  assign new_n322_ = pj1 & ~new_n321_;
  assign new_n323_ = pe1 & ~pf1;
  assign new_n324_ = new_n322_ & ~new_n323_;
  assign new_n325_ = ~new_n322_ & new_n323_;
  assign new_n326_ = ~new_n324_ & ~new_n325_;
  assign new_n327_ = ~pi1 & ~ph1;
  assign new_n328_ = new_n322_ & ~new_n326_;
  assign new_n329_ = new_n327_ & new_n328_;
  assign new_n330_ = ~ph1 & ~new_n329_;
  assign new_n331_ = ~pm1 & ~pl1;
  assign new_n332_ = ~pn1 & new_n331_;
  assign pv6 = pb | new_n332_;
  assign new_n334_ = ~new_n326_ & new_n327_;
  assign new_n335_ = new_n323_ & new_n334_;
  assign pn6 = pi1 | new_n335_;
  assign new_n337_ = ~pg1 & ~pn6;
  assign new_n338_ = new_n330_ & pv6;
  assign new_n339_ = new_n337_ & new_n338_;
  assign new_n340_ = ~new_n313_ & ~new_n318_;
  assign new_n341_ = ~pb & ~new_n339_;
  assign new_n342_ = new_n340_ & new_n341_;
  assign new_n343_ = ~pr1 & new_n337_;
  assign new_n344_ = ~new_n316_ & new_n337_;
  assign new_n345_ = ~new_n343_ & ~new_n344_;
  assign new_n346_ = new_n330_ & ~new_n345_;
  assign new_n347_ = pw0 & ~new_n346_;
  assign new_n348_ = px0 & new_n347_;
  assign new_n349_ = pv0 & new_n348_;
  assign new_n350_ = ~py0 & ~new_n349_;
  assign new_n351_ = py0 & new_n349_;
  assign new_n352_ = ~new_n350_ & ~new_n351_;
  assign pf6 = new_n342_ & new_n352_;
  assign new_n354_ = ~px0 & ~py0;
  assign new_n355_ = ~pz0 & new_n354_;
  assign new_n356_ = ~pp1 & ~new_n355_;
  assign new_n357_ = ~pr1 & new_n356_;
  assign new_n358_ = ~pa1 & ~pc1;
  assign new_n359_ = ~pb1 & new_n358_;
  assign new_n360_ = new_n355_ & new_n359_;
  assign new_n361_ = new_n356_ & ~new_n360_;
  assign new_n362_ = ~new_n354_ & ~new_n355_;
  assign new_n363_ = ~pr1 & new_n362_;
  assign new_n364_ = ~new_n360_ & new_n362_;
  assign new_n365_ = ~pv0 & pw0;
  assign new_n366_ = ~pq1 & ~pp1;
  assign new_n367_ = ~pr1 & new_n366_;
  assign new_n368_ = ~new_n360_ & new_n366_;
  assign new_n369_ = ~pq1 & ~new_n354_;
  assign new_n370_ = ~pr1 & new_n369_;
  assign new_n371_ = ~new_n360_ & new_n369_;
  assign new_n372_ = ~new_n370_ & ~new_n371_;
  assign new_n373_ = ~new_n367_ & ~new_n368_;
  assign new_n374_ = new_n372_ & new_n373_;
  assign new_n375_ = ~new_n357_ & ~new_n361_;
  assign new_n376_ = ~new_n363_ & new_n375_;
  assign new_n377_ = ~new_n364_ & new_n365_;
  assign new_n378_ = new_n376_ & new_n377_;
  assign new_n379_ = new_n374_ & new_n378_;
  assign new_n380_ = pv6 & new_n379_;
  assign new_n381_ = ~ph & ~new_n380_;
  assign new_n382_ = ps1 & pt1;
  assign new_n383_ = pu1 & new_n382_;
  assign new_n384_ = ~pk & ~new_n383_;
  assign new_n385_ = pw1 & ~new_n384_;
  assign new_n386_ = pv1 & new_n385_;
  assign new_n387_ = px1 & new_n386_;
  assign new_n388_ = ~pk & ~new_n387_;
  assign new_n389_ = py1 & ~new_n388_;
  assign new_n390_ = ~pi & new_n337_;
  assign new_n391_ = ~new_n389_ & ~new_n390_;
  assign new_n392_ = ~ps1 & ~pt1;
  assign new_n393_ = ~pu1 & new_n392_;
  assign new_n394_ = ~pk & ~new_n393_;
  assign new_n395_ = ~pw1 & ~new_n394_;
  assign new_n396_ = ~pv1 & new_n395_;
  assign new_n397_ = ~px1 & new_n396_;
  assign new_n398_ = ~pk & ~new_n397_;
  assign new_n399_ = ~py1 & ~new_n398_;
  assign new_n400_ = ~new_n389_ & ~new_n399_;
  assign new_n401_ = new_n390_ & ~new_n399_;
  assign new_n402_ = ~new_n391_ & ~new_n400_;
  assign new_n403_ = ~new_n401_ & new_n402_;
  assign new_n404_ = ~new_n381_ & new_n403_;
  assign new_n405_ = ~pz1 & new_n404_;
  assign new_n406_ = pz1 & ~new_n404_;
  assign new_n407_ = ~new_n405_ & ~new_n406_;
  assign new_n408_ = ~pd3 & new_n407_;
  assign new_n409_ = ~pn1 & new_n311_;
  assign new_n410_ = pl1 & new_n409_;
  assign new_n411_ = ~pv6 & ~new_n410_;
  assign new_n412_ = ~pd1 & ~pw0;
  assign new_n413_ = new_n360_ & new_n412_;
  assign new_n414_ = pv0 & new_n413_;
  assign new_n415_ = ~new_n410_ & ~new_n414_;
  assign new_n416_ = ~new_n411_ & ~new_n415_;
  assign new_n417_ = new_n407_ & ~new_n416_;
  assign new_n418_ = ~pd3 & new_n416_;
  assign new_n419_ = ~new_n408_ & ~new_n417_;
  assign new_n420_ = ~new_n418_ & new_n419_;
  assign pg7 = pb | new_n420_;
  assign new_n422_ = pv6 & ~new_n337_;
  assign new_n423_ = ~pg & ~new_n422_;
  assign new_n424_ = pm1 & ~pb;
  assign new_n425_ = ~pn1 & new_n424_;
  assign new_n426_ = ~pl1 & new_n425_;
  assign new_n427_ = ~pb & ~new_n426_;
  assign new_n428_ = ~new_n423_ & ~new_n427_;
  assign new_n429_ = pr1 & ~pv6;
  assign new_n430_ = ~pv0 & new_n429_;
  assign new_n431_ = ~new_n316_ & ~pv6;
  assign new_n432_ = new_n330_ & new_n337_;
  assign new_n433_ = ~pv0 & new_n413_;
  assign new_n434_ = ~new_n432_ & new_n433_;
  assign new_n435_ = pr1 & ~new_n434_;
  assign new_n436_ = ~pv0 & new_n435_;
  assign new_n437_ = ~new_n316_ & ~new_n434_;
  assign new_n438_ = ~new_n430_ & ~new_n431_;
  assign new_n439_ = ~new_n436_ & ~new_n437_;
  assign new_n440_ = new_n438_ & new_n439_;
  assign new_n441_ = ~pf & ~new_n440_;
  assign new_n442_ = pp1 & new_n316_;
  assign new_n443_ = ~pj & new_n442_;
  assign new_n444_ = pr2 & pq2;
  assign new_n445_ = pq1 & new_n316_;
  assign new_n446_ = ~pj & new_n445_;
  assign new_n447_ = ~new_n444_ & ~new_n446_;
  assign new_n448_ = ~new_n443_ & new_n447_;
  assign new_n449_ = ~ps2 & ~new_n443_;
  assign new_n450_ = ~new_n448_ & ~new_n449_;
  assign new_n451_ = pt2 & new_n450_;
  assign new_n452_ = ~pj & ~new_n451_;
  assign new_n453_ = pv2 & ~new_n452_;
  assign new_n454_ = ~new_n423_ & ~new_n453_;
  assign new_n455_ = ~pr2 & ~pq2;
  assign new_n456_ = ~new_n446_ & ~new_n455_;
  assign new_n457_ = ~new_n443_ & new_n456_;
  assign new_n458_ = ps2 & ~new_n443_;
  assign new_n459_ = ~new_n457_ & ~new_n458_;
  assign new_n460_ = ~pt2 & new_n459_;
  assign new_n461_ = ~pj & ~new_n460_;
  assign new_n462_ = pu2 & ~new_n461_;
  assign new_n463_ = ~new_n453_ & ~new_n462_;
  assign new_n464_ = new_n423_ & ~new_n462_;
  assign new_n465_ = ~new_n454_ & ~new_n463_;
  assign new_n466_ = ~new_n464_ & new_n465_;
  assign new_n467_ = ~new_n441_ & new_n466_;
  assign new_n468_ = ~pa3 & new_n467_;
  assign new_n469_ = pa3 & ~new_n467_;
  assign new_n470_ = ~new_n468_ & ~new_n469_;
  assign new_n471_ = new_n427_ & ~new_n470_;
  assign ph8 = new_n428_ | new_n471_;
  assign new_n473_ = ~pm5 & ~pz;
  assign new_n474_ = ~pn5 & new_n473_;
  assign new_n475_ = pl5 & new_n474_;
  assign new_n476_ = ~pm5 & ~pl5;
  assign new_n477_ = ~pn5 & new_n476_;
  assign pv10 = pz | new_n477_;
  assign new_n479_ = ~new_n475_ & ~pv10;
  assign new_n480_ = ~pt4 & ~pu4;
  assign new_n481_ = ~pv4 & new_n480_;
  assign new_n482_ = ~pw4 & ~py4;
  assign new_n483_ = ~px4 & new_n482_;
  assign new_n484_ = new_n481_ & new_n483_;
  assign new_n485_ = ~ps4 & ~pz4;
  assign new_n486_ = new_n484_ & new_n485_;
  assign new_n487_ = pr4 & new_n486_;
  assign new_n488_ = ~new_n475_ & ~new_n487_;
  assign new_n489_ = ~new_n479_ & ~new_n488_;
  assign new_n490_ = ~pr5 & ~new_n480_;
  assign new_n491_ = ~pq5 & new_n490_;
  assign new_n492_ = ~new_n480_ & ~new_n484_;
  assign new_n493_ = ~pq5 & new_n492_;
  assign new_n494_ = ~pp5 & ~pr5;
  assign new_n495_ = ~pq5 & new_n494_;
  assign new_n496_ = ~pp5 & ~new_n484_;
  assign new_n497_ = ~pq5 & new_n496_;
  assign new_n498_ = ~pr4 & ps4;
  assign new_n499_ = ~new_n480_ & ~new_n481_;
  assign new_n500_ = ~pr5 & new_n499_;
  assign new_n501_ = ~new_n484_ & new_n499_;
  assign new_n502_ = ~pr5 & ~new_n481_;
  assign new_n503_ = ~pp5 & new_n502_;
  assign new_n504_ = ~new_n481_ & ~new_n484_;
  assign new_n505_ = ~pp5 & new_n504_;
  assign new_n506_ = ~new_n503_ & ~new_n505_;
  assign new_n507_ = ~new_n500_ & ~new_n501_;
  assign new_n508_ = new_n506_ & new_n507_;
  assign new_n509_ = ~new_n491_ & ~new_n493_;
  assign new_n510_ = ~new_n495_ & new_n509_;
  assign new_n511_ = ~new_n497_ & new_n498_;
  assign new_n512_ = new_n510_ & new_n511_;
  assign new_n513_ = new_n508_ & new_n512_;
  assign new_n514_ = pv10 & new_n513_;
  assign new_n515_ = ~pf0 & ~new_n514_;
  assign new_n516_ = ~pg5 & ~po5;
  assign new_n517_ = po5 & ~pi5;
  assign new_n518_ = ~new_n516_ & ~new_n517_;
  assign new_n519_ = pg5 & ~new_n518_;
  assign new_n520_ = pa5 & ~pb5;
  assign new_n521_ = new_n519_ & ~new_n520_;
  assign new_n522_ = ~new_n519_ & new_n520_;
  assign new_n523_ = ~new_n521_ & ~new_n522_;
  assign new_n524_ = ~pe5 & ~pd5;
  assign new_n525_ = ~new_n523_ & new_n524_;
  assign new_n526_ = new_n520_ & new_n525_;
  assign pj10 = pe5 | new_n526_;
  assign new_n528_ = ~pc5 & ~pj10;
  assign new_n529_ = ~pg0 & new_n528_;
  assign new_n530_ = ~pv3 & ~pu3;
  assign new_n531_ = ~pw3 & new_n530_;
  assign new_n532_ = ~pi0 & ~new_n531_;
  assign new_n533_ = ~py3 & ~new_n532_;
  assign new_n534_ = ~px3 & new_n533_;
  assign new_n535_ = ~pz3 & new_n534_;
  assign new_n536_ = ~pi0 & ~new_n535_;
  assign new_n537_ = ~pa4 & ~new_n536_;
  assign new_n538_ = new_n529_ & ~new_n537_;
  assign new_n539_ = pv3 & pu3;
  assign new_n540_ = pw3 & new_n539_;
  assign new_n541_ = ~pi0 & ~new_n540_;
  assign new_n542_ = py3 & ~new_n541_;
  assign new_n543_ = px3 & new_n542_;
  assign new_n544_ = pz3 & new_n543_;
  assign new_n545_ = ~pi0 & ~new_n544_;
  assign new_n546_ = pa4 & ~new_n545_;
  assign new_n547_ = ~new_n529_ & ~new_n546_;
  assign new_n548_ = ~new_n537_ & ~new_n546_;
  assign new_n549_ = ~new_n538_ & ~new_n547_;
  assign new_n550_ = ~new_n548_ & new_n549_;
  assign new_n551_ = ~new_n515_ & new_n550_;
  assign new_n552_ = ~pb4 & new_n551_;
  assign new_n553_ = pb4 & ~new_n551_;
  assign new_n554_ = ~new_n552_ & ~new_n553_;
  assign new_n555_ = ~new_n489_ & new_n554_;
  assign new_n556_ = ~ps3 & new_n489_;
  assign new_n557_ = ~ps3 & new_n554_;
  assign new_n558_ = ~new_n555_ & ~new_n556_;
  assign new_n559_ = ~new_n557_ & new_n558_;
  assign pi9 = pz | new_n559_;
  assign new_n561_ = pk5 & ~pj5;
  assign new_n562_ = ~pz & ~new_n561_;
  assign new_n563_ = ~pz & ~pn5;
  assign new_n564_ = pm5 & pl5;
  assign new_n565_ = new_n563_ & new_n564_;
  assign new_n566_ = pj5 & new_n565_;
  assign new_n567_ = ~pj5 & ~new_n565_;
  assign new_n568_ = ~new_n566_ & ~new_n567_;
  assign pq10 = new_n562_ & new_n568_;
  assign new_n570_ = new_n388_ & ~new_n390_;
  assign new_n571_ = new_n388_ & new_n398_;
  assign new_n572_ = new_n390_ & new_n398_;
  assign new_n573_ = ~new_n570_ & ~new_n571_;
  assign new_n574_ = ~new_n572_ & new_n573_;
  assign new_n575_ = ~new_n381_ & new_n574_;
  assign new_n576_ = ~py1 & new_n575_;
  assign new_n577_ = py1 & ~new_n575_;
  assign new_n578_ = ~new_n576_ & ~new_n577_;
  assign new_n579_ = ~pc3 & new_n578_;
  assign new_n580_ = ~new_n416_ & new_n578_;
  assign new_n581_ = ~pc3 & new_n416_;
  assign new_n582_ = ~new_n579_ & ~new_n580_;
  assign new_n583_ = ~new_n581_ & new_n582_;
  assign pf7 = ~pb & new_n583_;
  assign new_n585_ = pw0 & py0;
  assign new_n586_ = pv0 & px0;
  assign new_n587_ = new_n585_ & new_n586_;
  assign new_n588_ = ~new_n346_ & new_n587_;
  assign new_n589_ = ~pz0 & ~new_n588_;
  assign new_n590_ = pz0 & new_n588_;
  assign new_n591_ = ~new_n589_ & ~new_n590_;
  assign pg6 = new_n342_ & new_n591_;
  assign new_n593_ = new_n529_ & new_n536_;
  assign new_n594_ = ~new_n529_ & new_n545_;
  assign new_n595_ = new_n536_ & new_n545_;
  assign new_n596_ = ~new_n593_ & ~new_n594_;
  assign new_n597_ = ~new_n595_ & new_n596_;
  assign new_n598_ = ~new_n515_ & new_n597_;
  assign new_n599_ = ~pa4 & new_n598_;
  assign new_n600_ = pa4 & ~new_n598_;
  assign new_n601_ = ~new_n599_ & ~new_n600_;
  assign new_n602_ = ~new_n489_ & new_n601_;
  assign new_n603_ = ~pr3 & new_n489_;
  assign new_n604_ = ~pr3 & new_n601_;
  assign new_n605_ = ~new_n602_ & ~new_n603_;
  assign new_n606_ = ~new_n604_ & new_n605_;
  assign ph9 = ~pz & new_n606_;
  assign new_n608_ = pa3 & new_n453_;
  assign new_n609_ = ~pj & ~new_n608_;
  assign new_n610_ = ~new_n423_ & new_n609_;
  assign new_n611_ = ~pa3 & new_n462_;
  assign new_n612_ = ~pj & ~new_n611_;
  assign new_n613_ = new_n609_ & new_n612_;
  assign new_n614_ = new_n423_ & new_n612_;
  assign new_n615_ = ~new_n610_ & ~new_n613_;
  assign new_n616_ = ~new_n614_ & new_n615_;
  assign new_n617_ = ~new_n441_ & new_n616_;
  assign new_n618_ = ~pb3 & new_n617_;
  assign new_n619_ = pb3 & ~new_n617_;
  assign new_n620_ = ~new_n618_ & ~new_n619_;
  assign new_n621_ = new_n427_ & ~new_n620_;
  assign pi8 = new_n428_ | new_n621_;
  assign new_n623_ = pv0 & ~new_n346_;
  assign new_n624_ = ~pw0 & ~new_n623_;
  assign new_n625_ = pw0 & new_n623_;
  assign new_n626_ = ~new_n624_ & ~new_n625_;
  assign pd6 = new_n342_ & new_n626_;
  assign new_n628_ = pv1 & ~new_n384_;
  assign new_n629_ = pw1 & new_n628_;
  assign new_n630_ = ~new_n390_ & ~new_n629_;
  assign new_n631_ = ~pw1 & ~pv1;
  assign new_n632_ = ~new_n394_ & new_n631_;
  assign new_n633_ = ~new_n629_ & ~new_n632_;
  assign new_n634_ = new_n390_ & ~new_n632_;
  assign new_n635_ = ~new_n630_ & ~new_n633_;
  assign new_n636_ = ~new_n634_ & new_n635_;
  assign new_n637_ = ~new_n381_ & new_n636_;
  assign new_n638_ = ~px1 & new_n637_;
  assign new_n639_ = px1 & ~new_n637_;
  assign new_n640_ = ~new_n638_ & ~new_n639_;
  assign new_n641_ = ~pb3 & new_n640_;
  assign new_n642_ = ~new_n416_ & new_n640_;
  assign new_n643_ = ~pb3 & new_n416_;
  assign new_n644_ = ~new_n641_ & ~new_n642_;
  assign new_n645_ = ~new_n643_ & new_n644_;
  assign pe7 = pb | new_n645_;
  assign new_n647_ = pb3 & ~new_n609_;
  assign new_n648_ = ~new_n423_ & ~new_n647_;
  assign new_n649_ = ~pb3 & ~new_n612_;
  assign new_n650_ = ~new_n647_ & ~new_n649_;
  assign new_n651_ = new_n423_ & ~new_n649_;
  assign new_n652_ = ~new_n648_ & ~new_n650_;
  assign new_n653_ = ~new_n651_ & new_n652_;
  assign new_n654_ = ~new_n441_ & new_n653_;
  assign new_n655_ = ~pc3 & ~new_n654_;
  assign new_n656_ = pc3 & new_n654_;
  assign new_n657_ = ~new_n655_ & ~new_n656_;
  assign pj8 = new_n427_ & new_n657_;
  assign pk9 = ~pd4 | pz;
  assign new_n660_ = pm5 & ~pz;
  assign new_n661_ = ~pn5 & new_n660_;
  assign new_n662_ = ~pl5 & new_n661_;
  assign new_n663_ = new_n520_ & new_n662_;
  assign new_n664_ = pq3 & pp3;
  assign new_n665_ = ps3 & new_n664_;
  assign new_n666_ = pr3 & new_n665_;
  assign new_n667_ = pt3 & new_n666_;
  assign new_n668_ = ~pr3 & ~pt3;
  assign new_n669_ = ~ps3 & ~pq3;
  assign new_n670_ = new_n668_ & new_n669_;
  assign new_n671_ = ~po3 & ~pp3;
  assign new_n672_ = pn3 & new_n671_;
  assign new_n673_ = new_n670_ & new_n672_;
  assign new_n674_ = new_n520_ & new_n667_;
  assign new_n675_ = ~new_n673_ & new_n674_;
  assign new_n676_ = new_n565_ & ~new_n675_;
  assign new_n677_ = ~new_n475_ & ~new_n663_;
  assign new_n678_ = ~new_n676_ & new_n677_;
  assign ps10 = ~pz & ~new_n678_;
  assign new_n680_ = ~new_n390_ & ~new_n628_;
  assign new_n681_ = ~pv1 & ~new_n394_;
  assign new_n682_ = ~new_n628_ & ~new_n681_;
  assign new_n683_ = new_n390_ & ~new_n681_;
  assign new_n684_ = ~new_n680_ & ~new_n682_;
  assign new_n685_ = ~new_n683_ & new_n684_;
  assign new_n686_ = ~new_n381_ & new_n685_;
  assign new_n687_ = ~pw1 & new_n686_;
  assign new_n688_ = pw1 & ~new_n686_;
  assign new_n689_ = ~new_n687_ & ~new_n688_;
  assign new_n690_ = ~pa3 & new_n689_;
  assign new_n691_ = ~new_n416_ & new_n689_;
  assign new_n692_ = ~pa3 & new_n416_;
  assign new_n693_ = ~new_n690_ & ~new_n691_;
  assign new_n694_ = ~new_n692_ & new_n693_;
  assign pd7 = pb | new_n694_;
  assign new_n696_ = pv0 & new_n347_;
  assign new_n697_ = ~px0 & ~new_n696_;
  assign new_n698_ = px0 & new_n696_;
  assign new_n699_ = ~new_n697_ & ~new_n698_;
  assign pe6 = new_n342_ & new_n699_;
  assign new_n701_ = ~pa4 & ~pb4;
  assign new_n702_ = ~new_n536_ & new_n701_;
  assign new_n703_ = new_n529_ & ~new_n702_;
  assign new_n704_ = pb4 & new_n546_;
  assign new_n705_ = ~new_n529_ & ~new_n704_;
  assign new_n706_ = ~new_n702_ & ~new_n704_;
  assign new_n707_ = ~new_n703_ & ~new_n705_;
  assign new_n708_ = ~new_n706_ & new_n707_;
  assign new_n709_ = ~new_n515_ & new_n708_;
  assign new_n710_ = ~pc4 & new_n709_;
  assign new_n711_ = pc4 & ~new_n709_;
  assign new_n712_ = ~new_n710_ & ~new_n711_;
  assign new_n713_ = ~new_n489_ & new_n712_;
  assign new_n714_ = ~pt3 & new_n489_;
  assign new_n715_ = ~pt3 & new_n712_;
  assign new_n716_ = ~new_n713_ & ~new_n714_;
  assign new_n717_ = ~new_n715_ & new_n716_;
  assign pj9 = pz | new_n717_;
  assign new_n719_ = pc3 & new_n647_;
  assign new_n720_ = ~new_n423_ & ~new_n719_;
  assign new_n721_ = ~pc3 & new_n649_;
  assign new_n722_ = ~new_n719_ & ~new_n721_;
  assign new_n723_ = new_n423_ & ~new_n721_;
  assign new_n724_ = ~new_n720_ & ~new_n722_;
  assign new_n725_ = ~new_n723_ & new_n724_;
  assign new_n726_ = ~new_n441_ & new_n725_;
  assign new_n727_ = ~pd3 & new_n726_;
  assign new_n728_ = pd3 & ~new_n726_;
  assign new_n729_ = ~new_n727_ & ~new_n728_;
  assign new_n730_ = new_n427_ & ~new_n729_;
  assign pk8 = new_n428_ | new_n730_;
  assign new_n732_ = ~pk5 & ~new_n566_;
  assign new_n733_ = pk5 & new_n566_;
  assign new_n734_ = ~new_n732_ & ~new_n733_;
  assign pr10 = new_n562_ & new_n734_;
  assign new_n736_ = pn0 & pq5;
  assign new_n737_ = pn5 & pp0;
  assign new_n738_ = ~pz & ~new_n662_;
  assign new_n739_ = po0 & ~new_n738_;
  assign new_n740_ = ~pj0 & ~pp5;
  assign new_n741_ = pd4 & pe4;
  assign new_n742_ = pf4 & new_n741_;
  assign new_n743_ = ~pj0 & pq5;
  assign new_n744_ = ~new_n742_ & ~new_n743_;
  assign new_n745_ = pi4 & ~new_n744_;
  assign new_n746_ = new_n740_ & ~new_n745_;
  assign new_n747_ = pg4 & pp4;
  assign new_n748_ = ~new_n746_ & new_n747_;
  assign new_n749_ = pq0 & new_n748_;
  assign new_n750_ = ~new_n736_ & ~new_n737_;
  assign new_n751_ = ~new_n739_ & ~new_n749_;
  assign new_n752_ = new_n750_ & new_n751_;
  assign new_n753_ = pl0 & pl3;
  assign new_n754_ = pk0 & new_n673_;
  assign new_n755_ = pm0 & new_n667_;
  assign new_n756_ = ~new_n753_ & ~new_n754_;
  assign new_n757_ = ~new_n755_ & new_n756_;
  assign new_n758_ = pg4 & pr0;
  assign new_n759_ = pv4 & pt0;
  assign new_n760_ = pr5 & ~pv10;
  assign new_n761_ = ~pr4 & new_n760_;
  assign new_n762_ = ~pv10 & ~new_n561_;
  assign new_n763_ = new_n519_ & ~new_n523_;
  assign new_n764_ = new_n524_ & new_n763_;
  assign new_n765_ = ~pd5 & ~new_n764_;
  assign new_n766_ = new_n528_ & new_n765_;
  assign new_n767_ = ~pr4 & new_n486_;
  assign new_n768_ = ~new_n766_ & new_n767_;
  assign new_n769_ = pr5 & ~new_n768_;
  assign new_n770_ = ~pr4 & new_n769_;
  assign new_n771_ = ~new_n561_ & ~new_n768_;
  assign new_n772_ = ~new_n761_ & ~new_n762_;
  assign new_n773_ = ~new_n770_ & ~new_n771_;
  assign new_n774_ = new_n772_ & new_n773_;
  assign new_n775_ = ~pd0 & ~new_n774_;
  assign new_n776_ = ps0 & new_n775_;
  assign new_n777_ = pl5 & pu0;
  assign new_n778_ = ~new_n758_ & ~new_n759_;
  assign new_n779_ = ~new_n776_ & ~new_n777_;
  assign new_n780_ = new_n778_ & new_n779_;
  assign new_n781_ = new_n752_ & new_n757_;
  assign pb6 = ~new_n780_ | ~new_n781_;
  assign new_n783_ = new_n384_ & ~new_n390_;
  assign new_n784_ = new_n384_ & new_n394_;
  assign new_n785_ = new_n390_ & new_n394_;
  assign new_n786_ = ~new_n783_ & ~new_n784_;
  assign new_n787_ = ~new_n785_ & new_n786_;
  assign new_n788_ = ~new_n381_ & new_n787_;
  assign new_n789_ = ~pv1 & new_n788_;
  assign new_n790_ = pv1 & ~new_n788_;
  assign new_n791_ = ~new_n789_ & ~new_n790_;
  assign new_n792_ = ~pz2 & new_n791_;
  assign new_n793_ = ~new_n416_ & new_n791_;
  assign new_n794_ = ~pz2 & new_n416_;
  assign new_n795_ = ~new_n792_ & ~new_n793_;
  assign new_n796_ = ~new_n794_ & new_n795_;
  assign pc7 = pb | new_n796_;
  assign new_n798_ = pd3 & new_n719_;
  assign new_n799_ = ~new_n423_ & ~new_n798_;
  assign new_n800_ = ~pc3 & ~pd3;
  assign new_n801_ = new_n649_ & new_n800_;
  assign new_n802_ = ~new_n798_ & ~new_n801_;
  assign new_n803_ = new_n423_ & ~new_n801_;
  assign new_n804_ = ~new_n799_ & ~new_n802_;
  assign new_n805_ = ~new_n803_ & new_n804_;
  assign new_n806_ = ~new_n441_ & new_n805_;
  assign new_n807_ = ~pe3 & new_n806_;
  assign new_n808_ = pe3 & ~new_n806_;
  assign new_n809_ = ~new_n807_ & ~new_n808_;
  assign new_n810_ = new_n427_ & ~new_n809_;
  assign pl8 = new_n428_ | new_n810_;
  assign new_n812_ = ~pf4 & ~new_n741_;
  assign new_n813_ = ~new_n742_ & ~new_n812_;
  assign pm9 = pz | new_n813_;
  assign new_n815_ = pn5 & new_n660_;
  assign new_n816_ = pl5 & new_n815_;
  assign new_n817_ = ~new_n667_ & ~new_n816_;
  assign new_n818_ = ~new_n520_ & ~new_n816_;
  assign new_n819_ = new_n673_ & ~new_n816_;
  assign new_n820_ = ~new_n565_ & ~new_n816_;
  assign new_n821_ = ~new_n817_ & ~new_n818_;
  assign new_n822_ = ~new_n819_ & ~new_n820_;
  assign new_n823_ = new_n821_ & new_n822_;
  assign new_n824_ = pn5 & new_n473_;
  assign new_n825_ = ~pl5 & new_n824_;
  assign new_n826_ = ~new_n475_ & ~new_n825_;
  assign new_n827_ = ~new_n673_ & new_n826_;
  assign new_n828_ = ~new_n565_ & new_n826_;
  assign new_n829_ = ~new_n827_ & ~new_n828_;
  assign new_n830_ = ~new_n823_ & ~new_n829_;
  assign pu10 = ~pz & ~new_n830_;
  assign new_n832_ = ~new_n382_ & ~new_n390_;
  assign new_n833_ = ~new_n382_ & ~new_n392_;
  assign new_n834_ = new_n390_ & ~new_n392_;
  assign new_n835_ = ~new_n832_ & ~new_n833_;
  assign new_n836_ = ~new_n834_ & new_n835_;
  assign new_n837_ = ~new_n381_ & new_n836_;
  assign new_n838_ = ~pu1 & new_n837_;
  assign new_n839_ = pu1 & ~new_n837_;
  assign new_n840_ = ~new_n838_ & ~new_n839_;
  assign new_n841_ = ~py2 & new_n840_;
  assign new_n842_ = ~new_n416_ & new_n840_;
  assign new_n843_ = ~py2 & new_n416_;
  assign new_n844_ = ~new_n841_ & ~new_n842_;
  assign new_n845_ = ~new_n843_ & new_n844_;
  assign pb7 = ~pb & new_n845_;
  assign new_n847_ = ~pv0 & new_n346_;
  assign new_n848_ = ~new_n623_ & ~new_n847_;
  assign pc6 = new_n342_ & new_n848_;
  assign new_n850_ = ~pd4 & ~pe4;
  assign new_n851_ = ~new_n741_ & ~new_n850_;
  assign pl9 = pz | new_n851_;
  assign new_n853_ = ~pf3 & new_n775_;
  assign new_n854_ = pf3 & ~new_n775_;
  assign new_n855_ = ~new_n853_ & ~new_n854_;
  assign pm8 = new_n738_ & new_n855_;
  assign new_n857_ = ~pm5 & ~new_n816_;
  assign new_n858_ = ~new_n565_ & new_n857_;
  assign new_n859_ = new_n520_ & new_n857_;
  assign new_n860_ = ~pn5 & ~new_n816_;
  assign new_n861_ = new_n520_ & new_n860_;
  assign new_n862_ = new_n673_ & new_n860_;
  assign new_n863_ = ~new_n565_ & new_n860_;
  assign new_n864_ = new_n673_ & new_n857_;
  assign new_n865_ = ~new_n858_ & ~new_n859_;
  assign new_n866_ = ~new_n861_ & new_n865_;
  assign new_n867_ = ~new_n862_ & ~new_n863_;
  assign new_n868_ = ~new_n864_ & new_n867_;
  assign new_n869_ = new_n866_ & new_n868_;
  assign new_n870_ = new_n565_ & new_n673_;
  assign new_n871_ = ~pr5 & new_n528_;
  assign new_n872_ = new_n528_ & ~new_n565_;
  assign new_n873_ = ~new_n871_ & ~new_n872_;
  assign new_n874_ = new_n765_ & ~new_n873_;
  assign new_n875_ = py4 & ~new_n874_;
  assign new_n876_ = pw4 & px4;
  assign new_n877_ = pv4 & new_n876_;
  assign new_n878_ = pu4 & ps4;
  assign new_n879_ = pt4 & pr4;
  assign new_n880_ = new_n878_ & new_n879_;
  assign new_n881_ = new_n877_ & new_n880_;
  assign new_n882_ = new_n875_ & new_n881_;
  assign new_n883_ = pz4 & new_n882_;
  assign new_n884_ = ~pz4 & ~new_n883_;
  assign new_n885_ = ~pa0 & new_n884_;
  assign new_n886_ = pr5 & ~new_n883_;
  assign new_n887_ = ~pa0 & new_n886_;
  assign new_n888_ = ~pr5 & ~pz4;
  assign new_n889_ = ~pa0 & new_n888_;
  assign new_n890_ = ~new_n885_ & ~new_n887_;
  assign new_n891_ = ~new_n889_ & new_n890_;
  assign new_n892_ = pv10 & new_n891_;
  assign new_n893_ = ~new_n870_ & ~new_n892_;
  assign new_n894_ = ~new_n662_ & ~new_n825_;
  assign new_n895_ = new_n893_ & new_n894_;
  assign new_n896_ = ~new_n869_ & new_n895_;
  assign pt10 = ~pz & ~new_n896_;
  assign new_n898_ = ~ps1 & ~new_n390_;
  assign new_n899_ = ps1 & new_n390_;
  assign new_n900_ = ~new_n898_ & ~new_n899_;
  assign new_n901_ = ~new_n381_ & new_n900_;
  assign new_n902_ = ~pt1 & new_n901_;
  assign new_n903_ = pt1 & ~new_n901_;
  assign new_n904_ = ~new_n902_ & ~new_n903_;
  assign new_n905_ = ~px2 & new_n904_;
  assign new_n906_ = ~new_n416_ & new_n904_;
  assign new_n907_ = ~px2 & new_n416_;
  assign new_n908_ = ~new_n905_ & ~new_n906_;
  assign new_n909_ = ~new_n907_ & new_n908_;
  assign pa7 = ~pb & new_n909_;
  assign new_n911_ = pv10 & ~new_n528_;
  assign new_n912_ = ~pe0 & ~new_n911_;
  assign new_n913_ = ~pf3 & ~new_n912_;
  assign new_n914_ = pf3 & new_n912_;
  assign new_n915_ = ~new_n913_ & ~new_n914_;
  assign new_n916_ = ~new_n775_ & new_n915_;
  assign new_n917_ = ~pg3 & ~new_n916_;
  assign new_n918_ = pg3 & new_n916_;
  assign new_n919_ = ~new_n917_ & ~new_n918_;
  assign pn8 = new_n738_ & new_n919_;
  assign new_n921_ = pl5 & pn5;
  assign new_n922_ = new_n473_ & new_n921_;
  assign new_n923_ = ~new_n748_ & ~new_n922_;
  assign new_n924_ = ~pv3 & ~new_n923_;
  assign new_n925_ = pg4 & ~new_n746_;
  assign new_n926_ = ~ph4 & new_n925_;
  assign new_n927_ = ph4 & ~new_n925_;
  assign new_n928_ = ~new_n926_ & ~new_n927_;
  assign new_n929_ = new_n923_ & new_n928_;
  assign new_n930_ = ~pv3 & new_n928_;
  assign new_n931_ = ~new_n924_ & ~new_n929_;
  assign new_n932_ = ~new_n930_ & new_n931_;
  assign po9 = pz | new_n932_;
  assign new_n934_ = ~pb0 & ~new_n825_;
  assign new_n935_ = ~pr5 & new_n934_;
  assign new_n936_ = ~pp5 & new_n935_;
  assign new_n937_ = ~pc0 & ~new_n816_;
  assign new_n938_ = new_n934_ & new_n937_;
  assign new_n939_ = ~pp5 & new_n938_;
  assign new_n940_ = ~pq5 & new_n937_;
  assign new_n941_ = ~pp5 & new_n940_;
  assign new_n942_ = ~pr5 & ~new_n937_;
  assign new_n943_ = ~pq5 & new_n942_;
  assign new_n944_ = ~pq5 & ~pr5;
  assign new_n945_ = ~pp5 & new_n944_;
  assign new_n946_ = ~new_n934_ & new_n937_;
  assign new_n947_ = ~pq5 & new_n946_;
  assign new_n948_ = new_n934_ & ~new_n937_;
  assign new_n949_ = ~pr5 & new_n948_;
  assign new_n950_ = ~pr5 & ~new_n934_;
  assign new_n951_ = ~pq5 & new_n950_;
  assign new_n952_ = ~new_n936_ & ~new_n939_;
  assign new_n953_ = ~new_n941_ & ~new_n943_;
  assign new_n954_ = new_n952_ & new_n953_;
  assign new_n955_ = ~new_n949_ & ~new_n951_;
  assign new_n956_ = ~new_n945_ & ~new_n947_;
  assign new_n957_ = new_n955_ & new_n956_;
  assign new_n958_ = new_n954_ & new_n957_;
  assign new_n959_ = ~pq5 & ~pp5;
  assign new_n960_ = ~new_n494_ & ~new_n944_;
  assign new_n961_ = ~new_n959_ & new_n960_;
  assign new_n962_ = ~pz & ~new_n961_;
  assign new_n963_ = pr5 & new_n962_;
  assign new_n964_ = pq5 & new_n962_;
  assign new_n965_ = pp5 & new_n962_;
  assign new_n966_ = ~new_n963_ & ~new_n964_;
  assign new_n967_ = ~new_n965_ & new_n966_;
  assign pw10 = new_n958_ | new_n967_;
  assign new_n969_ = pn0 & pp5;
  assign new_n970_ = pm5 & pp0;
  assign new_n971_ = po0 & pr5;
  assign new_n972_ = pm4 & pq0;
  assign new_n973_ = ~new_n969_ & ~new_n970_;
  assign new_n974_ = ~new_n971_ & ~new_n972_;
  assign new_n975_ = new_n973_ & new_n974_;
  assign new_n976_ = pl0 & pm3;
  assign new_n977_ = pk0 & pq3;
  assign new_n978_ = pf3 & pm0;
  assign new_n979_ = ~new_n976_ & ~new_n977_;
  assign new_n980_ = ~new_n978_ & new_n979_;
  assign new_n981_ = ph4 & pr0;
  assign new_n982_ = pw4 & pt0;
  assign new_n983_ = pd4 & ps0;
  assign new_n984_ = pu0 & pr4;
  assign new_n985_ = ~new_n981_ & ~new_n982_;
  assign new_n986_ = ~new_n983_ & ~new_n984_;
  assign new_n987_ = new_n985_ & new_n986_;
  assign new_n988_ = new_n975_ & new_n980_;
  assign pa6 = ~new_n987_ | ~new_n988_;
  assign new_n990_ = ~pu3 & ~new_n923_;
  assign new_n991_ = ~pg4 & ~new_n746_;
  assign new_n992_ = pg4 & new_n746_;
  assign new_n993_ = ~new_n991_ & ~new_n992_;
  assign new_n994_ = new_n923_ & new_n993_;
  assign new_n995_ = ~pu3 & new_n993_;
  assign new_n996_ = ~new_n990_ & ~new_n994_;
  assign new_n997_ = ~new_n995_ & new_n996_;
  assign pn9 = pz | new_n997_;
  assign new_n999_ = ~pg3 & ~pf3;
  assign new_n1000_ = pq5 & new_n565_;
  assign new_n1001_ = ~ph0 & new_n1000_;
  assign new_n1002_ = ~new_n999_ & ~new_n1001_;
  assign new_n1003_ = new_n912_ & new_n1002_;
  assign new_n1004_ = pg3 & pf3;
  assign new_n1005_ = ~new_n1001_ & ~new_n1004_;
  assign new_n1006_ = ~new_n912_ & new_n1005_;
  assign new_n1007_ = new_n1002_ & new_n1005_;
  assign new_n1008_ = ~new_n1003_ & ~new_n1006_;
  assign new_n1009_ = ~new_n1007_ & new_n1008_;
  assign new_n1010_ = ~new_n775_ & new_n1009_;
  assign new_n1011_ = ~ph3 & ~new_n1010_;
  assign new_n1012_ = ph3 & new_n1010_;
  assign new_n1013_ = ~new_n1011_ & ~new_n1012_;
  assign po8 = new_n738_ & new_n1013_;
  assign new_n1015_ = ~new_n738_ & ~new_n912_;
  assign new_n1016_ = pp5 & new_n565_;
  assign new_n1017_ = ~ph0 & new_n1016_;
  assign new_n1018_ = new_n1002_ & ~new_n1017_;
  assign new_n1019_ = ph3 & ~new_n1017_;
  assign new_n1020_ = ~new_n1018_ & ~new_n1019_;
  assign new_n1021_ = ~pi3 & new_n1020_;
  assign new_n1022_ = ~ph0 & ~new_n1021_;
  assign new_n1023_ = pj3 & ~new_n1022_;
  assign new_n1024_ = ~pp3 & new_n1023_;
  assign new_n1025_ = ~ph0 & ~new_n1024_;
  assign new_n1026_ = ~pq3 & ~new_n1025_;
  assign new_n1027_ = ~ps3 & ~pr3;
  assign new_n1028_ = new_n1026_ & new_n1027_;
  assign new_n1029_ = new_n912_ & ~new_n1028_;
  assign new_n1030_ = new_n1005_ & ~new_n1017_;
  assign new_n1031_ = ~ph3 & ~new_n1017_;
  assign new_n1032_ = ~new_n1030_ & ~new_n1031_;
  assign new_n1033_ = pi3 & new_n1032_;
  assign new_n1034_ = ~ph0 & ~new_n1033_;
  assign new_n1035_ = pk3 & ~new_n1034_;
  assign new_n1036_ = pp3 & new_n1035_;
  assign new_n1037_ = ~ph0 & ~new_n1036_;
  assign new_n1038_ = pq3 & ~new_n1037_;
  assign new_n1039_ = pr3 & new_n1038_;
  assign new_n1040_ = ps3 & new_n1039_;
  assign new_n1041_ = ~new_n912_ & ~new_n1040_;
  assign new_n1042_ = ~new_n1028_ & ~new_n1040_;
  assign new_n1043_ = ~new_n1029_ & ~new_n1041_;
  assign new_n1044_ = ~new_n1042_ & new_n1043_;
  assign new_n1045_ = ~new_n775_ & new_n1044_;
  assign new_n1046_ = ~pt3 & new_n1045_;
  assign new_n1047_ = pt3 & ~new_n1045_;
  assign new_n1048_ = ~new_n1046_ & ~new_n1047_;
  assign new_n1049_ = new_n738_ & ~new_n1048_;
  assign pa9 = new_n1015_ | new_n1049_;
  assign new_n1051_ = ~pp1 & ~pl;
  assign new_n1052_ = pb2 & pc2;
  assign new_n1053_ = pd2 & new_n1052_;
  assign new_n1054_ = pq1 & ~pl;
  assign new_n1055_ = ~new_n1053_ & ~new_n1054_;
  assign new_n1056_ = pg2 & ~new_n1055_;
  assign new_n1057_ = new_n1051_ & ~new_n1056_;
  assign new_n1058_ = pe2 & ~new_n1057_;
  assign new_n1059_ = pf2 & new_n1058_;
  assign new_n1060_ = ~ph2 & new_n1059_;
  assign new_n1061_ = ph2 & ~new_n1059_;
  assign new_n1062_ = ~new_n1060_ & ~new_n1061_;
  assign new_n1063_ = ~pu1 & new_n1062_;
  assign new_n1064_ = pe2 & pn2;
  assign new_n1065_ = ~new_n1057_ & new_n1064_;
  assign new_n1066_ = ~new_n313_ & ~new_n1065_;
  assign new_n1067_ = new_n1062_ & new_n1066_;
  assign new_n1068_ = ~pu1 & ~new_n1066_;
  assign new_n1069_ = ~new_n1063_ & ~new_n1067_;
  assign new_n1070_ = ~new_n1068_ & new_n1069_;
  assign po7 = pb | new_n1070_;
  assign new_n1072_ = ~pq5 & new_n935_;
  assign new_n1073_ = ~pr5 & new_n938_;
  assign new_n1074_ = ~pr5 & new_n937_;
  assign new_n1075_ = ~pp5 & new_n1074_;
  assign new_n1076_ = ~pq5 & ~new_n937_;
  assign new_n1077_ = ~pp5 & new_n1076_;
  assign new_n1078_ = ~pp5 & new_n946_;
  assign new_n1079_ = ~pq5 & new_n948_;
  assign new_n1080_ = ~pq5 & ~new_n934_;
  assign new_n1081_ = ~pp5 & new_n1080_;
  assign new_n1082_ = ~new_n1072_ & ~new_n1073_;
  assign new_n1083_ = ~new_n1075_ & ~new_n1077_;
  assign new_n1084_ = new_n1082_ & new_n1083_;
  assign new_n1085_ = ~new_n1079_ & ~new_n1081_;
  assign new_n1086_ = ~new_n945_ & ~new_n1078_;
  assign new_n1087_ = new_n1085_ & new_n1086_;
  assign new_n1088_ = new_n1084_ & new_n1087_;
  assign py10 = ~new_n967_ & new_n1088_;
  assign new_n1090_ = ~new_n423_ & new_n450_;
  assign new_n1091_ = new_n423_ & new_n459_;
  assign new_n1092_ = ~new_n1090_ & ~new_n1091_;
  assign new_n1093_ = ~new_n441_ & ~new_n1092_;
  assign new_n1094_ = ~pt2 & new_n1093_;
  assign new_n1095_ = pt2 & ~new_n1093_;
  assign new_n1096_ = ~new_n1094_ & ~new_n1095_;
  assign new_n1097_ = new_n427_ & ~new_n1096_;
  assign pa8 = new_n428_ | new_n1097_;
  assign new_n1099_ = ~pg2 & new_n1055_;
  assign new_n1100_ = ~new_n1056_ & ~new_n1099_;
  assign pn7 = pb | new_n1100_;
  assign new_n1102_ = ~pb & ~new_n313_;
  assign new_n1103_ = ~new_n323_ & new_n1102_;
  assign new_n1104_ = ~ph1 & new_n1102_;
  assign new_n1105_ = ~new_n1103_ & ~new_n1104_;
  assign new_n1106_ = ph1 & ~new_n1105_;
  assign po6 = new_n329_ | new_n1106_;
  assign new_n1108_ = ~pq5 & new_n934_;
  assign new_n1109_ = ~pp5 & new_n1108_;
  assign new_n1110_ = ~pq5 & new_n938_;
  assign new_n1111_ = ~pq5 & new_n1074_;
  assign new_n1112_ = ~pp5 & new_n942_;
  assign new_n1113_ = ~pr5 & new_n946_;
  assign new_n1114_ = ~pp5 & new_n948_;
  assign new_n1115_ = ~pp5 & new_n950_;
  assign new_n1116_ = ~new_n1109_ & ~new_n1110_;
  assign new_n1117_ = ~new_n1111_ & ~new_n1112_;
  assign new_n1118_ = new_n1116_ & new_n1117_;
  assign new_n1119_ = ~new_n1114_ & ~new_n1115_;
  assign new_n1120_ = ~new_n945_ & ~new_n1113_;
  assign new_n1121_ = new_n1119_ & new_n1120_;
  assign new_n1122_ = new_n1118_ & new_n1121_;
  assign px10 = ~new_n967_ & new_n1122_;
  assign new_n1124_ = ~pz2 & ~px2;
  assign new_n1125_ = ~pw2 & ~py2;
  assign new_n1126_ = new_n1124_ & new_n1125_;
  assign new_n1127_ = new_n423_ & new_n1126_;
  assign new_n1128_ = new_n427_ & new_n1126_;
  assign new_n1129_ = new_n423_ & ~new_n427_;
  assign new_n1130_ = ~new_n1127_ & ~new_n1128_;
  assign pb8 = new_n1129_ | ~new_n1130_;
  assign new_n1132_ = ~pu3 & ~new_n529_;
  assign new_n1133_ = pu3 & new_n529_;
  assign new_n1134_ = ~new_n1132_ & ~new_n1133_;
  assign new_n1135_ = ~new_n515_ & new_n1134_;
  assign new_n1136_ = ~pv3 & new_n1135_;
  assign new_n1137_ = pv3 & ~new_n1135_;
  assign new_n1138_ = ~new_n1136_ & ~new_n1137_;
  assign new_n1139_ = ~new_n489_ & new_n1138_;
  assign new_n1140_ = ~pm3 & new_n489_;
  assign new_n1141_ = ~pm3 & new_n1138_;
  assign new_n1142_ = ~new_n1139_ & ~new_n1140_;
  assign new_n1143_ = ~new_n1141_ & new_n1142_;
  assign pc9 = ~pz & new_n1143_;
  assign new_n1145_ = ~pf2 & new_n1058_;
  assign new_n1146_ = pf2 & ~new_n1058_;
  assign new_n1147_ = ~new_n1145_ & ~new_n1146_;
  assign new_n1148_ = ~pt1 & new_n1147_;
  assign new_n1149_ = new_n1066_ & new_n1147_;
  assign new_n1150_ = ~pt1 & ~new_n1066_;
  assign new_n1151_ = ~new_n1148_ & ~new_n1149_;
  assign new_n1152_ = ~new_n1150_ & new_n1151_;
  assign pm7 = pb | new_n1152_;
  assign new_n1154_ = ~pu3 & ~new_n515_;
  assign new_n1155_ = pu3 & new_n515_;
  assign new_n1156_ = ~new_n1154_ & ~new_n1155_;
  assign new_n1157_ = ~new_n489_ & new_n1156_;
  assign new_n1158_ = ~pl3 & new_n489_;
  assign new_n1159_ = ~pl3 & new_n1156_;
  assign new_n1160_ = ~new_n1157_ & ~new_n1158_;
  assign new_n1161_ = ~new_n1159_ & new_n1160_;
  assign pb9 = ~pz & new_n1161_;
  assign new_n1163_ = pz2 & px2;
  assign new_n1164_ = pw2 & py2;
  assign new_n1165_ = new_n1163_ & new_n1164_;
  assign pc8 = new_n427_ & new_n1165_;
  assign new_n1167_ = ~pe2 & ~new_n1057_;
  assign new_n1168_ = pe2 & new_n1057_;
  assign new_n1169_ = ~new_n1167_ & ~new_n1168_;
  assign new_n1170_ = ~ps1 & new_n1169_;
  assign new_n1171_ = new_n1066_ & new_n1169_;
  assign new_n1172_ = ~ps1 & ~new_n1066_;
  assign new_n1173_ = ~new_n1170_ & ~new_n1171_;
  assign new_n1174_ = ~new_n1172_ & new_n1173_;
  assign pl7 = pb | new_n1174_;
  assign new_n1176_ = ~new_n423_ & new_n452_;
  assign new_n1177_ = new_n452_ & new_n461_;
  assign new_n1178_ = new_n423_ & new_n461_;
  assign new_n1179_ = ~new_n1176_ & ~new_n1177_;
  assign new_n1180_ = ~new_n1178_ & new_n1179_;
  assign new_n1181_ = ~new_n441_ & new_n1180_;
  assign new_n1182_ = ~pw2 & ~new_n1181_;
  assign new_n1183_ = pw2 & new_n1181_;
  assign new_n1184_ = ~new_n1182_ & ~new_n1183_;
  assign pd8 = new_n427_ & new_n1184_;
  assign new_n1186_ = new_n529_ & new_n532_;
  assign new_n1187_ = ~new_n529_ & new_n541_;
  assign new_n1188_ = new_n532_ & new_n541_;
  assign new_n1189_ = ~new_n1186_ & ~new_n1187_;
  assign new_n1190_ = ~new_n1188_ & new_n1189_;
  assign new_n1191_ = ~new_n515_ & new_n1190_;
  assign new_n1192_ = ~px3 & new_n1191_;
  assign new_n1193_ = px3 & ~new_n1191_;
  assign new_n1194_ = ~new_n1192_ & ~new_n1193_;
  assign new_n1195_ = ~new_n489_ & new_n1194_;
  assign new_n1196_ = ~po3 & new_n489_;
  assign new_n1197_ = ~po3 & new_n1194_;
  assign new_n1198_ = ~new_n1195_ & ~new_n1196_;
  assign new_n1199_ = ~new_n1197_ & new_n1198_;
  assign pe9 = pz | new_n1199_;
  assign new_n1201_ = pa1 & pb1;
  assign new_n1202_ = pz0 & new_n1201_;
  assign new_n1203_ = ~new_n346_ & new_n1202_;
  assign new_n1204_ = new_n587_ & new_n1203_;
  assign new_n1205_ = ~pc1 & ~new_n1204_;
  assign new_n1206_ = pc1 & new_n1204_;
  assign new_n1207_ = ~new_n1205_ & ~new_n1206_;
  assign pj6 = new_n342_ & new_n1207_;
  assign new_n1209_ = ~pd2 & ~new_n1052_;
  assign new_n1210_ = ~new_n1053_ & ~new_n1209_;
  assign pk7 = pb | new_n1210_;
  assign new_n1212_ = new_n529_ & ~new_n530_;
  assign new_n1213_ = ~new_n529_ & ~new_n539_;
  assign new_n1214_ = ~new_n530_ & ~new_n539_;
  assign new_n1215_ = ~new_n1212_ & ~new_n1213_;
  assign new_n1216_ = ~new_n1214_ & new_n1215_;
  assign new_n1217_ = ~new_n515_ & new_n1216_;
  assign new_n1218_ = ~pw3 & new_n1217_;
  assign new_n1219_ = pw3 & ~new_n1217_;
  assign new_n1220_ = ~new_n1218_ & ~new_n1219_;
  assign new_n1221_ = ~new_n489_ & new_n1220_;
  assign new_n1222_ = ~pn3 & new_n489_;
  assign new_n1223_ = ~pn3 & new_n1220_;
  assign new_n1224_ = ~new_n1221_ & ~new_n1222_;
  assign new_n1225_ = ~new_n1223_ & new_n1224_;
  assign pd9 = ~pz & new_n1225_;
  assign new_n1227_ = pw2 & ~new_n452_;
  assign new_n1228_ = ~new_n423_ & ~new_n1227_;
  assign new_n1229_ = ~pw2 & ~new_n461_;
  assign new_n1230_ = ~new_n1227_ & ~new_n1229_;
  assign new_n1231_ = new_n423_ & ~new_n1229_;
  assign new_n1232_ = ~new_n1228_ & ~new_n1230_;
  assign new_n1233_ = ~new_n1231_ & new_n1232_;
  assign new_n1234_ = ~new_n441_ & new_n1233_;
  assign new_n1235_ = ~px2 & ~new_n1234_;
  assign new_n1236_ = px2 & new_n1234_;
  assign new_n1237_ = ~new_n1235_ & ~new_n1236_;
  assign pe8 = new_n427_ & new_n1237_;
  assign new_n1239_ = ~pb2 & ~pc2;
  assign new_n1240_ = ~new_n1052_ & ~new_n1239_;
  assign pj7 = pb | new_n1240_;
  assign new_n1242_ = pc1 & ~new_n346_;
  assign new_n1243_ = new_n587_ & new_n1202_;
  assign new_n1244_ = new_n1242_ & new_n1243_;
  assign new_n1245_ = pd1 & new_n1244_;
  assign new_n1246_ = ~pd1 & ~new_n1244_;
  assign new_n1247_ = ~new_n1245_ & ~new_n1246_;
  assign pk6 = new_n342_ & new_n1247_;
  assign new_n1249_ = px2 & new_n1227_;
  assign new_n1250_ = ~new_n423_ & ~new_n1249_;
  assign new_n1251_ = ~pw2 & ~px2;
  assign new_n1252_ = ~new_n461_ & new_n1251_;
  assign new_n1253_ = ~new_n1249_ & ~new_n1252_;
  assign new_n1254_ = new_n423_ & ~new_n1252_;
  assign new_n1255_ = ~new_n1250_ & ~new_n1253_;
  assign new_n1256_ = ~new_n1254_ & new_n1255_;
  assign new_n1257_ = ~new_n441_ & new_n1256_;
  assign new_n1258_ = ~py2 & ~new_n1257_;
  assign new_n1259_ = py2 & new_n1257_;
  assign new_n1260_ = ~new_n1258_ & ~new_n1259_;
  assign pf8 = new_n427_ & new_n1260_;
  assign new_n1262_ = ~py3 & ~px3;
  assign new_n1263_ = ~new_n532_ & new_n1262_;
  assign new_n1264_ = new_n529_ & ~new_n1263_;
  assign new_n1265_ = px3 & ~new_n541_;
  assign new_n1266_ = py3 & new_n1265_;
  assign new_n1267_ = ~new_n529_ & ~new_n1266_;
  assign new_n1268_ = ~new_n1263_ & ~new_n1266_;
  assign new_n1269_ = ~new_n1264_ & ~new_n1267_;
  assign new_n1270_ = ~new_n1268_ & new_n1269_;
  assign new_n1271_ = ~new_n515_ & new_n1270_;
  assign new_n1272_ = ~pz3 & new_n1271_;
  assign new_n1273_ = pz3 & ~new_n1271_;
  assign new_n1274_ = ~new_n1272_ & ~new_n1273_;
  assign new_n1275_ = ~new_n489_ & new_n1274_;
  assign new_n1276_ = ~pq3 & new_n489_;
  assign new_n1277_ = ~pq3 & new_n1274_;
  assign new_n1278_ = ~new_n1275_ & ~new_n1276_;
  assign new_n1279_ = ~new_n1277_ & new_n1278_;
  assign pg9 = pz | new_n1279_;
  assign new_n1281_ = pz0 & ~new_n346_;
  assign new_n1282_ = new_n587_ & new_n1281_;
  assign new_n1283_ = ~pa1 & ~new_n1282_;
  assign new_n1284_ = pa1 & new_n1282_;
  assign new_n1285_ = ~new_n1283_ & ~new_n1284_;
  assign ph6 = new_n342_ & new_n1285_;
  assign pi7 = ~pb2 | pb;
  assign new_n1288_ = ~px3 & ~new_n532_;
  assign new_n1289_ = new_n529_ & ~new_n1288_;
  assign new_n1290_ = ~new_n529_ & ~new_n1265_;
  assign new_n1291_ = ~new_n1265_ & ~new_n1288_;
  assign new_n1292_ = ~new_n1289_ & ~new_n1290_;
  assign new_n1293_ = ~new_n1291_ & new_n1292_;
  assign new_n1294_ = ~new_n515_ & new_n1293_;
  assign new_n1295_ = ~py3 & new_n1294_;
  assign new_n1296_ = py3 & ~new_n1294_;
  assign new_n1297_ = ~new_n1295_ & ~new_n1296_;
  assign new_n1298_ = ~new_n489_ & new_n1297_;
  assign new_n1299_ = ~pp3 & new_n489_;
  assign new_n1300_ = ~pp3 & new_n1297_;
  assign new_n1301_ = ~new_n1298_ & ~new_n1299_;
  assign new_n1302_ = ~new_n1300_ & new_n1301_;
  assign pf9 = pz | new_n1302_;
  assign new_n1304_ = px2 & ~new_n452_;
  assign new_n1305_ = pw2 & new_n1304_;
  assign new_n1306_ = py2 & new_n1305_;
  assign new_n1307_ = ~new_n423_ & ~new_n1306_;
  assign new_n1308_ = ~px2 & new_n1125_;
  assign new_n1309_ = ~new_n461_ & new_n1308_;
  assign new_n1310_ = ~new_n1306_ & ~new_n1309_;
  assign new_n1311_ = new_n423_ & ~new_n1309_;
  assign new_n1312_ = ~new_n1307_ & ~new_n1310_;
  assign new_n1313_ = ~new_n1311_ & new_n1312_;
  assign new_n1314_ = ~new_n441_ & new_n1313_;
  assign new_n1315_ = ~pz2 & new_n1314_;
  assign new_n1316_ = pz2 & ~new_n1314_;
  assign new_n1317_ = ~new_n1315_ & ~new_n1316_;
  assign new_n1318_ = new_n427_ & ~new_n1317_;
  assign pg8 = new_n428_ | new_n1318_;
  assign new_n1320_ = pz1 & new_n389_;
  assign new_n1321_ = ~new_n390_ & ~new_n1320_;
  assign new_n1322_ = ~py1 & ~pz1;
  assign new_n1323_ = ~new_n398_ & new_n1322_;
  assign new_n1324_ = ~new_n1320_ & ~new_n1323_;
  assign new_n1325_ = new_n390_ & ~new_n1323_;
  assign new_n1326_ = ~new_n1321_ & ~new_n1324_;
  assign new_n1327_ = ~new_n1325_ & new_n1326_;
  assign new_n1328_ = ~new_n381_ & new_n1327_;
  assign new_n1329_ = ~pa2 & new_n1328_;
  assign new_n1330_ = pa2 & ~new_n1328_;
  assign new_n1331_ = ~new_n1329_ & ~new_n1330_;
  assign new_n1332_ = ~pe3 & new_n1331_;
  assign new_n1333_ = ~new_n416_ & new_n1331_;
  assign new_n1334_ = ~pe3 & new_n416_;
  assign new_n1335_ = ~new_n1332_ & ~new_n1333_;
  assign new_n1336_ = ~new_n1334_ & new_n1335_;
  assign ph7 = pb | new_n1336_;
  assign new_n1338_ = pa1 & new_n1281_;
  assign new_n1339_ = new_n587_ & new_n1338_;
  assign new_n1340_ = ~pb1 & ~new_n1339_;
  assign new_n1341_ = pb1 & new_n1339_;
  assign new_n1342_ = ~new_n1340_ & ~new_n1341_;
  assign pi6 = new_n342_ & new_n1342_;
  assign new_n1344_ = pr4 & new_n565_;
  assign new_n1345_ = pr5 & new_n1344_;
  assign new_n1346_ = pv10 & new_n765_;
  assign new_n1347_ = new_n528_ & new_n1346_;
  assign new_n1348_ = ~new_n922_ & ~new_n1345_;
  assign new_n1349_ = ~pz & ~new_n1347_;
  assign new_n1350_ = new_n1348_ & new_n1349_;
  assign new_n1351_ = ps4 & ~new_n874_;
  assign new_n1352_ = pr4 & new_n1351_;
  assign new_n1353_ = ~pt4 & ~new_n1352_;
  assign new_n1354_ = pt4 & new_n1352_;
  assign new_n1355_ = ~new_n1353_ & ~new_n1354_;
  assign pa10 = new_n1350_ & new_n1355_;
  assign new_n1357_ = pp & py1;
  assign new_n1358_ = pr & ps1;
  assign new_n1359_ = pq & pv1;
  assign new_n1360_ = ps & pl2;
  assign new_n1361_ = ~new_n1357_ & ~new_n1358_;
  assign new_n1362_ = ~new_n1359_ & ~new_n1360_;
  assign new_n1363_ = new_n1361_ & new_n1362_;
  assign new_n1364_ = py2 & pn;
  assign new_n1365_ = pc3 & pm;
  assign new_n1366_ = pr2 & po;
  assign new_n1367_ = ~new_n1364_ & ~new_n1365_;
  assign new_n1368_ = ~new_n1366_ & new_n1367_;
  assign new_n1369_ = pt & ph2;
  assign new_n1370_ = pb1 & pv;
  assign new_n1371_ = pc2 & pu;
  assign new_n1372_ = pw & pw0;
  assign new_n1373_ = ~new_n1369_ & ~new_n1370_;
  assign new_n1374_ = ~new_n1371_ & ~new_n1372_;
  assign new_n1375_ = new_n1373_ & new_n1374_;
  assign new_n1376_ = new_n1363_ & new_n1368_;
  assign pu5 = ~new_n1375_ | ~new_n1376_;
  assign new_n1378_ = pj1 & new_n1065_;
  assign new_n1379_ = pp2 & ~new_n1378_;
  assign new_n1380_ = ~pa & new_n1378_;
  assign new_n1381_ = ~pa & pp2;
  assign new_n1382_ = ~new_n1379_ & ~new_n1380_;
  assign pw7 = new_n1381_ | ~new_n1382_;
  assign new_n1384_ = new_n912_ & new_n1025_;
  assign new_n1385_ = ~new_n912_ & new_n1037_;
  assign new_n1386_ = new_n1025_ & new_n1037_;
  assign new_n1387_ = ~new_n1384_ & ~new_n1385_;
  assign new_n1388_ = ~new_n1386_ & new_n1387_;
  assign new_n1389_ = ~new_n775_ & new_n1388_;
  assign new_n1390_ = ~pq3 & new_n1389_;
  assign new_n1391_ = pq3 & ~new_n1389_;
  assign new_n1392_ = ~new_n1390_ & ~new_n1391_;
  assign new_n1393_ = new_n738_ & ~new_n1392_;
  assign px8 = new_n1015_ | new_n1393_;
  assign new_n1395_ = ~pr4 & new_n874_;
  assign new_n1396_ = pr4 & ~new_n874_;
  assign new_n1397_ = ~new_n1395_ & ~new_n1396_;
  assign py9 = new_n1350_ & new_n1397_;
  assign new_n1399_ = pp & pz1;
  assign new_n1400_ = pr & pt1;
  assign new_n1401_ = pq & pw1;
  assign new_n1402_ = ps & pm2;
  assign new_n1403_ = ~new_n1399_ & ~new_n1400_;
  assign new_n1404_ = ~new_n1401_ & ~new_n1402_;
  assign new_n1405_ = new_n1403_ & new_n1404_;
  assign new_n1406_ = pz2 & pn;
  assign new_n1407_ = pd3 & pm;
  assign new_n1408_ = ps2 & po;
  assign new_n1409_ = ~new_n1406_ & ~new_n1407_;
  assign new_n1410_ = ~new_n1408_ & new_n1409_;
  assign new_n1411_ = pt & pi2;
  assign new_n1412_ = pc1 & pv;
  assign new_n1413_ = pu & pd2;
  assign new_n1414_ = pw & px0;
  assign new_n1415_ = ~new_n1411_ & ~new_n1412_;
  assign new_n1416_ = ~new_n1413_ & ~new_n1414_;
  assign new_n1417_ = new_n1415_ & new_n1416_;
  assign new_n1418_ = new_n1405_ & new_n1410_;
  assign pt5 = ~new_n1417_ | ~new_n1418_;
  assign new_n1420_ = ph2 & new_n1059_;
  assign new_n1421_ = pi2 & new_n1420_;
  assign new_n1422_ = pj2 & new_n1421_;
  assign new_n1423_ = ~pl & ~new_n1422_;
  assign new_n1424_ = pk2 & ~new_n1423_;
  assign new_n1425_ = pl2 & new_n1424_;
  assign new_n1426_ = pm2 & new_n1425_;
  assign new_n1427_ = ~po2 & new_n1426_;
  assign new_n1428_ = po2 & ~new_n1426_;
  assign new_n1429_ = ~new_n1427_ & ~new_n1428_;
  assign new_n1430_ = ~pa2 & new_n1429_;
  assign new_n1431_ = new_n1066_ & new_n1429_;
  assign new_n1432_ = ~pa2 & ~new_n1066_;
  assign new_n1433_ = ~new_n1430_ & ~new_n1431_;
  assign new_n1434_ = ~new_n1432_ & new_n1433_;
  assign pv7 = pb | new_n1434_;
  assign new_n1436_ = pn1 & new_n311_;
  assign new_n1437_ = ~pl1 & new_n1436_;
  assign new_n1438_ = ~pd & ~new_n1437_;
  assign new_n1439_ = ~pr1 & new_n1438_;
  assign new_n1440_ = ~pp1 & new_n1439_;
  assign new_n1441_ = pn1 & new_n424_;
  assign new_n1442_ = pl1 & new_n1441_;
  assign new_n1443_ = ~pe & ~new_n1442_;
  assign new_n1444_ = new_n1438_ & new_n1443_;
  assign new_n1445_ = ~pp1 & new_n1444_;
  assign new_n1446_ = ~pq1 & new_n1443_;
  assign new_n1447_ = ~pp1 & new_n1446_;
  assign new_n1448_ = ~pr1 & ~new_n1443_;
  assign new_n1449_ = ~pq1 & new_n1448_;
  assign new_n1450_ = ~pq1 & ~pr1;
  assign new_n1451_ = ~pp1 & new_n1450_;
  assign new_n1452_ = ~new_n1438_ & new_n1443_;
  assign new_n1453_ = ~pq1 & new_n1452_;
  assign new_n1454_ = new_n1438_ & ~new_n1443_;
  assign new_n1455_ = ~pr1 & new_n1454_;
  assign new_n1456_ = ~pr1 & ~new_n1438_;
  assign new_n1457_ = ~pq1 & new_n1456_;
  assign new_n1458_ = ~new_n1440_ & ~new_n1445_;
  assign new_n1459_ = ~new_n1447_ & ~new_n1449_;
  assign new_n1460_ = new_n1458_ & new_n1459_;
  assign new_n1461_ = ~new_n1455_ & ~new_n1457_;
  assign new_n1462_ = ~new_n1451_ & ~new_n1453_;
  assign new_n1463_ = new_n1461_ & new_n1462_;
  assign new_n1464_ = new_n1460_ & new_n1463_;
  assign new_n1465_ = ~pp1 & ~pr1;
  assign new_n1466_ = ~new_n1450_ & ~new_n1465_;
  assign new_n1467_ = ~new_n366_ & new_n1466_;
  assign new_n1468_ = ~pb & ~new_n1467_;
  assign new_n1469_ = pr1 & new_n1468_;
  assign new_n1470_ = pq1 & new_n1468_;
  assign new_n1471_ = pp1 & new_n1468_;
  assign new_n1472_ = ~new_n1469_ & ~new_n1470_;
  assign new_n1473_ = ~new_n1471_ & new_n1472_;
  assign pw6 = new_n1464_ | new_n1473_;
  assign new_n1475_ = ~pc4 & ~new_n923_;
  assign new_n1476_ = ph4 & new_n925_;
  assign new_n1477_ = pj4 & new_n1476_;
  assign new_n1478_ = pk4 & new_n1477_;
  assign new_n1479_ = pl4 & new_n1478_;
  assign new_n1480_ = ~pj0 & ~new_n1479_;
  assign new_n1481_ = pm4 & ~new_n1480_;
  assign new_n1482_ = pn4 & new_n1481_;
  assign new_n1483_ = po4 & new_n1482_;
  assign new_n1484_ = ~pq4 & new_n1483_;
  assign new_n1485_ = pq4 & ~new_n1483_;
  assign new_n1486_ = ~new_n1484_ & ~new_n1485_;
  assign new_n1487_ = new_n923_ & new_n1486_;
  assign new_n1488_ = ~pc4 & new_n1486_;
  assign new_n1489_ = ~new_n1475_ & ~new_n1487_;
  assign new_n1490_ = ~new_n1488_ & new_n1489_;
  assign px9 = pz | new_n1490_;
  assign new_n1492_ = new_n912_ & ~new_n1026_;
  assign new_n1493_ = ~new_n912_ & ~new_n1038_;
  assign new_n1494_ = ~new_n1026_ & ~new_n1038_;
  assign new_n1495_ = ~new_n1492_ & ~new_n1493_;
  assign new_n1496_ = ~new_n1494_ & new_n1495_;
  assign new_n1497_ = ~new_n775_ & new_n1496_;
  assign new_n1498_ = ~pr3 & ~new_n1497_;
  assign new_n1499_ = pr3 & new_n1497_;
  assign new_n1500_ = ~new_n1498_ & ~new_n1499_;
  assign py8 = new_n738_ & new_n1500_;
  assign new_n1502_ = ~new_n874_ & new_n880_;
  assign new_n1503_ = ~pv4 & ~new_n1502_;
  assign new_n1504_ = pv4 & new_n1502_;
  assign new_n1505_ = ~new_n1503_ & ~new_n1504_;
  assign pc10 = new_n1350_ & new_n1505_;
  assign new_n1507_ = ~pm1 & ~new_n1442_;
  assign new_n1508_ = ~new_n316_ & new_n1507_;
  assign new_n1509_ = new_n323_ & new_n1507_;
  assign new_n1510_ = ~pn1 & ~new_n1442_;
  assign new_n1511_ = new_n323_ & new_n1510_;
  assign new_n1512_ = ~pc3 & ~pe3;
  assign new_n1513_ = ~pb3 & ~pd3;
  assign new_n1514_ = new_n1512_ & new_n1513_;
  assign new_n1515_ = ~pa3 & ~pz2;
  assign new_n1516_ = py2 & new_n1515_;
  assign new_n1517_ = new_n1514_ & new_n1516_;
  assign new_n1518_ = new_n1510_ & new_n1517_;
  assign new_n1519_ = ~new_n316_ & new_n1510_;
  assign new_n1520_ = new_n1507_ & new_n1517_;
  assign new_n1521_ = ~new_n1508_ & ~new_n1509_;
  assign new_n1522_ = ~new_n1511_ & new_n1521_;
  assign new_n1523_ = ~new_n1518_ & ~new_n1519_;
  assign new_n1524_ = ~new_n1520_ & new_n1523_;
  assign new_n1525_ = new_n1522_ & new_n1524_;
  assign new_n1526_ = new_n316_ & new_n1517_;
  assign new_n1527_ = ~pd1 & ~new_n1245_;
  assign new_n1528_ = ~pc & new_n1527_;
  assign new_n1529_ = pr1 & ~new_n1245_;
  assign new_n1530_ = ~pc & new_n1529_;
  assign new_n1531_ = ~pd1 & ~pr1;
  assign new_n1532_ = ~pc & new_n1531_;
  assign new_n1533_ = ~new_n1528_ & ~new_n1530_;
  assign new_n1534_ = ~new_n1532_ & new_n1533_;
  assign new_n1535_ = pv6 & new_n1534_;
  assign new_n1536_ = ~new_n1526_ & ~new_n1535_;
  assign new_n1537_ = ~new_n426_ & ~new_n1437_;
  assign new_n1538_ = new_n1536_ & new_n1537_;
  assign new_n1539_ = ~new_n1525_ & new_n1538_;
  assign pt6 = ~pb & ~new_n1539_;
  assign new_n1541_ = ~pb & ~new_n1066_;
  assign new_n1542_ = pj2 & pi2;
  assign new_n1543_ = pk2 & new_n1542_;
  assign new_n1544_ = pf2 & ph2;
  assign new_n1545_ = pl2 & pm2;
  assign new_n1546_ = po2 & new_n1545_;
  assign new_n1547_ = ~new_n1541_ & new_n1543_;
  assign new_n1548_ = new_n1544_ & new_n1547_;
  assign pu7 = new_n1546_ & new_n1548_;
  assign new_n1550_ = pp & pq1;
  assign new_n1551_ = pr & pn1;
  assign new_n1552_ = pq & ~new_n427_;
  assign new_n1553_ = ps & new_n1065_;
  assign new_n1554_ = ~new_n1550_ & ~new_n1551_;
  assign new_n1555_ = ~new_n1552_ & ~new_n1553_;
  assign new_n1556_ = new_n1554_ & new_n1555_;
  assign new_n1557_ = pw2 & pn;
  assign new_n1558_ = pm & new_n1517_;
  assign new_n1559_ = pc3 & pd3;
  assign new_n1560_ = pe3 & new_n1559_;
  assign new_n1561_ = po & new_n1560_;
  assign new_n1562_ = ~new_n1557_ & ~new_n1558_;
  assign new_n1563_ = ~new_n1561_ & new_n1562_;
  assign new_n1564_ = pt & pe2;
  assign new_n1565_ = pv & pz0;
  assign new_n1566_ = pu & new_n441_;
  assign new_n1567_ = pw & pl1;
  assign new_n1568_ = ~new_n1564_ & ~new_n1565_;
  assign new_n1569_ = ~new_n1566_ & ~new_n1567_;
  assign new_n1570_ = new_n1568_ & new_n1569_;
  assign new_n1571_ = new_n1556_ & new_n1563_;
  assign pw5 = ~new_n1570_ | ~new_n1571_;
  assign new_n1573_ = ~pr3 & new_n1026_;
  assign new_n1574_ = new_n912_ & ~new_n1573_;
  assign new_n1575_ = ~new_n912_ & ~new_n1039_;
  assign new_n1576_ = ~new_n1039_ & ~new_n1573_;
  assign new_n1577_ = ~new_n1574_ & ~new_n1575_;
  assign new_n1578_ = ~new_n1576_ & new_n1577_;
  assign new_n1579_ = ~new_n775_ & new_n1578_;
  assign new_n1580_ = ~ps3 & new_n1579_;
  assign new_n1581_ = ps3 & ~new_n1579_;
  assign new_n1582_ = ~new_n1580_ & ~new_n1581_;
  assign new_n1583_ = new_n738_ & ~new_n1582_;
  assign pz8 = new_n1015_ | new_n1583_;
  assign new_n1585_ = pt4 & new_n1351_;
  assign new_n1586_ = pr4 & new_n1585_;
  assign new_n1587_ = ~pu4 & ~new_n1586_;
  assign new_n1588_ = pu4 & new_n1586_;
  assign new_n1589_ = ~new_n1587_ & ~new_n1588_;
  assign pb10 = new_n1350_ & new_n1589_;
  assign new_n1591_ = ~pm2 & new_n1425_;
  assign new_n1592_ = pm2 & ~new_n1425_;
  assign new_n1593_ = ~new_n1591_ & ~new_n1592_;
  assign new_n1594_ = ~pz1 & new_n1593_;
  assign new_n1595_ = new_n1066_ & new_n1593_;
  assign new_n1596_ = ~pz1 & ~new_n1066_;
  assign new_n1597_ = ~new_n1594_ & ~new_n1595_;
  assign new_n1598_ = ~new_n1596_ & new_n1597_;
  assign pt7 = pb | new_n1598_;
  assign new_n1600_ = ~new_n1442_ & ~new_n1560_;
  assign new_n1601_ = ~new_n323_ & ~new_n1442_;
  assign new_n1602_ = ~new_n1442_ & new_n1517_;
  assign new_n1603_ = ~new_n316_ & ~new_n1442_;
  assign new_n1604_ = ~new_n1600_ & ~new_n1601_;
  assign new_n1605_ = ~new_n1602_ & ~new_n1603_;
  assign new_n1606_ = new_n1604_ & new_n1605_;
  assign new_n1607_ = ~new_n410_ & ~new_n1437_;
  assign new_n1608_ = ~new_n1517_ & new_n1607_;
  assign new_n1609_ = ~new_n316_ & new_n1607_;
  assign new_n1610_ = ~new_n1608_ & ~new_n1609_;
  assign new_n1611_ = ~new_n1606_ & ~new_n1610_;
  assign pu6 = ~pb & ~new_n1611_;
  assign new_n1613_ = pp & pp1;
  assign new_n1614_ = pr & pm1;
  assign new_n1615_ = pq & pr1;
  assign new_n1616_ = ps & pk2;
  assign new_n1617_ = ~new_n1613_ & ~new_n1614_;
  assign new_n1618_ = ~new_n1615_ & ~new_n1616_;
  assign new_n1619_ = new_n1617_ & new_n1618_;
  assign new_n1620_ = px2 & pn;
  assign new_n1621_ = pb3 & pm;
  assign new_n1622_ = pq2 & po;
  assign new_n1623_ = ~new_n1620_ & ~new_n1621_;
  assign new_n1624_ = ~new_n1622_ & new_n1623_;
  assign new_n1625_ = pf2 & pt;
  assign new_n1626_ = pa1 & pv;
  assign new_n1627_ = pb2 & pu;
  assign new_n1628_ = pw & pv0;
  assign new_n1629_ = ~new_n1625_ & ~new_n1626_;
  assign new_n1630_ = ~new_n1627_ & ~new_n1628_;
  assign new_n1631_ = new_n1629_ & new_n1630_;
  assign new_n1632_ = new_n1619_ & new_n1624_;
  assign pv5 = ~new_n1631_ | ~new_n1632_;
  assign new_n1634_ = ~ps4 & ~new_n1396_;
  assign new_n1635_ = ps4 & new_n1396_;
  assign new_n1636_ = ~new_n1634_ & ~new_n1635_;
  assign pz9 = new_n1350_ & new_n1636_;
  assign new_n1638_ = pv4 & ~new_n874_;
  assign new_n1639_ = pw4 & new_n1638_;
  assign new_n1640_ = new_n880_ & new_n1639_;
  assign new_n1641_ = ~px4 & ~new_n1640_;
  assign new_n1642_ = px4 & new_n1640_;
  assign new_n1643_ = ~new_n1641_ & ~new_n1642_;
  assign pe10 = new_n1350_ & new_n1643_;
  assign new_n1645_ = ~pl2 & new_n1424_;
  assign new_n1646_ = pl2 & ~new_n1424_;
  assign new_n1647_ = ~new_n1645_ & ~new_n1646_;
  assign new_n1648_ = ~py1 & new_n1647_;
  assign new_n1649_ = new_n1066_ & new_n1647_;
  assign new_n1650_ = ~py1 & ~new_n1066_;
  assign new_n1651_ = ~new_n1648_ & ~new_n1649_;
  assign new_n1652_ = ~new_n1650_ & new_n1651_;
  assign ps7 = pb | new_n1652_;
  assign new_n1654_ = new_n880_ & new_n1638_;
  assign new_n1655_ = ~pw4 & ~new_n1654_;
  assign new_n1656_ = pw4 & new_n1654_;
  assign new_n1657_ = ~new_n1655_ & ~new_n1656_;
  assign pd10 = new_n1350_ & new_n1657_;
  assign new_n1659_ = ~pk2 & ~new_n1423_;
  assign new_n1660_ = pk2 & new_n1423_;
  assign new_n1661_ = ~new_n1659_ & ~new_n1660_;
  assign new_n1662_ = ~px1 & new_n1661_;
  assign new_n1663_ = new_n1066_ & new_n1661_;
  assign new_n1664_ = ~px1 & ~new_n1066_;
  assign new_n1665_ = ~new_n1662_ & ~new_n1663_;
  assign new_n1666_ = ~new_n1664_ & new_n1665_;
  assign pr7 = pb | new_n1666_;
  assign new_n1668_ = new_n323_ & new_n426_;
  assign new_n1669_ = new_n323_ & new_n1560_;
  assign new_n1670_ = ~new_n1517_ & new_n1669_;
  assign new_n1671_ = new_n316_ & ~new_n1670_;
  assign new_n1672_ = ~new_n410_ & ~new_n1668_;
  assign new_n1673_ = ~new_n1671_ & new_n1672_;
  assign ps6 = ~pb & ~new_n1673_;
  assign new_n1675_ = ~pz4 & ~new_n882_;
  assign new_n1676_ = ~new_n883_ & ~new_n1675_;
  assign pg10 = new_n1350_ & new_n1676_;
  assign new_n1678_ = ~pi1 & new_n1102_;
  assign new_n1679_ = ~new_n322_ & new_n1102_;
  assign new_n1680_ = ~new_n1678_ & ~new_n1679_;
  assign new_n1681_ = pi1 & ~new_n1680_;
  assign pp6 = new_n335_ | new_n1681_;
  assign new_n1683_ = ~pj2 & new_n1421_;
  assign new_n1684_ = pj2 & ~new_n1421_;
  assign new_n1685_ = ~new_n1683_ & ~new_n1684_;
  assign new_n1686_ = ~pw1 & new_n1685_;
  assign new_n1687_ = new_n1066_ & new_n1685_;
  assign new_n1688_ = ~pw1 & ~new_n1066_;
  assign new_n1689_ = ~new_n1686_ & ~new_n1687_;
  assign new_n1690_ = ~new_n1688_ & new_n1689_;
  assign pq7 = pb | new_n1690_;
  assign new_n1692_ = pp & pa2;
  assign new_n1693_ = pr & pu1;
  assign new_n1694_ = pq & px1;
  assign new_n1695_ = ps & po2;
  assign new_n1696_ = ~new_n1692_ & ~new_n1693_;
  assign new_n1697_ = ~new_n1694_ & ~new_n1695_;
  assign new_n1698_ = new_n1696_ & new_n1697_;
  assign new_n1699_ = pa3 & pn;
  assign new_n1700_ = pe3 & pm;
  assign new_n1701_ = pt2 & po;
  assign new_n1702_ = ~new_n1699_ & ~new_n1700_;
  assign new_n1703_ = ~new_n1701_ & new_n1702_;
  assign new_n1704_ = pt & pj2;
  assign new_n1705_ = pd1 & pv;
  assign new_n1706_ = pg2 & pu;
  assign new_n1707_ = pw & py0;
  assign new_n1708_ = ~new_n1704_ & ~new_n1705_;
  assign new_n1709_ = ~new_n1706_ & ~new_n1707_;
  assign new_n1710_ = new_n1708_ & new_n1709_;
  assign new_n1711_ = new_n1698_ & new_n1703_;
  assign ps5 = ~new_n1710_ | ~new_n1711_;
  assign new_n1713_ = ~new_n874_ & new_n877_;
  assign new_n1714_ = new_n880_ & new_n1713_;
  assign new_n1715_ = ~py4 & ~new_n1714_;
  assign new_n1716_ = py4 & new_n1714_;
  assign new_n1717_ = ~new_n1715_ & ~new_n1716_;
  assign pf10 = new_n1350_ & new_n1717_;
  assign new_n1719_ = ~pi2 & new_n1420_;
  assign new_n1720_ = pi2 & ~new_n1420_;
  assign new_n1721_ = ~new_n1719_ & ~new_n1720_;
  assign new_n1722_ = ~pv1 & new_n1721_;
  assign new_n1723_ = new_n1066_ & new_n1721_;
  assign new_n1724_ = ~pv1 & ~new_n1066_;
  assign new_n1725_ = ~new_n1722_ & ~new_n1723_;
  assign new_n1726_ = ~new_n1724_ & new_n1725_;
  assign pp7 = pb | new_n1726_;
  assign new_n1728_ = ~new_n313_ & ~new_n410_;
  assign new_n1729_ = ~pj1 & ~new_n1065_;
  assign new_n1730_ = ~new_n1378_ & ~new_n1729_;
  assign new_n1731_ = ~pb & new_n1730_;
  assign pq6 = ~new_n1728_ | new_n1731_;
  assign new_n1733_ = ~new_n912_ & new_n1032_;
  assign new_n1734_ = new_n912_ & new_n1020_;
  assign new_n1735_ = ~new_n1733_ & ~new_n1734_;
  assign new_n1736_ = ~new_n775_ & ~new_n1735_;
  assign new_n1737_ = ~pi3 & new_n1736_;
  assign new_n1738_ = pi3 & ~new_n1736_;
  assign new_n1739_ = ~new_n1737_ & ~new_n1738_;
  assign new_n1740_ = new_n738_ & ~new_n1739_;
  assign pp8 = new_n1015_ | new_n1740_;
  assign new_n1742_ = ~pw3 & ~new_n923_;
  assign new_n1743_ = ~pj4 & new_n1476_;
  assign new_n1744_ = pj4 & ~new_n1476_;
  assign new_n1745_ = ~new_n1743_ & ~new_n1744_;
  assign new_n1746_ = new_n923_ & new_n1745_;
  assign new_n1747_ = ~pw3 & new_n1745_;
  assign new_n1748_ = ~new_n1742_ & ~new_n1746_;
  assign new_n1749_ = ~new_n1747_ & new_n1748_;
  assign pq9 = pz | new_n1749_;
  assign new_n1751_ = ~pi4 & new_n744_;
  assign new_n1752_ = ~new_n745_ & ~new_n1751_;
  assign pp9 = pz | new_n1752_;
  assign new_n1754_ = ~po3 & ~pm3;
  assign new_n1755_ = ~pn3 & ~pl3;
  assign new_n1756_ = new_n1754_ & new_n1755_;
  assign new_n1757_ = new_n738_ & new_n1756_;
  assign new_n1758_ = ~new_n738_ & new_n912_;
  assign new_n1759_ = new_n912_ & new_n1756_;
  assign new_n1760_ = ~new_n1757_ & ~new_n1758_;
  assign pq8 = new_n1759_ | ~new_n1760_;
  assign new_n1762_ = ~pz & ~new_n922_;
  assign new_n1763_ = ~new_n520_ & new_n1762_;
  assign new_n1764_ = ~pd5 & new_n1762_;
  assign new_n1765_ = ~new_n1763_ & ~new_n1764_;
  assign new_n1766_ = pd5 & ~new_n1765_;
  assign pk10 = new_n764_ | new_n1766_;
  assign new_n1768_ = po3 & pm3;
  assign new_n1769_ = pn3 & pl3;
  assign new_n1770_ = new_n1768_ & new_n1769_;
  assign pr8 = new_n738_ & new_n1770_;
  assign new_n1772_ = ~py3 & ~new_n923_;
  assign new_n1773_ = ~pl4 & new_n1478_;
  assign new_n1774_ = pl4 & ~new_n1478_;
  assign new_n1775_ = ~new_n1773_ & ~new_n1774_;
  assign new_n1776_ = new_n923_ & new_n1775_;
  assign new_n1777_ = ~py3 & new_n1775_;
  assign new_n1778_ = ~new_n1772_ & ~new_n1776_;
  assign new_n1779_ = ~new_n1777_ & new_n1778_;
  assign ps9 = pz | new_n1779_;
  assign new_n1781_ = ~px3 & ~new_n923_;
  assign new_n1782_ = ~pk4 & new_n1477_;
  assign new_n1783_ = pk4 & ~new_n1477_;
  assign new_n1784_ = ~new_n1782_ & ~new_n1783_;
  assign new_n1785_ = new_n923_ & new_n1784_;
  assign new_n1786_ = ~px3 & new_n1784_;
  assign new_n1787_ = ~new_n1781_ & ~new_n1785_;
  assign new_n1788_ = ~new_n1786_ & new_n1787_;
  assign pr9 = pz | new_n1788_;
  assign new_n1790_ = new_n912_ & new_n1022_;
  assign new_n1791_ = ~new_n912_ & new_n1034_;
  assign new_n1792_ = new_n1022_ & new_n1034_;
  assign new_n1793_ = ~new_n1790_ & ~new_n1791_;
  assign new_n1794_ = ~new_n1792_ & new_n1793_;
  assign new_n1795_ = ~new_n775_ & new_n1794_;
  assign new_n1796_ = ~pl3 & ~new_n1795_;
  assign new_n1797_ = pl3 & new_n1795_;
  assign new_n1798_ = ~new_n1796_ & ~new_n1797_;
  assign ps8 = new_n738_ & new_n1798_;
  assign new_n1800_ = ~new_n475_ & ~new_n922_;
  assign new_n1801_ = ~pg5 & ~pf5;
  assign new_n1802_ = ~pf5 & ~new_n1801_;
  assign new_n1803_ = ~pz & new_n1802_;
  assign new_n1804_ = ~ph5 & ~new_n748_;
  assign new_n1805_ = ph5 & new_n748_;
  assign new_n1806_ = ~new_n1804_ & ~new_n1805_;
  assign new_n1807_ = ~pz & new_n1806_;
  assign po10 = ~new_n1800_ | new_n1807_;
  assign new_n1809_ = ~ph5 & po10;
  assign new_n1810_ = ~new_n1801_ & new_n1809_;
  assign new_n1811_ = ~pz & new_n1810_;
  assign new_n1812_ = ~pf5 & ~new_n1809_;
  assign new_n1813_ = ~pz & new_n1812_;
  assign new_n1814_ = ~new_n1803_ & ~new_n1811_;
  assign new_n1815_ = ~new_n1813_ & new_n1814_;
  assign pm10 = new_n1800_ & new_n1815_;
  assign new_n1817_ = ~pl3 & ~new_n1022_;
  assign new_n1818_ = new_n912_ & ~new_n1817_;
  assign new_n1819_ = pl3 & ~new_n1034_;
  assign new_n1820_ = ~new_n912_ & ~new_n1819_;
  assign new_n1821_ = ~new_n1817_ & ~new_n1819_;
  assign new_n1822_ = ~new_n1818_ & ~new_n1820_;
  assign new_n1823_ = ~new_n1821_ & new_n1822_;
  assign new_n1824_ = ~new_n775_ & new_n1823_;
  assign new_n1825_ = ~pm3 & ~new_n1824_;
  assign new_n1826_ = pm3 & new_n1824_;
  assign new_n1827_ = ~new_n1825_ & ~new_n1826_;
  assign pt8 = new_n738_ & new_n1827_;
  assign new_n1829_ = ~pa4 & ~new_n923_;
  assign new_n1830_ = ~pn4 & new_n1481_;
  assign new_n1831_ = pn4 & ~new_n1481_;
  assign new_n1832_ = ~new_n1830_ & ~new_n1831_;
  assign new_n1833_ = new_n923_ & new_n1832_;
  assign new_n1834_ = ~pa4 & new_n1832_;
  assign new_n1835_ = ~new_n1829_ & ~new_n1833_;
  assign new_n1836_ = ~new_n1834_ & new_n1835_;
  assign pu9 = pz | new_n1836_;
  assign new_n1838_ = pb4 & pn0;
  assign new_n1839_ = pp0 & pv3;
  assign new_n1840_ = po0 & py3;
  assign new_n1841_ = po4 & pq0;
  assign new_n1842_ = ~new_n1838_ & ~new_n1839_;
  assign new_n1843_ = ~new_n1840_ & ~new_n1841_;
  assign new_n1844_ = new_n1842_ & new_n1843_;
  assign new_n1845_ = pl0 & po3;
  assign new_n1846_ = pk0 & ps3;
  assign new_n1847_ = ph3 & pm0;
  assign new_n1848_ = ~new_n1845_ & ~new_n1846_;
  assign new_n1849_ = ~new_n1847_ & new_n1848_;
  assign new_n1850_ = pk4 & pr0;
  assign new_n1851_ = pt0 & py4;
  assign new_n1852_ = pf4 & ps0;
  assign new_n1853_ = pt4 & pu0;
  assign new_n1854_ = ~new_n1850_ & ~new_n1851_;
  assign new_n1855_ = ~new_n1852_ & ~new_n1853_;
  assign new_n1856_ = new_n1854_ & new_n1855_;
  assign new_n1857_ = new_n1844_ & new_n1849_;
  assign py5 = ~new_n1856_ | ~new_n1857_;
  assign new_n1859_ = ~ps1 & ~new_n381_;
  assign new_n1860_ = ps1 & new_n381_;
  assign new_n1861_ = ~new_n1859_ & ~new_n1860_;
  assign new_n1862_ = ~pw2 & new_n1861_;
  assign new_n1863_ = ~new_n416_ & new_n1861_;
  assign new_n1864_ = ~pw2 & new_n416_;
  assign new_n1865_ = ~new_n1862_ & ~new_n1863_;
  assign new_n1866_ = ~new_n1864_ & new_n1865_;
  assign pz6 = ~pb & new_n1866_;
  assign new_n1868_ = ~pe5 & new_n1762_;
  assign new_n1869_ = ~new_n519_ & new_n1762_;
  assign new_n1870_ = ~new_n1868_ & ~new_n1869_;
  assign new_n1871_ = pe5 & ~new_n1870_;
  assign pl10 = new_n526_ | new_n1871_;
  assign new_n1873_ = ~pz3 & ~new_n923_;
  assign new_n1874_ = ~pm4 & ~new_n1480_;
  assign new_n1875_ = pm4 & new_n1480_;
  assign new_n1876_ = ~new_n1874_ & ~new_n1875_;
  assign new_n1877_ = new_n923_ & new_n1876_;
  assign new_n1878_ = ~pz3 & new_n1876_;
  assign new_n1879_ = ~new_n1873_ & ~new_n1877_;
  assign new_n1880_ = ~new_n1878_ & new_n1879_;
  assign pt9 = pz | new_n1880_;
  assign new_n1882_ = ~pm3 & ~pl3;
  assign new_n1883_ = ~new_n1022_ & new_n1882_;
  assign new_n1884_ = new_n912_ & ~new_n1883_;
  assign new_n1885_ = pm3 & new_n1819_;
  assign new_n1886_ = ~new_n912_ & ~new_n1885_;
  assign new_n1887_ = ~new_n1883_ & ~new_n1885_;
  assign new_n1888_ = ~new_n1884_ & ~new_n1886_;
  assign new_n1889_ = ~new_n1887_ & new_n1888_;
  assign new_n1890_ = ~new_n775_ & new_n1889_;
  assign new_n1891_ = ~pn3 & ~new_n1890_;
  assign new_n1892_ = pn3 & new_n1890_;
  assign new_n1893_ = ~new_n1891_ & ~new_n1892_;
  assign pu8 = new_n738_ & new_n1893_;
  assign new_n1895_ = pc4 & pn0;
  assign new_n1896_ = pp0 & pw3;
  assign new_n1897_ = po0 & pz3;
  assign new_n1898_ = pq0 & pq4;
  assign new_n1899_ = ~new_n1895_ & ~new_n1896_;
  assign new_n1900_ = ~new_n1897_ & ~new_n1898_;
  assign new_n1901_ = new_n1899_ & new_n1900_;
  assign new_n1902_ = pl0 & pp3;
  assign new_n1903_ = pk0 & pt3;
  assign new_n1904_ = pi3 & pm0;
  assign new_n1905_ = ~new_n1902_ & ~new_n1903_;
  assign new_n1906_ = ~new_n1904_ & new_n1905_;
  assign new_n1907_ = pl4 & pr0;
  assign new_n1908_ = pt0 & pz4;
  assign new_n1909_ = pi4 & ps0;
  assign new_n1910_ = pu4 & pu0;
  assign new_n1911_ = ~new_n1907_ & ~new_n1908_;
  assign new_n1912_ = ~new_n1909_ & ~new_n1910_;
  assign new_n1913_ = new_n1911_ & new_n1912_;
  assign new_n1914_ = new_n1901_ & new_n1906_;
  assign px5 = ~new_n1913_ | ~new_n1914_;
  assign new_n1916_ = ~new_n423_ & new_n447_;
  assign new_n1917_ = new_n447_ & new_n456_;
  assign new_n1918_ = new_n423_ & new_n456_;
  assign new_n1919_ = ~new_n1916_ & ~new_n1917_;
  assign new_n1920_ = ~new_n1918_ & new_n1919_;
  assign new_n1921_ = ~new_n441_ & new_n1920_;
  assign new_n1922_ = ~ps2 & ~new_n1921_;
  assign new_n1923_ = ps2 & new_n1921_;
  assign new_n1924_ = ~new_n1922_ & ~new_n1923_;
  assign pz7 = new_n427_ & new_n1924_;
  assign new_n1926_ = ~pm3 & new_n1755_;
  assign new_n1927_ = ~new_n1022_ & new_n1926_;
  assign new_n1928_ = new_n912_ & ~new_n1927_;
  assign new_n1929_ = pm3 & ~new_n1034_;
  assign new_n1930_ = pl3 & new_n1929_;
  assign new_n1931_ = pn3 & new_n1930_;
  assign new_n1932_ = ~new_n912_ & ~new_n1931_;
  assign new_n1933_ = ~new_n1927_ & ~new_n1931_;
  assign new_n1934_ = ~new_n1928_ & ~new_n1932_;
  assign new_n1935_ = ~new_n1933_ & new_n1934_;
  assign new_n1936_ = ~new_n775_ & new_n1935_;
  assign new_n1937_ = ~po3 & new_n1936_;
  assign new_n1938_ = po3 & ~new_n1936_;
  assign new_n1939_ = ~new_n1937_ & ~new_n1938_;
  assign new_n1940_ = new_n738_ & ~new_n1939_;
  assign pv8 = new_n1015_ | new_n1940_;
  assign new_n1942_ = ~pz & ~new_n923_;
  assign new_n1943_ = pl4 & pk4;
  assign new_n1944_ = pm4 & new_n1943_;
  assign new_n1945_ = ph4 & pj4;
  assign new_n1946_ = pn4 & po4;
  assign new_n1947_ = pq4 & new_n1946_;
  assign new_n1948_ = ~new_n1942_ & new_n1944_;
  assign new_n1949_ = new_n1945_ & new_n1948_;
  assign pw9 = new_n1947_ & new_n1949_;
  assign new_n1951_ = ~pq1 & new_n1438_;
  assign new_n1952_ = ~pp1 & new_n1951_;
  assign new_n1953_ = ~pq1 & new_n1444_;
  assign new_n1954_ = ~pr1 & new_n1443_;
  assign new_n1955_ = ~pq1 & new_n1954_;
  assign new_n1956_ = ~pp1 & new_n1448_;
  assign new_n1957_ = ~pr1 & new_n1452_;
  assign new_n1958_ = ~pp1 & new_n1454_;
  assign new_n1959_ = ~pp1 & new_n1456_;
  assign new_n1960_ = ~new_n1952_ & ~new_n1953_;
  assign new_n1961_ = ~new_n1955_ & ~new_n1956_;
  assign new_n1962_ = new_n1960_ & new_n1961_;
  assign new_n1963_ = ~new_n1958_ & ~new_n1959_;
  assign new_n1964_ = ~new_n1451_ & ~new_n1957_;
  assign new_n1965_ = new_n1963_ & new_n1964_;
  assign new_n1966_ = new_n1962_ & new_n1965_;
  assign px6 = ~new_n1473_ & new_n1966_;
  assign new_n1968_ = ~pq2 & ~new_n423_;
  assign new_n1969_ = pq2 & new_n423_;
  assign new_n1970_ = ~new_n1968_ & ~new_n1969_;
  assign new_n1971_ = ~new_n441_ & new_n1970_;
  assign new_n1972_ = ~pr2 & ~new_n1971_;
  assign new_n1973_ = pr2 & new_n1971_;
  assign new_n1974_ = ~new_n1972_ & ~new_n1973_;
  assign py7 = new_n427_ & new_n1974_;
  assign new_n1976_ = new_n1800_ & ~new_n1809_;
  assign new_n1977_ = ~pg5 & new_n1976_;
  assign new_n1978_ = new_n1800_ & new_n1809_;
  assign new_n1979_ = ~pf5 & new_n1978_;
  assign new_n1980_ = ~pg5 & new_n1800_;
  assign new_n1981_ = ~pf5 & new_n1980_;
  assign new_n1982_ = ~new_n1977_ & ~new_n1979_;
  assign new_n1983_ = ~new_n1981_ & new_n1982_;
  assign pn10 = ~pz & new_n1983_;
  assign new_n1985_ = ~pb4 & ~new_n923_;
  assign new_n1986_ = ~po4 & new_n1482_;
  assign new_n1987_ = po4 & ~new_n1482_;
  assign new_n1988_ = ~new_n1986_ & ~new_n1987_;
  assign new_n1989_ = new_n923_ & new_n1988_;
  assign new_n1990_ = ~pb4 & new_n1988_;
  assign new_n1991_ = ~new_n1985_ & ~new_n1989_;
  assign new_n1992_ = ~new_n1990_ & new_n1991_;
  assign pv9 = pz | new_n1992_;
  assign new_n1994_ = new_n912_ & ~new_n1023_;
  assign new_n1995_ = ~new_n912_ & ~new_n1035_;
  assign new_n1996_ = ~new_n1023_ & ~new_n1035_;
  assign new_n1997_ = ~new_n1994_ & ~new_n1995_;
  assign new_n1998_ = ~new_n1996_ & new_n1997_;
  assign new_n1999_ = ~new_n775_ & new_n1998_;
  assign new_n2000_ = ~pp3 & new_n1999_;
  assign new_n2001_ = pp3 & ~new_n1999_;
  assign new_n2002_ = ~new_n2000_ & ~new_n2001_;
  assign new_n2003_ = new_n738_ & ~new_n2002_;
  assign pw8 = new_n1015_ | new_n2003_;
  assign new_n2005_ = ~pq2 & new_n441_;
  assign new_n2006_ = pq2 & ~new_n441_;
  assign new_n2007_ = ~new_n2005_ & ~new_n2006_;
  assign px7 = new_n427_ & new_n2007_;
  assign new_n2009_ = ~pq1 & new_n1439_;
  assign new_n2010_ = ~pr1 & new_n1444_;
  assign new_n2011_ = ~pp1 & new_n1954_;
  assign new_n2012_ = ~pq1 & ~new_n1443_;
  assign new_n2013_ = ~pp1 & new_n2012_;
  assign new_n2014_ = ~pp1 & new_n1452_;
  assign new_n2015_ = ~pq1 & new_n1454_;
  assign new_n2016_ = ~pq1 & ~new_n1438_;
  assign new_n2017_ = ~pp1 & new_n2016_;
  assign new_n2018_ = ~new_n2009_ & ~new_n2010_;
  assign new_n2019_ = ~new_n2011_ & ~new_n2013_;
  assign new_n2020_ = new_n2018_ & new_n2019_;
  assign new_n2021_ = ~new_n2015_ & ~new_n2017_;
  assign new_n2022_ = ~new_n1451_ & ~new_n2014_;
  assign new_n2023_ = new_n2021_ & new_n2022_;
  assign new_n2024_ = new_n2020_ & new_n2023_;
  assign py6 = ~new_n1473_ & new_n2024_;
  assign new_n2026_ = pa4 & pn0;
  assign new_n2027_ = pp0 & pu3;
  assign new_n2028_ = po0 & px3;
  assign new_n2029_ = pn4 & pq0;
  assign new_n2030_ = ~new_n2026_ & ~new_n2027_;
  assign new_n2031_ = ~new_n2028_ & ~new_n2029_;
  assign new_n2032_ = new_n2030_ & new_n2031_;
  assign new_n2033_ = pl0 & pn3;
  assign new_n2034_ = pk0 & pr3;
  assign new_n2035_ = pg3 & pm0;
  assign new_n2036_ = ~new_n2033_ & ~new_n2034_;
  assign new_n2037_ = ~new_n2035_ & new_n2036_;
  assign new_n2038_ = pj4 & pr0;
  assign new_n2039_ = pt0 & px4;
  assign new_n2040_ = pe4 & ps0;
  assign new_n2041_ = pu0 & ps4;
  assign new_n2042_ = ~new_n2038_ & ~new_n2039_;
  assign new_n2043_ = ~new_n2040_ & ~new_n2041_;
  assign new_n2044_ = new_n2042_ & new_n2043_;
  assign new_n2045_ = new_n2032_ & new_n2037_;
  assign pz5 = ~new_n2044_ | ~new_n2045_;
  assign pp10 = pg5;
  assign pl6 = pa;
  assign pm6 = pe1;
  assign pr6 = pj1;
  assign pi10 = pa5;
  assign ph10 = py;
endmodule

