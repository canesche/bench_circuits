module top ( 
    i_50_, i_40_, i_30_, i_20_, i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_27_,
    i_14_, i_3_, i_39_, i_28_, i_13_, i_4_, i_25_, i_12_, i_1_, i_26_,
    i_11_, i_2_, i_49_, i_23_, i_18_, i_24_, i_17_, i_0_, i_21_, i_16_,
    i_22_, i_15_, i_45_, i_32_, i_46_, i_31_, i_47_, i_34_, i_48_, i_33_,
    i_19_, i_41_, i_36_, i_53_, i_42_, i_35_, i_52_, i_43_, i_38_, i_29_,
    i_51_, i_44_, i_37_,
    o_1_, o_19_, o_2_, o_0_, o_29_, o_39_, o_38_, o_25_, o_12_, o_37_,
    o_26_, o_11_, o_36_, o_27_, o_14_, o_35_, o_28_, o_13_, o_34_, o_21_,
    o_16_, o_40_, o_33_, o_22_, o_15_, o_32_, o_23_, o_18_, o_31_, o_24_,
    o_17_, o_43_, o_30_, o_44_, o_41_, o_42_, o_20_, o_47_, o_48_, o_45_,
    o_10_, o_46_, o_9_, o_49_, o_7_, o_8_, o_5_, o_6_, o_3_, o_4_  );
  input  i_50_, i_40_, i_30_, i_20_, i_9_, i_10_, i_7_, i_8_, i_5_, i_6_,
    i_27_, i_14_, i_3_, i_39_, i_28_, i_13_, i_4_, i_25_, i_12_, i_1_,
    i_26_, i_11_, i_2_, i_49_, i_23_, i_18_, i_24_, i_17_, i_0_, i_21_,
    i_16_, i_22_, i_15_, i_45_, i_32_, i_46_, i_31_, i_47_, i_34_, i_48_,
    i_33_, i_19_, i_41_, i_36_, i_53_, i_42_, i_35_, i_52_, i_43_, i_38_,
    i_29_, i_51_, i_44_, i_37_;
  output o_1_, o_19_, o_2_, o_0_, o_29_, o_39_, o_38_, o_25_, o_12_, o_37_,
    o_26_, o_11_, o_36_, o_27_, o_14_, o_35_, o_28_, o_13_, o_34_, o_21_,
    o_16_, o_40_, o_33_, o_22_, o_15_, o_32_, o_23_, o_18_, o_31_, o_24_,
    o_17_, o_43_, o_30_, o_44_, o_41_, o_42_, o_20_, o_47_, o_48_, o_45_,
    o_10_, o_46_, o_9_, o_49_, o_7_, o_8_, o_5_, o_6_, o_3_, o_4_;
  wire new_n105_, new_n106_, new_n107_, new_n108_, new_n109_, new_n110_,
    new_n111_, new_n112_, new_n113_, new_n114_, new_n115_, new_n116_,
    new_n117_, new_n118_, new_n119_, new_n120_, new_n121_, new_n122_,
    new_n123_, new_n124_, new_n125_, new_n126_, new_n127_, new_n128_,
    new_n129_, new_n130_, new_n131_, new_n132_, new_n133_, new_n134_,
    new_n135_, new_n136_, new_n137_, new_n138_, new_n139_, new_n140_,
    new_n141_, new_n142_, new_n143_, new_n144_, new_n145_, new_n146_,
    new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_,
    new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_,
    new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_,
    new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_,
    new_n171_, new_n172_, new_n173_, new_n174_, new_n175_, new_n176_,
    new_n177_, new_n178_, new_n179_, new_n180_, new_n181_, new_n182_,
    new_n183_, new_n184_, new_n185_, new_n186_, new_n187_, new_n188_,
    new_n189_, new_n190_, new_n191_, new_n192_, new_n193_, new_n194_,
    new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_,
    new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_,
    new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_,
    new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_,
    new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_,
    new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_,
    new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_,
    new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_,
    new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_,
    new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_,
    new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_,
    new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_,
    new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_,
    new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_,
    new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_,
    new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_,
    new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_,
    new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_,
    new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_,
    new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_,
    new_n339_, new_n340_, new_n341_, new_n342_, new_n343_, new_n344_,
    new_n345_, new_n346_, new_n347_, new_n348_, new_n349_, new_n350_,
    new_n351_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_,
    new_n357_, new_n358_, new_n359_, new_n360_, new_n361_, new_n362_,
    new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_,
    new_n369_, new_n370_, new_n371_, new_n372_, new_n373_, new_n374_,
    new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n380_,
    new_n381_, new_n382_, new_n383_, new_n384_, new_n385_, new_n386_,
    new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n392_,
    new_n393_, new_n394_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_,
    new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_,
    new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n456_,
    new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_,
    new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_,
    new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_,
    new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_,
    new_n481_, new_n482_, new_n483_, new_n484_, new_n486_, new_n487_,
    new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_,
    new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n500_,
    new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_,
    new_n507_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n791_, new_n792_, new_n793_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n804_, new_n805_, new_n807_, new_n808_, new_n809_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n854_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n919_,
    new_n920_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n939_, new_n940_, new_n941_, new_n942_,
    new_n943_, new_n944_, new_n945_, new_n946_, new_n947_, new_n948_,
    new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n961_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n968_, new_n969_, new_n971_,
    new_n972_, new_n973_, new_n974_, new_n975_, new_n977_, new_n978_,
    new_n981_, new_n982_, new_n983_, new_n984_, new_n985_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_,
    new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_,
    new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_,
    new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_,
    new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_,
    new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_,
    new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_,
    new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_,
    new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_,
    new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_,
    new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_,
    new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_,
    new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_,
    new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_,
    new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_,
    new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_,
    new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_,
    new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_,
    new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_,
    new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_,
    new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_,
    new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_,
    new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_,
    new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_,
    new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_,
    new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_,
    new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_,
    new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_,
    new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_,
    new_n1168_, new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_,
    new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_,
    new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_,
    new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_,
    new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_,
    new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_,
    new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_,
    new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_,
    new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_,
    new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_,
    new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_,
    new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_,
    new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_,
    new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_,
    new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_,
    new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_,
    new_n1266_, new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_,
    new_n1272_, new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_,
    new_n1278_, new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_,
    new_n1284_, new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_,
    new_n1290_, new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_,
    new_n1296_, new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_,
    new_n1302_, new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_,
    new_n1308_, new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_,
    new_n1314_, new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_,
    new_n1320_, new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_,
    new_n1326_, new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_,
    new_n1332_, new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_,
    new_n1338_, new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_,
    new_n1344_, new_n1345_, new_n1346_, new_n1348_, new_n1349_, new_n1350_,
    new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_,
    new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_,
    new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_,
    new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_,
    new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_,
    new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_,
    new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_,
    new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_, new_n1398_,
    new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_,
    new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_,
    new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_,
    new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_,
    new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_,
    new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_,
    new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_,
    new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_, new_n1446_,
    new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_, new_n1452_,
    new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_, new_n1458_,
    new_n1459_, new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1465_,
    new_n1466_, new_n1467_, new_n1468_, new_n1469_, new_n1470_, new_n1471_,
    new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_, new_n1477_,
    new_n1478_, new_n1479_, new_n1480_, new_n1481_, new_n1482_, new_n1483_,
    new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_, new_n1489_,
    new_n1490_, new_n1491_, new_n1492_, new_n1493_, new_n1494_, new_n1495_,
    new_n1496_, new_n1497_, new_n1498_, new_n1499_, new_n1500_, new_n1501_,
    new_n1502_, new_n1503_, new_n1504_, new_n1505_, new_n1506_, new_n1507_,
    new_n1508_, new_n1509_, new_n1510_, new_n1511_, new_n1512_, new_n1513_,
    new_n1514_, new_n1515_, new_n1516_, new_n1517_, new_n1518_, new_n1519_,
    new_n1520_, new_n1521_, new_n1522_, new_n1523_, new_n1524_, new_n1525_,
    new_n1526_, new_n1527_, new_n1528_, new_n1529_, new_n1530_, new_n1531_,
    new_n1532_, new_n1533_, new_n1534_, new_n1535_, new_n1536_, new_n1537_,
    new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1542_, new_n1543_,
    new_n1544_, new_n1545_, new_n1546_, new_n1547_, new_n1548_, new_n1549_,
    new_n1550_, new_n1551_, new_n1552_, new_n1553_, new_n1554_, new_n1555_,
    new_n1556_, new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1561_,
    new_n1562_, new_n1563_, new_n1564_, new_n1565_, new_n1566_, new_n1567_,
    new_n1568_, new_n1569_, new_n1570_, new_n1571_, new_n1572_, new_n1573_,
    new_n1574_, new_n1575_, new_n1576_, new_n1577_, new_n1578_, new_n1579_,
    new_n1580_, new_n1581_, new_n1583_, new_n1584_, new_n1585_, new_n1586_,
    new_n1587_, new_n1588_, new_n1589_, new_n1590_, new_n1591_, new_n1592_,
    new_n1593_, new_n1594_, new_n1595_, new_n1596_, new_n1597_, new_n1598_,
    new_n1599_, new_n1600_, new_n1601_, new_n1602_, new_n1603_, new_n1604_,
    new_n1605_, new_n1606_, new_n1607_, new_n1608_, new_n1609_, new_n1610_,
    new_n1611_, new_n1612_, new_n1613_, new_n1614_, new_n1615_, new_n1616_,
    new_n1617_, new_n1618_, new_n1619_, new_n1620_, new_n1621_, new_n1622_,
    new_n1623_, new_n1624_, new_n1625_, new_n1626_, new_n1627_, new_n1628_,
    new_n1629_, new_n1630_, new_n1631_, new_n1632_, new_n1633_, new_n1634_,
    new_n1635_, new_n1636_, new_n1637_, new_n1638_, new_n1639_, new_n1640_,
    new_n1641_, new_n1642_, new_n1643_, new_n1644_, new_n1645_, new_n1646_,
    new_n1647_, new_n1648_, new_n1649_, new_n1650_, new_n1651_, new_n1652_,
    new_n1653_, new_n1654_, new_n1655_, new_n1656_, new_n1657_, new_n1658_,
    new_n1659_, new_n1660_, new_n1661_, new_n1662_, new_n1663_, new_n1664_,
    new_n1665_, new_n1666_, new_n1667_, new_n1668_, new_n1669_, new_n1670_,
    new_n1671_, new_n1672_, new_n1673_, new_n1674_, new_n1675_, new_n1676_,
    new_n1677_, new_n1678_, new_n1679_, new_n1680_, new_n1681_, new_n1682_,
    new_n1683_, new_n1684_, new_n1685_, new_n1686_, new_n1687_, new_n1688_,
    new_n1689_, new_n1690_, new_n1691_, new_n1692_, new_n1693_, new_n1694_,
    new_n1695_, new_n1696_, new_n1697_, new_n1698_, new_n1699_, new_n1700_,
    new_n1701_, new_n1702_, new_n1703_, new_n1704_, new_n1705_, new_n1706_;
  assign new_n105_ = ~i_50_ & i_51_;
  assign new_n106_ = ~i_49_ & new_n105_;
  assign new_n107_ = ~i_53_ & ~i_52_;
  assign new_n108_ = i_46_ & ~i_47_;
  assign new_n109_ = i_37_ & new_n108_;
  assign new_n110_ = new_n106_ & new_n107_;
  assign new_n111_ = new_n109_ & new_n110_;
  assign new_n112_ = i_50_ & ~i_49_;
  assign new_n113_ = i_48_ & new_n112_;
  assign new_n114_ = ~i_51_ & new_n107_;
  assign new_n115_ = i_4_ & new_n108_;
  assign new_n116_ = new_n113_ & new_n114_;
  assign new_n117_ = new_n115_ & new_n116_;
  assign new_n118_ = i_50_ & i_51_;
  assign new_n119_ = ~i_49_ & new_n118_;
  assign new_n120_ = i_53_ & ~i_52_;
  assign new_n121_ = ~i_47_ & i_48_;
  assign new_n122_ = i_46_ & new_n121_;
  assign new_n123_ = new_n119_ & new_n120_;
  assign new_n124_ = new_n122_ & new_n123_;
  assign new_n125_ = ~new_n111_ & ~new_n117_;
  assign new_n126_ = ~new_n124_ & new_n125_;
  assign new_n127_ = i_53_ & i_52_;
  assign new_n128_ = i_47_ & ~i_48_;
  assign new_n129_ = ~i_46_ & new_n128_;
  assign new_n130_ = new_n119_ & new_n127_;
  assign new_n131_ = new_n129_ & new_n130_;
  assign new_n132_ = i_49_ & new_n105_;
  assign new_n133_ = ~i_46_ & i_47_;
  assign new_n134_ = i_20_ & new_n133_;
  assign new_n135_ = ~i_52_ & new_n132_;
  assign new_n136_ = new_n134_ & new_n135_;
  assign new_n137_ = ~i_48_ & new_n112_;
  assign new_n138_ = ~i_53_ & ~i_51_;
  assign new_n139_ = ~i_28_ & new_n133_;
  assign new_n140_ = new_n137_ & new_n138_;
  assign new_n141_ = new_n139_ & new_n140_;
  assign new_n142_ = ~new_n131_ & ~new_n136_;
  assign new_n143_ = ~new_n141_ & new_n142_;
  assign new_n144_ = ~i_50_ & i_49_;
  assign new_n145_ = i_48_ & new_n144_;
  assign new_n146_ = ~i_53_ & i_51_;
  assign new_n147_ = i_1_ & new_n133_;
  assign new_n148_ = new_n145_ & new_n146_;
  assign new_n149_ = new_n147_ & new_n148_;
  assign new_n150_ = ~i_43_ & new_n133_;
  assign new_n151_ = new_n148_ & new_n150_;
  assign new_n152_ = ~i_50_ & ~i_51_;
  assign new_n153_ = ~i_49_ & new_n152_;
  assign new_n154_ = i_47_ & i_48_;
  assign new_n155_ = ~i_46_ & new_n154_;
  assign new_n156_ = new_n127_ & new_n153_;
  assign new_n157_ = new_n155_ & new_n156_;
  assign new_n158_ = ~new_n149_ & ~new_n151_;
  assign new_n159_ = ~new_n157_ & new_n158_;
  assign new_n160_ = new_n126_ & new_n143_;
  assign new_n161_ = new_n159_ & new_n160_;
  assign new_n162_ = ~i_53_ & i_52_;
  assign new_n163_ = i_51_ & new_n162_;
  assign new_n164_ = i_3_ & new_n108_;
  assign new_n165_ = new_n113_ & new_n163_;
  assign new_n166_ = new_n164_ & new_n165_;
  assign new_n167_ = ~i_50_ & ~i_49_;
  assign new_n168_ = i_48_ & new_n167_;
  assign new_n169_ = new_n114_ & new_n168_;
  assign new_n170_ = new_n147_ & new_n169_;
  assign new_n171_ = i_50_ & i_49_;
  assign new_n172_ = ~i_48_ & new_n171_;
  assign new_n173_ = ~i_51_ & new_n127_;
  assign new_n174_ = new_n172_ & new_n173_;
  assign new_n175_ = new_n147_ & new_n174_;
  assign new_n176_ = ~new_n166_ & ~new_n170_;
  assign new_n177_ = ~new_n175_ & new_n176_;
  assign new_n178_ = ~i_51_ & new_n120_;
  assign new_n179_ = ~i_1_ & new_n133_;
  assign new_n180_ = new_n168_ & new_n178_;
  assign new_n181_ = new_n179_ & new_n180_;
  assign new_n182_ = i_49_ & i_48_;
  assign new_n183_ = i_47_ & new_n182_;
  assign new_n184_ = ~i_52_ & i_51_;
  assign new_n185_ = ~i_46_ & i_43_;
  assign new_n186_ = ~i_1_ & new_n185_;
  assign new_n187_ = new_n183_ & new_n184_;
  assign new_n188_ = new_n186_ & new_n187_;
  assign new_n189_ = new_n150_ & new_n180_;
  assign new_n190_ = ~new_n181_ & ~new_n188_;
  assign new_n191_ = ~new_n189_ & new_n190_;
  assign new_n192_ = ~i_48_ & new_n105_;
  assign new_n193_ = ~i_29_ & new_n133_;
  assign new_n194_ = new_n120_ & new_n192_;
  assign new_n195_ = new_n193_ & new_n194_;
  assign new_n196_ = i_51_ & new_n120_;
  assign new_n197_ = i_43_ & new_n133_;
  assign new_n198_ = new_n172_ & new_n196_;
  assign new_n199_ = new_n197_ & new_n198_;
  assign new_n200_ = ~i_50_ & i_52_;
  assign new_n201_ = ~i_49_ & new_n200_;
  assign new_n202_ = ~i_13_ & new_n133_;
  assign new_n203_ = i_53_ & new_n201_;
  assign new_n204_ = new_n202_ & new_n203_;
  assign new_n205_ = ~new_n195_ & ~new_n199_;
  assign new_n206_ = ~new_n204_ & new_n205_;
  assign new_n207_ = new_n177_ & new_n191_;
  assign new_n208_ = new_n206_ & new_n207_;
  assign new_n209_ = ~i_51_ & new_n162_;
  assign new_n210_ = i_16_ & new_n108_;
  assign new_n211_ = new_n168_ & new_n209_;
  assign new_n212_ = new_n210_ & new_n211_;
  assign new_n213_ = ~i_48_ & new_n167_;
  assign new_n214_ = i_51_ & new_n127_;
  assign new_n215_ = i_39_ & new_n108_;
  assign new_n216_ = new_n213_ & new_n214_;
  assign new_n217_ = new_n215_ & new_n216_;
  assign new_n218_ = ~i_49_ & ~i_51_;
  assign new_n219_ = i_48_ & new_n218_;
  assign new_n220_ = ~i_53_ & new_n219_;
  assign new_n221_ = new_n179_ & new_n220_;
  assign new_n222_ = ~new_n212_ & ~new_n217_;
  assign new_n223_ = ~new_n221_ & new_n222_;
  assign new_n224_ = ~i_48_ & new_n144_;
  assign new_n225_ = i_52_ & ~i_51_;
  assign new_n226_ = i_38_ & new_n133_;
  assign new_n227_ = new_n224_ & new_n225_;
  assign new_n228_ = new_n226_ & new_n227_;
  assign new_n229_ = new_n120_ & new_n153_;
  assign new_n230_ = new_n122_ & new_n229_;
  assign new_n231_ = new_n127_ & new_n132_;
  assign new_n232_ = new_n129_ & new_n231_;
  assign new_n233_ = ~new_n228_ & ~new_n230_;
  assign new_n234_ = ~new_n232_ & new_n233_;
  assign new_n235_ = ~i_48_ & new_n225_;
  assign new_n236_ = ~i_31_ & new_n133_;
  assign new_n237_ = ~i_53_ & new_n235_;
  assign new_n238_ = new_n236_ & new_n237_;
  assign new_n239_ = i_51_ & new_n107_;
  assign new_n240_ = ~i_11_ & new_n133_;
  assign new_n241_ = new_n172_ & new_n239_;
  assign new_n242_ = new_n240_ & new_n241_;
  assign new_n243_ = new_n106_ & new_n127_;
  assign new_n244_ = new_n129_ & new_n243_;
  assign new_n245_ = ~new_n238_ & ~new_n242_;
  assign new_n246_ = ~new_n244_ & new_n245_;
  assign new_n247_ = new_n223_ & new_n234_;
  assign new_n248_ = new_n246_ & new_n247_;
  assign new_n249_ = new_n161_ & new_n208_;
  assign new_n250_ = new_n248_ & new_n249_;
  assign new_n251_ = ~i_9_ & new_n133_;
  assign new_n252_ = new_n114_ & new_n213_;
  assign new_n253_ = new_n251_ & new_n252_;
  assign new_n254_ = new_n174_ & new_n179_;
  assign new_n255_ = new_n113_ & new_n178_;
  assign new_n256_ = new_n115_ & new_n255_;
  assign new_n257_ = ~new_n253_ & ~new_n254_;
  assign new_n258_ = ~new_n256_ & new_n257_;
  assign new_n259_ = i_43_ & ~i_38_;
  assign new_n260_ = i_1_ & new_n259_;
  assign new_n261_ = new_n155_ & new_n178_;
  assign new_n262_ = new_n260_ & new_n261_;
  assign new_n263_ = ~i_46_ & ~i_47_;
  assign new_n264_ = i_41_ & new_n263_;
  assign new_n265_ = new_n178_ & new_n213_;
  assign new_n266_ = new_n264_ & new_n265_;
  assign new_n267_ = ~i_47_ & new_n167_;
  assign new_n268_ = i_46_ & ~i_43_;
  assign new_n269_ = ~i_38_ & new_n268_;
  assign new_n270_ = new_n239_ & new_n267_;
  assign new_n271_ = new_n269_ & new_n270_;
  assign new_n272_ = new_n168_ & new_n214_;
  assign new_n273_ = new_n115_ & new_n272_;
  assign new_n274_ = ~new_n266_ & ~new_n271_;
  assign new_n275_ = ~new_n273_ & new_n274_;
  assign new_n276_ = new_n258_ & ~new_n262_;
  assign new_n277_ = new_n275_ & new_n276_;
  assign new_n278_ = i_53_ & i_51_;
  assign new_n279_ = i_29_ & new_n133_;
  assign new_n280_ = new_n213_ & new_n278_;
  assign new_n281_ = new_n279_ & new_n280_;
  assign new_n282_ = new_n113_ & new_n209_;
  assign new_n283_ = new_n115_ & new_n282_;
  assign new_n284_ = i_48_ & new_n171_;
  assign new_n285_ = i_29_ & new_n263_;
  assign new_n286_ = new_n178_ & new_n284_;
  assign new_n287_ = new_n285_ & new_n286_;
  assign new_n288_ = ~new_n281_ & ~new_n283_;
  assign new_n289_ = ~new_n287_ & new_n288_;
  assign new_n290_ = new_n150_ & new_n198_;
  assign new_n291_ = ~i_38_ & new_n133_;
  assign new_n292_ = new_n173_ & new_n224_;
  assign new_n293_ = new_n291_ & new_n292_;
  assign new_n294_ = ~i_48_ & new_n152_;
  assign new_n295_ = ~i_39_ & new_n133_;
  assign new_n296_ = new_n120_ & new_n294_;
  assign new_n297_ = new_n295_ & new_n296_;
  assign new_n298_ = ~new_n290_ & ~new_n293_;
  assign new_n299_ = ~new_n297_ & new_n298_;
  assign new_n300_ = new_n180_ & new_n226_;
  assign new_n301_ = i_49_ & new_n118_;
  assign new_n302_ = ~i_46_ & new_n121_;
  assign new_n303_ = new_n127_ & new_n301_;
  assign new_n304_ = new_n302_ & new_n303_;
  assign new_n305_ = i_49_ & new_n152_;
  assign new_n306_ = new_n127_ & new_n305_;
  assign new_n307_ = new_n155_ & new_n306_;
  assign new_n308_ = ~new_n300_ & ~new_n304_;
  assign new_n309_ = ~new_n307_ & new_n308_;
  assign new_n310_ = new_n289_ & new_n299_;
  assign new_n311_ = new_n309_ & new_n310_;
  assign new_n312_ = new_n277_ & new_n311_;
  assign new_n313_ = i_50_ & ~i_52_;
  assign new_n314_ = ~i_49_ & new_n313_;
  assign new_n315_ = i_53_ & new_n314_;
  assign new_n316_ = new_n129_ & new_n315_;
  assign new_n317_ = i_50_ & ~i_51_;
  assign new_n318_ = ~i_49_ & new_n317_;
  assign new_n319_ = new_n162_ & new_n318_;
  assign new_n320_ = new_n129_ & new_n319_;
  assign new_n321_ = i_49_ & new_n317_;
  assign new_n322_ = new_n127_ & new_n321_;
  assign new_n323_ = new_n155_ & new_n322_;
  assign new_n324_ = ~new_n316_ & ~new_n320_;
  assign new_n325_ = ~new_n323_ & new_n324_;
  assign new_n326_ = ~i_52_ & ~i_51_;
  assign new_n327_ = i_49_ & new_n326_;
  assign new_n328_ = i_53_ & new_n327_;
  assign new_n329_ = new_n155_ & new_n328_;
  assign new_n330_ = ~i_50_ & new_n326_;
  assign new_n331_ = i_49_ & i_47_;
  assign new_n332_ = ~i_46_ & new_n331_;
  assign new_n333_ = i_53_ & new_n330_;
  assign new_n334_ = new_n332_ & new_n333_;
  assign new_n335_ = new_n162_ & new_n305_;
  assign new_n336_ = new_n129_ & new_n335_;
  assign new_n337_ = ~new_n329_ & ~new_n334_;
  assign new_n338_ = ~new_n336_ & new_n337_;
  assign new_n339_ = new_n106_ & new_n162_;
  assign new_n340_ = new_n302_ & new_n339_;
  assign new_n341_ = new_n107_ & new_n119_;
  assign new_n342_ = new_n129_ & new_n341_;
  assign new_n343_ = i_49_ & new_n184_;
  assign new_n344_ = i_53_ & new_n343_;
  assign new_n345_ = new_n155_ & new_n344_;
  assign new_n346_ = ~new_n340_ & ~new_n342_;
  assign new_n347_ = ~new_n345_ & new_n346_;
  assign new_n348_ = new_n325_ & new_n338_;
  assign new_n349_ = new_n347_ & new_n348_;
  assign new_n350_ = new_n122_ & new_n341_;
  assign new_n351_ = new_n155_ & new_n335_;
  assign new_n352_ = new_n107_ & new_n305_;
  assign new_n353_ = new_n155_ & new_n352_;
  assign new_n354_ = ~new_n350_ & ~new_n351_;
  assign new_n355_ = ~new_n353_ & new_n354_;
  assign new_n356_ = new_n106_ & new_n120_;
  assign new_n357_ = new_n122_ & new_n356_;
  assign new_n358_ = new_n127_ & new_n318_;
  assign new_n359_ = new_n129_ & new_n358_;
  assign new_n360_ = new_n122_ & new_n156_;
  assign new_n361_ = ~new_n357_ & ~new_n359_;
  assign new_n362_ = ~new_n360_ & new_n361_;
  assign new_n363_ = new_n120_ & new_n132_;
  assign new_n364_ = new_n129_ & new_n363_;
  assign new_n365_ = new_n120_ & new_n318_;
  assign new_n366_ = new_n155_ & new_n365_;
  assign new_n367_ = i_39_ & new_n263_;
  assign new_n368_ = new_n163_ & new_n284_;
  assign new_n369_ = new_n367_ & new_n368_;
  assign new_n370_ = ~new_n364_ & ~new_n366_;
  assign new_n371_ = ~new_n369_ & new_n370_;
  assign new_n372_ = new_n355_ & new_n362_;
  assign new_n373_ = new_n371_ & new_n372_;
  assign new_n374_ = new_n132_ & new_n162_;
  assign new_n375_ = new_n155_ & new_n374_;
  assign new_n376_ = ~i_47_ & ~i_48_;
  assign new_n377_ = i_46_ & new_n376_;
  assign new_n378_ = new_n110_ & new_n377_;
  assign new_n379_ = ~i_49_ & i_51_;
  assign new_n380_ = new_n155_ & new_n379_;
  assign new_n381_ = ~new_n375_ & ~new_n378_;
  assign new_n382_ = ~new_n380_ & new_n381_;
  assign new_n383_ = i_50_ & new_n326_;
  assign new_n384_ = ~i_53_ & new_n383_;
  assign new_n385_ = new_n155_ & new_n384_;
  assign new_n386_ = ~i_49_ & new_n225_;
  assign new_n387_ = ~i_53_ & new_n386_;
  assign new_n388_ = new_n155_ & new_n387_;
  assign new_n389_ = new_n162_ & new_n321_;
  assign new_n390_ = new_n129_ & new_n389_;
  assign new_n391_ = ~new_n385_ & ~new_n388_;
  assign new_n392_ = ~new_n390_ & new_n391_;
  assign new_n393_ = new_n302_ & new_n356_;
  assign new_n394_ = new_n107_ & new_n301_;
  assign o_33_ = new_n155_ & new_n394_;
  assign new_n396_ = new_n162_ & new_n301_;
  assign new_n397_ = new_n129_ & new_n396_;
  assign new_n398_ = ~new_n393_ & ~o_33_;
  assign new_n399_ = ~new_n397_ & new_n398_;
  assign new_n400_ = new_n382_ & new_n392_;
  assign new_n401_ = new_n399_ & new_n400_;
  assign new_n402_ = new_n349_ & new_n373_;
  assign new_n403_ = new_n401_ & new_n402_;
  assign new_n404_ = new_n250_ & new_n312_;
  assign o_1_ = ~new_n403_ | ~new_n404_;
  assign new_n406_ = ~i_46_ & new_n376_;
  assign new_n407_ = new_n319_ & new_n406_;
  assign new_n408_ = ~i_25_ & ~i_11_;
  assign new_n409_ = ~i_10_ & new_n408_;
  assign new_n410_ = new_n321_ & new_n377_;
  assign new_n411_ = new_n409_ & new_n410_;
  assign new_n412_ = new_n162_ & new_n411_;
  assign new_n413_ = i_10_ & new_n108_;
  assign new_n414_ = new_n172_ & new_n209_;
  assign new_n415_ = new_n413_ & new_n414_;
  assign new_n416_ = ~new_n407_ & ~new_n412_;
  assign new_n417_ = ~new_n415_ & new_n416_;
  assign new_n418_ = new_n155_ & new_n243_;
  assign new_n419_ = new_n123_ & new_n406_;
  assign new_n420_ = new_n339_ & new_n406_;
  assign new_n421_ = ~new_n418_ & ~new_n419_;
  assign new_n422_ = ~new_n420_ & new_n421_;
  assign new_n423_ = i_25_ & new_n108_;
  assign new_n424_ = new_n414_ & new_n423_;
  assign new_n425_ = i_11_ & new_n108_;
  assign new_n426_ = new_n414_ & new_n425_;
  assign new_n427_ = new_n120_ & new_n305_;
  assign new_n428_ = new_n406_ & new_n427_;
  assign new_n429_ = ~new_n424_ & ~new_n426_;
  assign new_n430_ = ~new_n428_ & new_n429_;
  assign new_n431_ = new_n107_ & new_n132_;
  assign new_n432_ = new_n377_ & new_n431_;
  assign new_n433_ = ~new_n342_ & ~new_n366_;
  assign new_n434_ = ~new_n432_ & new_n433_;
  assign new_n435_ = new_n422_ & new_n430_;
  assign new_n436_ = new_n434_ & new_n435_;
  assign o_19_ = ~new_n417_ | ~new_n436_;
  assign new_n438_ = ~i_49_ & i_48_;
  assign new_n439_ = ~i_47_ & new_n438_;
  assign new_n440_ = ~i_50_ & new_n184_;
  assign new_n441_ = i_46_ & i_38_;
  assign new_n442_ = ~i_37_ & new_n441_;
  assign new_n443_ = new_n439_ & new_n440_;
  assign new_n444_ = new_n442_ & new_n443_;
  assign new_n445_ = ~i_53_ & new_n444_;
  assign new_n446_ = i_46_ & i_43_;
  assign new_n447_ = ~i_37_ & new_n446_;
  assign new_n448_ = new_n443_ & new_n447_;
  assign new_n449_ = ~i_53_ & new_n448_;
  assign new_n450_ = ~new_n262_ & ~new_n449_;
  assign new_n451_ = ~new_n254_ & new_n450_;
  assign new_n452_ = ~new_n445_ & new_n451_;
  assign new_n453_ = new_n129_ & new_n374_;
  assign new_n454_ = new_n107_ & new_n321_;
  assign o_14_ = new_n302_ & new_n454_;
  assign new_n456_ = ~new_n453_ & ~o_14_;
  assign new_n457_ = ~new_n217_ & new_n456_;
  assign new_n458_ = new_n120_ & new_n321_;
  assign new_n459_ = new_n129_ & new_n458_;
  assign new_n460_ = i_30_ & new_n263_;
  assign new_n461_ = new_n163_ & new_n172_;
  assign new_n462_ = new_n460_ & new_n461_;
  assign new_n463_ = ~new_n459_ & ~new_n462_;
  assign new_n464_ = ~new_n157_ & new_n463_;
  assign new_n465_ = new_n335_ & new_n377_;
  assign new_n466_ = ~new_n212_ & ~new_n465_;
  assign new_n467_ = ~new_n221_ & new_n466_;
  assign new_n468_ = new_n457_ & new_n464_;
  assign new_n469_ = new_n467_ & new_n468_;
  assign new_n470_ = i_35_ & new_n263_;
  assign new_n471_ = new_n241_ & new_n470_;
  assign new_n472_ = ~i_20_ & new_n133_;
  assign new_n473_ = new_n224_ & new_n239_;
  assign new_n474_ = new_n472_ & new_n473_;
  assign new_n475_ = ~i_29_ & new_n263_;
  assign new_n476_ = new_n225_ & new_n284_;
  assign new_n477_ = new_n475_ & new_n476_;
  assign new_n478_ = ~new_n471_ & ~new_n474_;
  assign new_n479_ = ~new_n477_ & new_n478_;
  assign new_n480_ = ~i_3_ & new_n263_;
  assign new_n481_ = new_n272_ & new_n480_;
  assign new_n482_ = ~i_20_ & new_n263_;
  assign new_n483_ = new_n145_ & new_n225_;
  assign new_n484_ = new_n482_ & new_n483_;
  assign o_27_ = new_n229_ & new_n302_;
  assign new_n486_ = ~new_n481_ & ~new_n484_;
  assign new_n487_ = ~o_27_ & new_n486_;
  assign new_n488_ = new_n156_ & new_n302_;
  assign new_n489_ = new_n158_ & ~new_n488_;
  assign new_n490_ = new_n479_ & new_n487_;
  assign new_n491_ = new_n489_ & new_n490_;
  assign new_n492_ = new_n162_ & new_n284_;
  assign new_n493_ = new_n285_ & new_n492_;
  assign new_n494_ = ~i_7_ & new_n263_;
  assign new_n495_ = new_n239_ & new_n284_;
  assign new_n496_ = new_n494_ & new_n495_;
  assign new_n497_ = ~new_n351_ & ~new_n493_;
  assign new_n498_ = ~new_n496_ & new_n497_;
  assign o_36_ = new_n302_ & new_n306_;
  assign new_n500_ = i_19_ & new_n263_;
  assign new_n501_ = new_n145_ & new_n196_;
  assign new_n502_ = new_n500_ & new_n501_;
  assign new_n503_ = ~i_52_ & new_n321_;
  assign new_n504_ = new_n155_ & new_n503_;
  assign new_n505_ = ~o_36_ & ~new_n502_;
  assign new_n506_ = ~new_n504_ & new_n505_;
  assign new_n507_ = new_n155_ & new_n231_;
  assign o_37_ = new_n302_ & new_n352_;
  assign new_n509_ = ~new_n350_ & ~new_n507_;
  assign new_n510_ = ~o_37_ & new_n509_;
  assign new_n511_ = new_n498_ & new_n506_;
  assign new_n512_ = new_n510_ & new_n511_;
  assign new_n513_ = new_n469_ & new_n491_;
  assign new_n514_ = new_n512_ & new_n513_;
  assign new_n515_ = ~new_n300_ & ~new_n307_;
  assign new_n516_ = ~new_n188_ & new_n515_;
  assign new_n517_ = i_7_ & new_n263_;
  assign new_n518_ = new_n495_ & new_n517_;
  assign new_n519_ = ~i_17_ & new_n263_;
  assign new_n520_ = new_n145_ & new_n214_;
  assign new_n521_ = new_n519_ & new_n520_;
  assign new_n522_ = ~new_n283_ & ~new_n518_;
  assign new_n523_ = ~new_n521_ & new_n522_;
  assign new_n524_ = ~new_n181_ & ~new_n189_;
  assign new_n525_ = ~new_n170_ & new_n524_;
  assign new_n526_ = new_n516_ & new_n523_;
  assign new_n527_ = new_n525_ & new_n526_;
  assign new_n528_ = i_37_ & new_n263_;
  assign new_n529_ = new_n169_ & new_n528_;
  assign new_n530_ = i_48_ & new_n379_;
  assign new_n531_ = i_20_ & new_n263_;
  assign new_n532_ = new_n127_ & new_n530_;
  assign new_n533_ = new_n531_ & new_n532_;
  assign new_n534_ = ~new_n529_ & ~new_n533_;
  assign new_n535_ = ~new_n290_ & new_n534_;
  assign new_n536_ = i_3_ & new_n376_;
  assign new_n537_ = new_n303_ & new_n536_;
  assign new_n538_ = i_3_ & new_n263_;
  assign new_n539_ = new_n272_ & new_n538_;
  assign new_n540_ = ~new_n256_ & ~new_n537_;
  assign new_n541_ = ~new_n539_ & new_n540_;
  assign new_n542_ = ~i_16_ & new_n108_;
  assign new_n543_ = new_n211_ & new_n542_;
  assign new_n544_ = i_28_ & new_n133_;
  assign new_n545_ = new_n114_ & new_n137_;
  assign new_n546_ = new_n544_ & new_n545_;
  assign new_n547_ = ~i_4_ & new_n108_;
  assign new_n548_ = new_n282_ & new_n547_;
  assign new_n549_ = ~new_n543_ & ~new_n546_;
  assign new_n550_ = ~new_n548_ & new_n549_;
  assign new_n551_ = new_n535_ & new_n541_;
  assign new_n552_ = new_n550_ & new_n551_;
  assign new_n553_ = ~i_3_ & new_n108_;
  assign new_n554_ = new_n165_ & new_n553_;
  assign new_n555_ = new_n145_ & new_n209_;
  assign new_n556_ = new_n531_ & new_n555_;
  assign new_n557_ = new_n174_ & new_n531_;
  assign new_n558_ = ~new_n554_ & ~new_n556_;
  assign new_n559_ = ~new_n557_ & new_n558_;
  assign new_n560_ = new_n113_ & new_n326_;
  assign new_n561_ = new_n547_ & new_n560_;
  assign new_n562_ = i_44_ & new_n263_;
  assign new_n563_ = new_n198_ & new_n562_;
  assign new_n564_ = new_n272_ & new_n547_;
  assign new_n565_ = ~new_n561_ & ~new_n563_;
  assign new_n566_ = ~new_n564_ & new_n565_;
  assign new_n567_ = i_8_ & new_n263_;
  assign new_n568_ = new_n414_ & new_n567_;
  assign new_n569_ = ~i_46_ & i_48_;
  assign new_n570_ = ~i_29_ & new_n569_;
  assign new_n571_ = new_n328_ & new_n570_;
  assign new_n572_ = i_29_ & new_n569_;
  assign new_n573_ = new_n365_ & new_n572_;
  assign new_n574_ = ~new_n568_ & ~new_n571_;
  assign new_n575_ = ~new_n573_ & new_n574_;
  assign new_n576_ = new_n559_ & new_n566_;
  assign new_n577_ = new_n575_ & new_n576_;
  assign new_n578_ = new_n527_ & new_n552_;
  assign new_n579_ = new_n577_ & new_n578_;
  assign new_n580_ = new_n129_ & new_n339_;
  assign new_n581_ = ~i_46_ & new_n182_;
  assign new_n582_ = new_n333_ & new_n581_;
  assign new_n583_ = new_n122_ & new_n130_;
  assign new_n584_ = ~new_n580_ & ~new_n582_;
  assign new_n585_ = ~new_n583_ & new_n584_;
  assign new_n586_ = new_n377_ & new_n458_;
  assign new_n587_ = ~i_41_ & new_n569_;
  assign new_n588_ = new_n120_ & new_n301_;
  assign new_n589_ = new_n587_ & new_n588_;
  assign new_n590_ = i_42_ & new_n263_;
  assign new_n591_ = new_n214_ & new_n284_;
  assign new_n592_ = new_n590_ & new_n591_;
  assign new_n593_ = ~new_n586_ & ~new_n589_;
  assign new_n594_ = ~new_n592_ & new_n593_;
  assign new_n595_ = ~i_39_ & new_n263_;
  assign new_n596_ = new_n368_ & new_n595_;
  assign new_n597_ = new_n302_ & new_n322_;
  assign new_n598_ = ~new_n323_ & ~new_n596_;
  assign new_n599_ = ~new_n597_ & new_n598_;
  assign new_n600_ = new_n585_ & new_n594_;
  assign new_n601_ = new_n599_ & new_n600_;
  assign new_n602_ = i_8_ & new_n569_;
  assign new_n603_ = new_n384_ & new_n602_;
  assign o_38_ = new_n302_ & new_n431_;
  assign new_n605_ = ~new_n603_ & ~o_38_;
  assign new_n606_ = ~new_n366_ & new_n605_;
  assign new_n607_ = new_n153_ & new_n162_;
  assign new_n608_ = new_n302_ & new_n607_;
  assign new_n609_ = new_n229_ & new_n406_;
  assign new_n610_ = ~new_n353_ & ~new_n608_;
  assign new_n611_ = ~new_n609_ & new_n610_;
  assign new_n612_ = new_n155_ & new_n358_;
  assign new_n613_ = new_n129_ & new_n303_;
  assign new_n614_ = ~new_n369_ & ~new_n612_;
  assign new_n615_ = ~new_n613_ & new_n614_;
  assign new_n616_ = new_n606_ & new_n611_;
  assign new_n617_ = new_n615_ & new_n616_;
  assign new_n618_ = ~new_n378_ & ~new_n385_;
  assign new_n619_ = ~new_n375_ & new_n618_;
  assign new_n620_ = new_n129_ & new_n352_;
  assign new_n621_ = ~new_n345_ & ~new_n620_;
  assign new_n622_ = ~new_n388_ & new_n621_;
  assign new_n623_ = i_52_ & i_51_;
  assign new_n624_ = i_50_ & new_n623_;
  assign new_n625_ = ~i_46_ & new_n438_;
  assign new_n626_ = ~i_53_ & new_n624_;
  assign new_n627_ = new_n625_ & new_n626_;
  assign new_n628_ = ~new_n380_ & ~o_33_;
  assign new_n629_ = ~new_n627_ & new_n628_;
  assign new_n630_ = new_n619_ & new_n622_;
  assign new_n631_ = new_n629_ & new_n630_;
  assign new_n632_ = new_n601_ & new_n617_;
  assign new_n633_ = new_n631_ & new_n632_;
  assign new_n634_ = new_n514_ & new_n579_;
  assign new_n635_ = new_n633_ & new_n634_;
  assign o_2_ = ~new_n452_ | ~new_n635_;
  assign new_n637_ = i_24_ & new_n108_;
  assign new_n638_ = new_n184_ & new_n224_;
  assign new_n639_ = new_n637_ & new_n638_;
  assign new_n640_ = new_n231_ & new_n377_;
  assign new_n641_ = ~new_n639_ & ~new_n640_;
  assign new_n642_ = ~new_n459_ & new_n641_;
  assign new_n643_ = i_21_ & new_n108_;
  assign new_n644_ = new_n137_ & new_n163_;
  assign new_n645_ = new_n643_ & new_n644_;
  assign new_n646_ = new_n322_ & new_n377_;
  assign new_n647_ = ~new_n474_ & ~new_n645_;
  assign new_n648_ = ~new_n646_ & new_n647_;
  assign new_n649_ = new_n339_ & new_n377_;
  assign new_n650_ = ~i_21_ & new_n108_;
  assign new_n651_ = ~i_53_ & new_n137_;
  assign new_n652_ = new_n650_ & new_n651_;
  assign new_n653_ = ~new_n453_ & ~new_n649_;
  assign new_n654_ = ~new_n652_ & new_n653_;
  assign new_n655_ = new_n642_ & new_n648_;
  assign new_n656_ = new_n654_ & new_n655_;
  assign new_n657_ = new_n130_ & new_n377_;
  assign new_n658_ = ~new_n564_ & ~new_n657_;
  assign new_n659_ = ~new_n554_ & new_n658_;
  assign new_n660_ = i_41_ & new_n108_;
  assign new_n661_ = new_n137_ & new_n178_;
  assign new_n662_ = new_n660_ & new_n661_;
  assign new_n663_ = ~new_n424_ & ~new_n662_;
  assign new_n664_ = ~new_n561_ & new_n663_;
  assign new_n665_ = i_40_ & new_n263_;
  assign new_n666_ = new_n168_ & new_n239_;
  assign new_n667_ = new_n665_ & new_n666_;
  assign new_n668_ = new_n377_ & new_n427_;
  assign new_n669_ = new_n306_ & new_n377_;
  assign new_n670_ = ~new_n667_ & ~new_n668_;
  assign new_n671_ = ~new_n669_ & new_n670_;
  assign new_n672_ = new_n659_ & new_n664_;
  assign new_n673_ = new_n671_ & new_n672_;
  assign new_n674_ = ~i_46_ & ~i_48_;
  assign new_n675_ = i_13_ & new_n674_;
  assign new_n676_ = new_n156_ & new_n675_;
  assign new_n677_ = new_n110_ & new_n129_;
  assign new_n678_ = new_n352_ & new_n377_;
  assign new_n679_ = ~new_n676_ & ~new_n677_;
  assign new_n680_ = ~new_n678_ & new_n679_;
  assign new_n681_ = ~i_50_ & new_n225_;
  assign new_n682_ = ~i_49_ & ~i_48_;
  assign new_n683_ = ~i_47_ & new_n682_;
  assign new_n684_ = i_53_ & new_n681_;
  assign new_n685_ = new_n683_ & new_n684_;
  assign new_n686_ = ~i_34_ & new_n263_;
  assign new_n687_ = new_n145_ & new_n163_;
  assign new_n688_ = new_n686_ & new_n687_;
  assign new_n689_ = ~new_n465_ & ~new_n685_;
  assign new_n690_ = ~new_n688_ & new_n689_;
  assign new_n691_ = new_n122_ & new_n358_;
  assign new_n692_ = new_n129_ & new_n454_;
  assign new_n693_ = ~new_n691_ & ~new_n692_;
  assign new_n694_ = ~new_n507_ & new_n693_;
  assign new_n695_ = new_n680_ & new_n690_;
  assign new_n696_ = new_n694_ & new_n695_;
  assign new_n697_ = new_n656_ & new_n673_;
  assign new_n698_ = new_n696_ & new_n697_;
  assign new_n699_ = i_6_ & new_n108_;
  assign new_n700_ = new_n198_ & new_n699_;
  assign new_n701_ = i_9_ & new_n133_;
  assign new_n702_ = new_n107_ & new_n294_;
  assign new_n703_ = new_n701_ & new_n702_;
  assign new_n704_ = i_20_ & new_n108_;
  assign new_n705_ = new_n169_ & new_n704_;
  assign new_n706_ = ~new_n700_ & ~new_n703_;
  assign new_n707_ = ~new_n705_ & new_n706_;
  assign new_n708_ = i_39_ & new_n133_;
  assign new_n709_ = new_n265_ & new_n708_;
  assign new_n710_ = ~new_n445_ & ~new_n449_;
  assign new_n711_ = ~new_n709_ & new_n710_;
  assign new_n712_ = new_n303_ & new_n377_;
  assign new_n713_ = ~i_41_ & new_n108_;
  assign new_n714_ = new_n661_ & new_n713_;
  assign new_n715_ = ~i_39_ & new_n108_;
  assign new_n716_ = new_n213_ & new_n623_;
  assign new_n717_ = new_n715_ & new_n716_;
  assign new_n718_ = ~new_n712_ & ~new_n714_;
  assign new_n719_ = ~new_n717_ & new_n718_;
  assign new_n720_ = new_n707_ & new_n711_;
  assign new_n721_ = new_n719_ & new_n720_;
  assign new_n722_ = ~i_28_ & ~i_25_;
  assign new_n723_ = ~i_22_ & new_n722_;
  assign new_n724_ = new_n119_ & new_n377_;
  assign new_n725_ = new_n723_ & new_n724_;
  assign new_n726_ = new_n120_ & new_n725_;
  assign new_n727_ = ~new_n412_ & ~new_n726_;
  assign new_n728_ = ~i_24_ & new_n108_;
  assign new_n729_ = new_n196_ & new_n224_;
  assign new_n730_ = new_n728_ & new_n729_;
  assign new_n731_ = ~new_n518_ & ~new_n548_;
  assign new_n732_ = ~new_n730_ & new_n731_;
  assign new_n733_ = i_31_ & new_n133_;
  assign new_n734_ = new_n209_ & new_n213_;
  assign new_n735_ = new_n733_ & new_n734_;
  assign new_n736_ = new_n549_ & ~new_n735_;
  assign new_n737_ = new_n196_ & new_n284_;
  assign new_n738_ = new_n264_ & new_n737_;
  assign new_n739_ = ~new_n415_ & ~new_n738_;
  assign new_n740_ = ~new_n426_ & new_n739_;
  assign new_n741_ = new_n732_ & new_n736_;
  assign new_n742_ = new_n740_ & new_n741_;
  assign new_n743_ = new_n721_ & new_n727_;
  assign new_n744_ = new_n742_ & new_n743_;
  assign new_n745_ = i_11_ & new_n133_;
  assign new_n746_ = new_n107_ & new_n172_;
  assign new_n747_ = new_n745_ & new_n746_;
  assign new_n748_ = ~i_49_ & new_n138_;
  assign new_n749_ = new_n377_ & new_n748_;
  assign new_n750_ = i_17_ & new_n263_;
  assign new_n751_ = new_n231_ & new_n750_;
  assign new_n752_ = ~new_n747_ & ~new_n749_;
  assign new_n753_ = ~new_n751_ & new_n752_;
  assign new_n754_ = ~new_n580_ & ~new_n586_;
  assign new_n755_ = ~new_n583_ & new_n754_;
  assign new_n756_ = new_n377_ & new_n396_;
  assign new_n757_ = new_n119_ & new_n162_;
  assign new_n758_ = new_n129_ & new_n757_;
  assign new_n759_ = new_n374_ & new_n377_;
  assign new_n760_ = ~new_n756_ & ~new_n758_;
  assign new_n761_ = ~new_n759_ & new_n760_;
  assign new_n762_ = new_n753_ & new_n755_;
  assign new_n763_ = new_n761_ & new_n762_;
  assign new_n764_ = i_22_ & new_n108_;
  assign new_n765_ = new_n137_ & new_n184_;
  assign new_n766_ = new_n764_ & new_n765_;
  assign new_n767_ = new_n377_ & new_n454_;
  assign new_n768_ = i_28_ & new_n108_;
  assign new_n769_ = new_n765_ & new_n768_;
  assign new_n770_ = ~new_n766_ & ~new_n767_;
  assign new_n771_ = ~new_n769_ & new_n770_;
  assign new_n772_ = new_n122_ & new_n339_;
  assign new_n773_ = new_n356_ & new_n377_;
  assign new_n774_ = ~new_n772_ & ~new_n773_;
  assign new_n775_ = ~new_n612_ & new_n774_;
  assign new_n776_ = new_n423_ & new_n765_;
  assign new_n777_ = new_n155_ & new_n389_;
  assign new_n778_ = ~new_n613_ & ~new_n776_;
  assign new_n779_ = ~new_n777_ & new_n778_;
  assign new_n780_ = new_n771_ & new_n775_;
  assign new_n781_ = new_n779_ & new_n780_;
  assign o_46_ = new_n155_ & new_n303_;
  assign new_n783_ = new_n155_ & new_n396_;
  assign new_n784_ = ~new_n432_ & ~o_46_;
  assign new_n785_ = ~new_n783_ & new_n784_;
  assign new_n786_ = new_n229_ & new_n377_;
  assign new_n787_ = new_n358_ & new_n377_;
  assign new_n788_ = ~new_n620_ & ~new_n786_;
  assign new_n789_ = ~new_n787_ & new_n788_;
  assign o_42_ = new_n231_ & new_n406_;
  assign new_n791_ = i_50_ & new_n184_;
  assign new_n792_ = ~i_53_ & new_n791_;
  assign new_n793_ = new_n377_ & new_n792_;
  assign o_43_ = new_n363_ & new_n406_;
  assign new_n795_ = ~o_42_ & ~new_n793_;
  assign new_n796_ = ~o_43_ & new_n795_;
  assign new_n797_ = new_n785_ & new_n789_;
  assign new_n798_ = new_n796_ & new_n797_;
  assign new_n799_ = new_n763_ & new_n781_;
  assign new_n800_ = new_n798_ & new_n799_;
  assign new_n801_ = new_n698_ & new_n744_;
  assign o_0_ = ~new_n800_ | ~new_n801_;
  assign o_29_ = new_n155_ & new_n588_;
  assign new_n804_ = ~i_24_ & new_n263_;
  assign new_n805_ = new_n255_ & new_n804_;
  assign o_39_ = new_n393_ | new_n805_;
  assign new_n807_ = ~i_19_ & new_n263_;
  assign new_n808_ = new_n501_ & new_n807_;
  assign new_n809_ = new_n505_ & ~o_38_;
  assign o_25_ = new_n808_ | ~new_n809_;
  assign new_n811_ = ~new_n507_ & ~new_n692_;
  assign new_n812_ = ~new_n329_ & new_n811_;
  assign new_n813_ = i_53_ & new_n791_;
  assign new_n814_ = new_n129_ & new_n813_;
  assign new_n815_ = ~new_n157_ & ~new_n453_;
  assign new_n816_ = ~new_n814_ & new_n815_;
  assign new_n817_ = ~new_n336_ & ~new_n613_;
  assign new_n818_ = ~new_n620_ & new_n817_;
  assign new_n819_ = new_n812_ & new_n816_;
  assign o_12_ = ~new_n818_ | ~new_n819_;
  assign new_n821_ = ~new_n359_ & ~new_n465_;
  assign o_26_ = new_n612_ | ~new_n821_;
  assign new_n823_ = new_n341_ & new_n377_;
  assign new_n824_ = new_n110_ & new_n406_;
  assign new_n825_ = new_n358_ & new_n406_;
  assign new_n826_ = ~new_n824_ & ~new_n825_;
  assign new_n827_ = ~new_n580_ & new_n826_;
  assign new_n828_ = ~i_16_ & new_n263_;
  assign new_n829_ = new_n644_ & new_n828_;
  assign new_n830_ = i_16_ & new_n263_;
  assign new_n831_ = new_n644_ & new_n830_;
  assign new_n832_ = ~new_n640_ & ~new_n829_;
  assign new_n833_ = ~new_n831_ & new_n832_;
  assign new_n834_ = ~new_n340_ & ~new_n390_;
  assign new_n835_ = ~new_n393_ & new_n834_;
  assign new_n836_ = new_n827_ & new_n833_;
  assign new_n837_ = new_n835_ & new_n836_;
  assign o_11_ = new_n823_ | ~new_n837_;
  assign new_n839_ = new_n302_ & new_n319_;
  assign new_n840_ = new_n302_ & new_n341_;
  assign new_n841_ = ~new_n839_ & ~new_n840_;
  assign new_n842_ = ~new_n459_ & new_n841_;
  assign new_n843_ = ~new_n597_ & ~new_n608_;
  assign new_n844_ = ~new_n759_ & new_n843_;
  assign o_35_ = ~new_n842_ | ~new_n844_;
  assign new_n846_ = ~new_n364_ & ~new_n507_;
  assign new_n847_ = ~new_n613_ & new_n846_;
  assign new_n848_ = ~new_n131_ & ~new_n453_;
  assign new_n849_ = ~new_n375_ & ~new_n620_;
  assign new_n850_ = ~new_n397_ & new_n849_;
  assign new_n851_ = new_n847_ & new_n848_;
  assign o_28_ = ~new_n850_ | ~new_n851_;
  assign o_13_ = new_n156_ & new_n406_;
  assign new_n854_ = ~new_n334_ & ~new_n353_;
  assign o_34_ = new_n336_ | ~new_n854_;
  assign o_21_ = new_n773_ | new_n783_;
  assign new_n857_ = ~new_n242_ & ~new_n692_;
  assign new_n858_ = ~new_n777_ & new_n857_;
  assign new_n859_ = ~new_n199_ & ~o_13_;
  assign new_n860_ = ~new_n649_ & new_n859_;
  assign new_n861_ = ~new_n747_ & ~new_n758_;
  assign new_n862_ = ~new_n787_ & new_n861_;
  assign new_n863_ = new_n858_ & new_n860_;
  assign new_n864_ = new_n862_ & new_n863_;
  assign o_16_ = new_n290_ | ~new_n864_;
  assign new_n866_ = ~new_n242_ & ~new_n814_;
  assign new_n867_ = ~new_n692_ & new_n866_;
  assign new_n868_ = ~new_n504_ & ~new_n747_;
  assign new_n869_ = ~new_n342_ & new_n868_;
  assign new_n870_ = ~new_n230_ & new_n867_;
  assign o_40_ = ~new_n869_ | ~new_n870_;
  assign new_n872_ = i_25_ & new_n263_;
  assign new_n873_ = new_n137_ & new_n239_;
  assign new_n874_ = new_n872_ & new_n873_;
  assign new_n875_ = ~new_n175_ & ~new_n307_;
  assign new_n876_ = ~new_n874_ & new_n875_;
  assign new_n877_ = new_n114_ & new_n224_;
  assign new_n878_ = new_n872_ & new_n877_;
  assign new_n879_ = ~i_25_ & new_n263_;
  assign new_n880_ = new_n877_ & new_n879_;
  assign new_n881_ = ~new_n808_ & ~new_n878_;
  assign new_n882_ = ~new_n880_ & new_n881_;
  assign new_n883_ = new_n873_ & new_n879_;
  assign new_n884_ = ~new_n502_ & ~new_n883_;
  assign new_n885_ = ~new_n767_ & new_n884_;
  assign new_n886_ = new_n876_ & new_n882_;
  assign new_n887_ = new_n885_ & new_n886_;
  assign o_22_ = new_n254_ | ~new_n887_;
  assign new_n889_ = ~i_37_ & new_n263_;
  assign new_n890_ = new_n169_ & new_n889_;
  assign new_n891_ = i_50_ & new_n225_;
  assign new_n892_ = ~i_49_ & ~i_47_;
  assign new_n893_ = i_46_ & new_n892_;
  assign new_n894_ = ~i_53_ & new_n891_;
  assign new_n895_ = new_n893_ & new_n894_;
  assign new_n896_ = ~new_n529_ & ~new_n890_;
  assign new_n897_ = ~new_n895_ & new_n896_;
  assign new_n898_ = ~new_n273_ & ~new_n537_;
  assign new_n899_ = ~new_n539_ & new_n898_;
  assign new_n900_ = ~i_52_ & new_n106_;
  assign new_n901_ = new_n155_ & new_n900_;
  assign new_n902_ = ~new_n166_ & ~new_n561_;
  assign new_n903_ = ~new_n901_ & new_n902_;
  assign new_n904_ = new_n897_ & new_n899_;
  assign new_n905_ = new_n903_ & new_n904_;
  assign new_n906_ = ~new_n117_ & ~new_n230_;
  assign new_n907_ = ~new_n351_ & new_n906_;
  assign new_n908_ = ~new_n554_ & ~new_n564_;
  assign new_n909_ = ~new_n481_ & new_n908_;
  assign new_n910_ = ~i_3_ & new_n376_;
  assign new_n911_ = new_n303_ & new_n910_;
  assign new_n912_ = ~new_n336_ & ~new_n911_;
  assign new_n913_ = ~new_n627_ & new_n912_;
  assign new_n914_ = new_n907_ & new_n909_;
  assign new_n915_ = new_n913_ & new_n914_;
  assign new_n916_ = ~new_n256_ & new_n905_;
  assign o_15_ = ~new_n915_ | ~new_n916_;
  assign o_32_ = o_37_ | new_n712_;
  assign new_n919_ = ~i_49_ & i_47_;
  assign new_n920_ = ~i_46_ & new_n919_;
  assign o_23_ = new_n626_ & new_n920_;
  assign new_n922_ = ~new_n657_ & ~new_n668_;
  assign new_n923_ = ~new_n350_ & new_n922_;
  assign new_n924_ = i_23_ & new_n133_;
  assign new_n925_ = new_n116_ & new_n924_;
  assign new_n926_ = ~new_n320_ & ~new_n772_;
  assign new_n927_ = ~new_n342_ & new_n926_;
  assign new_n928_ = new_n923_ & ~new_n925_;
  assign o_18_ = ~new_n927_ | ~new_n928_;
  assign o_31_ = new_n374_ & new_n406_;
  assign o_24_ = new_n390_ | new_n759_;
  assign new_n932_ = new_n216_ & new_n830_;
  assign new_n933_ = new_n216_ & new_n828_;
  assign new_n934_ = ~new_n543_ & ~new_n932_;
  assign new_n935_ = ~new_n933_ & new_n934_;
  assign new_n936_ = ~new_n212_ & ~new_n829_;
  assign new_n937_ = ~new_n831_ & new_n936_;
  assign o_17_ = ~new_n935_ | ~new_n937_;
  assign new_n939_ = ~new_n878_ & ~new_n880_;
  assign new_n940_ = ~new_n428_ & ~new_n730_;
  assign new_n941_ = ~new_n669_ & new_n940_;
  assign new_n942_ = new_n939_ & new_n941_;
  assign new_n943_ = new_n365_ & new_n406_;
  assign new_n944_ = ~new_n772_ & ~new_n943_;
  assign new_n945_ = ~new_n767_ & new_n944_;
  assign new_n946_ = ~new_n640_ & ~new_n646_;
  assign new_n947_ = ~new_n639_ & new_n946_;
  assign new_n948_ = ~i_53_ & new_n318_;
  assign new_n949_ = new_n406_ & new_n948_;
  assign new_n950_ = ~new_n759_ & ~new_n949_;
  assign new_n951_ = ~new_n432_ & new_n950_;
  assign new_n952_ = new_n945_ & new_n947_;
  assign new_n953_ = new_n951_ & new_n952_;
  assign o_30_ = ~new_n942_ | ~new_n953_;
  assign new_n955_ = new_n302_ & new_n358_;
  assign new_n956_ = ~i_52_ & new_n119_;
  assign new_n957_ = new_n302_ & new_n956_;
  assign new_n958_ = ~new_n488_ & ~new_n955_;
  assign new_n959_ = ~new_n957_ & new_n958_;
  assign o_44_ = new_n839_ | ~new_n959_;
  assign new_n961_ = ~new_n244_ & ~new_n418_;
  assign o_41_ = new_n678_ | ~new_n961_;
  assign new_n963_ = i_34_ & new_n263_;
  assign new_n964_ = new_n687_ & new_n963_;
  assign new_n965_ = ~new_n502_ & ~new_n808_;
  assign new_n966_ = ~new_n688_ & new_n965_;
  assign o_20_ = new_n964_ | ~new_n966_;
  assign new_n968_ = ~i_40_ & new_n263_;
  assign new_n969_ = new_n666_ & new_n968_;
  assign o_47_ = new_n667_ | new_n969_;
  assign new_n971_ = i_47_ & new_n682_;
  assign new_n972_ = ~i_46_ & ~i_43_;
  assign new_n973_ = i_27_ & new_n972_;
  assign new_n974_ = new_n440_ & new_n971_;
  assign new_n975_ = new_n973_ & new_n974_;
  assign o_48_ = ~i_53_ & new_n975_;
  assign new_n977_ = ~new_n340_ & ~new_n580_;
  assign new_n978_ = ~new_n393_ & new_n977_;
  assign o_10_ = ~new_n826_ | ~new_n978_;
  assign o_9_ = new_n323_ | new_n609_;
  assign new_n981_ = new_n356_ & new_n406_;
  assign new_n982_ = ~new_n669_ & ~new_n981_;
  assign new_n983_ = ~new_n244_ & new_n982_;
  assign new_n984_ = ~new_n359_ & ~new_n691_;
  assign new_n985_ = ~new_n759_ & new_n984_;
  assign o_49_ = ~new_n983_ | ~new_n985_;
  assign new_n987_ = ~i_23_ & new_n133_;
  assign new_n988_ = new_n137_ & new_n326_;
  assign new_n989_ = new_n987_ & new_n988_;
  assign new_n990_ = ~new_n290_ & ~new_n529_;
  assign new_n991_ = ~new_n989_ & new_n990_;
  assign new_n992_ = ~i_26_ & new_n133_;
  assign new_n993_ = new_n560_ & new_n992_;
  assign new_n994_ = new_n197_ & new_n560_;
  assign new_n995_ = ~new_n273_ & ~new_n993_;
  assign new_n996_ = ~new_n994_ & new_n995_;
  assign new_n997_ = new_n172_ & new_n178_;
  assign new_n998_ = new_n528_ & new_n997_;
  assign new_n999_ = ~i_0_ & new_n133_;
  assign new_n1000_ = new_n988_ & new_n999_;
  assign new_n1001_ = ~i_32_ & new_n263_;
  assign new_n1002_ = new_n734_ & new_n1001_;
  assign new_n1003_ = ~new_n998_ & ~new_n1000_;
  assign new_n1004_ = ~new_n1002_ & new_n1003_;
  assign new_n1005_ = new_n991_ & new_n996_;
  assign new_n1006_ = new_n1004_ & new_n1005_;
  assign new_n1007_ = i_14_ & new_n108_;
  assign new_n1008_ = new_n173_ & new_n213_;
  assign new_n1009_ = new_n1007_ & new_n1008_;
  assign new_n1010_ = ~new_n412_ & ~new_n1009_;
  assign new_n1011_ = ~new_n253_ & new_n1010_;
  assign new_n1012_ = i_45_ & new_n133_;
  assign new_n1013_ = new_n113_ & new_n214_;
  assign new_n1014_ = new_n1012_ & new_n1013_;
  assign new_n1015_ = ~new_n880_ & ~new_n933_;
  assign new_n1016_ = ~new_n1014_ & new_n1015_;
  assign new_n1017_ = new_n197_ & new_n765_;
  assign new_n1018_ = ~new_n546_ & ~new_n1017_;
  assign new_n1019_ = ~new_n543_ & new_n1018_;
  assign new_n1020_ = i_49_ & i_51_;
  assign new_n1021_ = ~i_48_ & new_n1020_;
  assign new_n1022_ = ~i_20_ & new_n108_;
  assign new_n1023_ = ~i_53_ & new_n1021_;
  assign new_n1024_ = new_n1022_ & new_n1023_;
  assign new_n1025_ = new_n113_ & new_n239_;
  assign new_n1026_ = new_n992_ & new_n1025_;
  assign new_n1027_ = ~new_n287_ & ~new_n1024_;
  assign new_n1028_ = ~new_n1026_ & new_n1027_;
  assign new_n1029_ = new_n1016_ & new_n1019_;
  assign new_n1030_ = new_n1028_ & new_n1029_;
  assign new_n1031_ = new_n1006_ & new_n1011_;
  assign new_n1032_ = new_n1030_ & new_n1031_;
  assign new_n1033_ = i_47_ & new_n112_;
  assign new_n1034_ = i_26_ & ~i_46_;
  assign new_n1035_ = i_1_ & new_n1034_;
  assign new_n1036_ = new_n146_ & new_n1033_;
  assign new_n1037_ = new_n1035_ & new_n1036_;
  assign new_n1038_ = i_48_ & new_n225_;
  assign new_n1039_ = i_5_ & new_n133_;
  assign new_n1040_ = ~i_53_ & new_n1038_;
  assign new_n1041_ = new_n1039_ & new_n1040_;
  assign new_n1042_ = ~i_49_ & new_n326_;
  assign new_n1043_ = ~i_33_ & new_n376_;
  assign new_n1044_ = ~i_53_ & new_n1042_;
  assign new_n1045_ = new_n1043_ & new_n1044_;
  assign new_n1046_ = ~new_n1037_ & ~new_n1041_;
  assign new_n1047_ = ~new_n1045_ & new_n1046_;
  assign new_n1048_ = i_26_ & new_n121_;
  assign new_n1049_ = i_52_ & new_n153_;
  assign new_n1050_ = new_n1048_ & new_n1049_;
  assign new_n1051_ = ~i_50_ & ~i_52_;
  assign new_n1052_ = ~i_49_ & new_n1051_;
  assign new_n1053_ = ~i_29_ & new_n121_;
  assign new_n1054_ = i_53_ & new_n1052_;
  assign new_n1055_ = new_n1053_ & new_n1054_;
  assign new_n1056_ = ~new_n166_ & ~new_n1050_;
  assign new_n1057_ = ~new_n1055_ & new_n1056_;
  assign new_n1058_ = i_49_ & ~i_46_;
  assign new_n1059_ = i_18_ & new_n1058_;
  assign new_n1060_ = new_n384_ & new_n1059_;
  assign new_n1061_ = ~i_49_ & new_n184_;
  assign new_n1062_ = ~i_53_ & new_n1061_;
  assign new_n1063_ = new_n1039_ & new_n1062_;
  assign new_n1064_ = ~new_n1060_ & ~new_n1063_;
  assign new_n1065_ = ~new_n564_ & new_n1064_;
  assign new_n1066_ = new_n1047_ & new_n1057_;
  assign new_n1067_ = new_n1065_ & new_n1066_;
  assign new_n1068_ = ~new_n181_ & ~new_n300_;
  assign new_n1069_ = ~new_n189_ & new_n1068_;
  assign new_n1070_ = i_27_ & new_n108_;
  assign new_n1071_ = i_52_ & new_n137_;
  assign new_n1072_ = new_n1070_ & new_n1071_;
  assign new_n1073_ = new_n179_ & new_n1025_;
  assign new_n1074_ = ~new_n1072_ & ~new_n1073_;
  assign new_n1075_ = ~new_n738_ & new_n1074_;
  assign new_n1076_ = ~i_14_ & new_n263_;
  assign new_n1077_ = new_n178_ & new_n224_;
  assign new_n1078_ = new_n1076_ & new_n1077_;
  assign new_n1079_ = i_2_ & new_n133_;
  assign new_n1080_ = i_52_ & new_n284_;
  assign new_n1081_ = new_n1079_ & new_n1080_;
  assign new_n1082_ = ~new_n662_ & ~new_n1078_;
  assign new_n1083_ = ~new_n1081_ & new_n1082_;
  assign new_n1084_ = new_n1069_ & new_n1075_;
  assign new_n1085_ = new_n1083_ & new_n1084_;
  assign new_n1086_ = i_48_ & new_n105_;
  assign new_n1087_ = i_27_ & new_n133_;
  assign new_n1088_ = new_n162_ & new_n1086_;
  assign new_n1089_ = new_n1087_ & new_n1088_;
  assign new_n1090_ = i_53_ & new_n1042_;
  assign new_n1091_ = new_n122_ & new_n1090_;
  assign new_n1092_ = ~new_n1089_ & ~new_n1091_;
  assign new_n1093_ = ~new_n883_ & new_n1092_;
  assign new_n1094_ = i_3_ & new_n569_;
  assign new_n1095_ = new_n626_ & new_n1094_;
  assign new_n1096_ = ~new_n829_ & ~new_n1095_;
  assign new_n1097_ = ~new_n556_ & new_n1096_;
  assign new_n1098_ = ~new_n141_ & ~new_n568_;
  assign new_n1099_ = ~new_n667_ & new_n1098_;
  assign new_n1100_ = new_n1093_ & new_n1097_;
  assign new_n1101_ = new_n1099_ & new_n1100_;
  assign new_n1102_ = new_n1067_ & new_n1085_;
  assign new_n1103_ = new_n1101_ & new_n1102_;
  assign new_n1104_ = new_n1032_ & new_n1103_;
  assign new_n1105_ = ~o_38_ & ~new_n772_;
  assign new_n1106_ = ~new_n603_ & new_n1105_;
  assign new_n1107_ = ~new_n353_ & ~new_n773_;
  assign new_n1108_ = ~new_n608_ & new_n1107_;
  assign new_n1109_ = ~i_35_ & new_n674_;
  assign new_n1110_ = new_n394_ & new_n1109_;
  assign new_n1111_ = ~new_n369_ & ~new_n1110_;
  assign new_n1112_ = ~new_n767_ & new_n1111_;
  assign new_n1113_ = new_n1106_ & new_n1108_;
  assign new_n1114_ = new_n1112_ & new_n1113_;
  assign new_n1115_ = ~new_n360_ & ~new_n493_;
  assign new_n1116_ = ~new_n496_ & new_n1115_;
  assign new_n1117_ = ~new_n692_ & ~new_n824_;
  assign new_n1118_ = ~new_n357_ & new_n1117_;
  assign new_n1119_ = ~i_45_ & new_n133_;
  assign new_n1120_ = new_n113_ & new_n623_;
  assign new_n1121_ = new_n1119_ & new_n1120_;
  assign new_n1122_ = ~i_8_ & new_n674_;
  assign new_n1123_ = new_n389_ & new_n1122_;
  assign new_n1124_ = ~o_37_ & ~new_n1121_;
  assign new_n1125_ = ~new_n1123_ & new_n1124_;
  assign new_n1126_ = new_n1116_ & new_n1118_;
  assign new_n1127_ = new_n1125_ & new_n1126_;
  assign new_n1128_ = new_n137_ & new_n278_;
  assign new_n1129_ = new_n1076_ & new_n1128_;
  assign new_n1130_ = new_n817_ & ~new_n1129_;
  assign new_n1131_ = ~new_n766_ & ~new_n769_;
  assign new_n1132_ = ~new_n776_ & new_n1131_;
  assign new_n1133_ = ~new_n586_ & ~new_n777_;
  assign new_n1134_ = ~new_n592_ & new_n1133_;
  assign new_n1135_ = new_n1130_ & new_n1132_;
  assign new_n1136_ = new_n1134_ & new_n1135_;
  assign new_n1137_ = new_n1114_ & new_n1127_;
  assign new_n1138_ = new_n1136_ & new_n1137_;
  assign new_n1139_ = ~i_41_ & new_n263_;
  assign new_n1140_ = new_n638_ & new_n1139_;
  assign new_n1141_ = ~new_n652_ & ~o_23_;
  assign new_n1142_ = ~new_n1140_ & new_n1141_;
  assign new_n1143_ = i_49_ & new_n225_;
  assign new_n1144_ = ~i_14_ & new_n674_;
  assign new_n1145_ = ~i_53_ & new_n1143_;
  assign new_n1146_ = new_n1144_ & new_n1145_;
  assign new_n1147_ = ~new_n228_ & ~new_n1146_;
  assign new_n1148_ = ~new_n217_ & new_n1147_;
  assign new_n1149_ = ~new_n212_ & ~o_31_;
  assign new_n1150_ = ~new_n221_ & new_n1149_;
  assign new_n1151_ = new_n1142_ & new_n1148_;
  assign new_n1152_ = new_n1150_ & new_n1151_;
  assign new_n1153_ = ~new_n471_ & ~new_n645_;
  assign new_n1154_ = ~new_n151_ & new_n1153_;
  assign new_n1155_ = ~new_n117_ & ~new_n481_;
  assign new_n1156_ = ~new_n474_ & new_n1155_;
  assign new_n1157_ = ~new_n149_ & ~new_n462_;
  assign new_n1158_ = ~o_14_ & new_n1157_;
  assign new_n1159_ = new_n1154_ & new_n1156_;
  assign new_n1160_ = new_n1158_ & new_n1159_;
  assign new_n1161_ = ~new_n502_ & ~new_n688_;
  assign new_n1162_ = ~new_n420_ & new_n1161_;
  assign new_n1163_ = ~new_n242_ & ~new_n831_;
  assign new_n1164_ = ~new_n238_ & new_n1163_;
  assign new_n1165_ = new_n1162_ & new_n1164_;
  assign new_n1166_ = new_n680_ & new_n1165_;
  assign new_n1167_ = new_n1152_ & new_n1160_;
  assign new_n1168_ = new_n1166_ & new_n1167_;
  assign new_n1169_ = ~new_n340_ & ~new_n787_;
  assign new_n1170_ = ~new_n432_ & new_n1169_;
  assign new_n1171_ = ~new_n342_ & ~new_n949_;
  assign new_n1172_ = ~new_n620_ & new_n1171_;
  assign new_n1173_ = ~new_n388_ & ~o_46_;
  assign new_n1174_ = ~new_n783_ & new_n1173_;
  assign new_n1175_ = new_n1170_ & new_n1172_;
  assign new_n1176_ = new_n1174_ & new_n1175_;
  assign new_n1177_ = ~new_n596_ & ~new_n747_;
  assign new_n1178_ = ~new_n751_ & new_n1177_;
  assign new_n1179_ = ~new_n580_ & ~new_n749_;
  assign new_n1180_ = ~new_n320_ & new_n1179_;
  assign new_n1181_ = ~new_n759_ & ~new_n911_;
  assign new_n1182_ = ~new_n786_ & new_n1181_;
  assign new_n1183_ = new_n1178_ & new_n1180_;
  assign new_n1184_ = new_n1182_ & new_n1183_;
  assign new_n1185_ = ~new_n375_ & ~new_n793_;
  assign new_n1186_ = ~o_42_ & new_n1185_;
  assign new_n1187_ = new_n406_ & new_n684_;
  assign new_n1188_ = ~new_n385_ & ~new_n390_;
  assign new_n1189_ = ~new_n1187_ & new_n1188_;
  assign new_n1190_ = ~new_n393_ & ~o_43_;
  assign new_n1191_ = ~new_n397_ & new_n1190_;
  assign new_n1192_ = new_n1186_ & new_n1189_;
  assign new_n1193_ = new_n1191_ & new_n1192_;
  assign new_n1194_ = new_n1176_ & new_n1184_;
  assign new_n1195_ = new_n1193_ & new_n1194_;
  assign new_n1196_ = new_n1138_ & new_n1168_;
  assign new_n1197_ = new_n1195_ & new_n1196_;
  assign o_7_ = ~new_n1104_ | ~new_n1197_;
  assign new_n1199_ = i_32_ & new_n263_;
  assign new_n1200_ = new_n734_ & new_n1199_;
  assign new_n1201_ = ~new_n714_ & ~new_n1200_;
  assign new_n1202_ = new_n406_ & new_n458_;
  assign new_n1203_ = ~new_n955_ & ~new_n1202_;
  assign new_n1204_ = ~new_n580_ & new_n1203_;
  assign new_n1205_ = ~new_n840_ & ~new_n1002_;
  assign new_n1206_ = ~new_n662_ & new_n1205_;
  assign new_n1207_ = ~new_n390_ & ~new_n793_;
  assign new_n1208_ = ~new_n393_ & new_n1207_;
  assign new_n1209_ = new_n1204_ & new_n1206_;
  assign new_n1210_ = new_n1208_ & new_n1209_;
  assign o_8_ = ~new_n1201_ | ~new_n1210_;
  assign new_n1212_ = ~new_n445_ & ~new_n726_;
  assign new_n1213_ = i_21_ & new_n133_;
  assign new_n1214_ = new_n168_ & new_n196_;
  assign new_n1215_ = new_n1213_ & new_n1214_;
  assign new_n1216_ = ~new_n449_ & ~new_n1200_;
  assign new_n1217_ = ~new_n1215_ & new_n1216_;
  assign new_n1218_ = new_n1212_ & new_n1217_;
  assign new_n1219_ = ~new_n293_ & ~new_n714_;
  assign new_n1220_ = ~new_n998_ & new_n1219_;
  assign new_n1221_ = ~new_n256_ & ~new_n700_;
  assign new_n1222_ = ~new_n705_ & new_n1221_;
  assign new_n1223_ = ~new_n735_ & ~new_n933_;
  assign new_n1224_ = ~new_n518_ & new_n1223_;
  assign new_n1225_ = new_n1220_ & new_n1222_;
  assign new_n1226_ = new_n1224_ & new_n1225_;
  assign new_n1227_ = new_n1218_ & new_n1226_;
  assign new_n1228_ = new_n264_ & new_n473_;
  assign new_n1229_ = ~new_n166_ & ~new_n563_;
  assign new_n1230_ = ~new_n1228_ & new_n1229_;
  assign new_n1231_ = ~new_n170_ & ~new_n189_;
  assign new_n1232_ = ~new_n1078_ & new_n1231_;
  assign new_n1233_ = i_12_ & new_n1058_;
  assign new_n1234_ = ~i_53_ & new_n440_;
  assign new_n1235_ = new_n1233_ & new_n1234_;
  assign new_n1236_ = ~new_n175_ & ~new_n1037_;
  assign new_n1237_ = ~new_n1235_ & new_n1236_;
  assign new_n1238_ = new_n1230_ & new_n1232_;
  assign new_n1239_ = new_n1237_ & new_n1238_;
  assign new_n1240_ = ~new_n415_ & ~new_n426_;
  assign new_n1241_ = ~o_29_ & new_n1240_;
  assign new_n1242_ = ~i_48_ & new_n218_;
  assign new_n1243_ = ~i_36_ & new_n108_;
  assign new_n1244_ = i_52_ & new_n1242_;
  assign new_n1245_ = new_n1243_ & new_n1244_;
  assign new_n1246_ = ~new_n287_ & ~new_n730_;
  assign new_n1247_ = ~new_n1245_ & new_n1246_;
  assign new_n1248_ = ~new_n300_ & ~new_n424_;
  assign new_n1249_ = ~new_n181_ & new_n1248_;
  assign new_n1250_ = new_n1241_ & new_n1247_;
  assign new_n1251_ = new_n1249_ & new_n1250_;
  assign new_n1252_ = ~new_n204_ & ~new_n554_;
  assign new_n1253_ = ~new_n557_ & new_n1252_;
  assign new_n1254_ = ~new_n195_ & ~new_n564_;
  assign new_n1255_ = ~new_n874_ & new_n1254_;
  assign new_n1256_ = ~new_n883_ & ~new_n1089_;
  assign new_n1257_ = ~new_n568_ & new_n1256_;
  assign new_n1258_ = new_n1253_ & new_n1255_;
  assign new_n1259_ = new_n1257_ & new_n1258_;
  assign new_n1260_ = new_n1239_ & new_n1251_;
  assign new_n1261_ = new_n1259_ & new_n1260_;
  assign new_n1262_ = new_n1227_ & new_n1261_;
  assign new_n1263_ = ~new_n350_ & ~new_n773_;
  assign new_n1264_ = ~new_n609_ & new_n1263_;
  assign new_n1265_ = ~new_n357_ & ~new_n496_;
  assign new_n1266_ = ~new_n1121_ & new_n1265_;
  assign new_n1267_ = ~new_n364_ & ~new_n612_;
  assign new_n1268_ = ~new_n1110_ & new_n1267_;
  assign new_n1269_ = new_n1264_ & new_n1266_;
  assign new_n1270_ = new_n1268_ & new_n1269_;
  assign new_n1271_ = ~new_n420_ & ~new_n825_;
  assign new_n1272_ = ~o_36_ & new_n1271_;
  assign new_n1273_ = ~new_n359_ & new_n1161_;
  assign new_n1274_ = ~new_n676_ & ~new_n692_;
  assign new_n1275_ = ~new_n824_ & new_n1274_;
  assign new_n1276_ = new_n1272_ & new_n1273_;
  assign new_n1277_ = new_n1275_ & new_n1276_;
  assign new_n1278_ = ~i_50_ & i_47_;
  assign new_n1279_ = ~i_46_ & new_n1278_;
  assign new_n1280_ = new_n239_ & new_n1279_;
  assign new_n1281_ = ~new_n1129_ & ~new_n1280_;
  assign new_n1282_ = ~new_n777_ & new_n1281_;
  assign new_n1283_ = ~new_n589_ & ~new_n592_;
  assign new_n1284_ = ~new_n580_ & new_n1283_;
  assign new_n1285_ = new_n1132_ & new_n1282_;
  assign new_n1286_ = new_n1284_ & new_n1285_;
  assign new_n1287_ = new_n1270_ & new_n1277_;
  assign new_n1288_ = new_n1286_ & new_n1287_;
  assign new_n1289_ = ~new_n157_ & ~new_n639_;
  assign new_n1290_ = ~new_n230_ & new_n1289_;
  assign new_n1291_ = ~i_44_ & new_n263_;
  assign new_n1292_ = new_n198_ & new_n1291_;
  assign new_n1293_ = ~new_n462_ & ~new_n488_;
  assign new_n1294_ = ~new_n1292_ & new_n1293_;
  assign new_n1295_ = new_n335_ & new_n406_;
  assign new_n1296_ = new_n322_ & new_n482_;
  assign new_n1297_ = ~new_n1295_ & ~new_n1296_;
  assign new_n1298_ = ~new_n465_ & new_n1297_;
  assign new_n1299_ = new_n1290_ & new_n1294_;
  assign new_n1300_ = new_n1298_ & new_n1299_;
  assign new_n1301_ = ~new_n669_ & new_n1155_;
  assign new_n1302_ = i_48_ & new_n118_;
  assign new_n1303_ = new_n120_ & new_n1302_;
  assign new_n1304_ = new_n150_ & new_n1303_;
  assign new_n1305_ = ~new_n419_ & ~new_n484_;
  assign new_n1306_ = ~new_n1304_ & new_n1305_;
  assign new_n1307_ = ~new_n418_ & ~new_n645_;
  assign new_n1308_ = ~new_n477_ & new_n1307_;
  assign new_n1309_ = new_n1301_ & new_n1306_;
  assign new_n1310_ = new_n1308_ & new_n1309_;
  assign new_n1311_ = ~o_31_ & ~new_n981_;
  assign new_n1312_ = ~new_n831_ & new_n1311_;
  assign new_n1313_ = ~new_n814_ & ~new_n1140_;
  assign new_n1314_ = ~new_n212_ & new_n1313_;
  assign new_n1315_ = ~new_n242_ & ~new_n244_;
  assign new_n1316_ = ~new_n685_ & new_n1315_;
  assign new_n1317_ = new_n1312_ & new_n1314_;
  assign new_n1318_ = new_n1316_ & new_n1317_;
  assign new_n1319_ = new_n1300_ & new_n1310_;
  assign new_n1320_ = new_n1318_ & new_n1319_;
  assign new_n1321_ = ~new_n342_ & ~new_n620_;
  assign new_n1322_ = ~new_n787_ & new_n1321_;
  assign new_n1323_ = ~new_n597_ & ~new_n759_;
  assign new_n1324_ = ~new_n786_ & new_n1323_;
  assign new_n1325_ = new_n1322_ & new_n1324_;
  assign new_n1326_ = new_n785_ & new_n1325_;
  assign new_n1327_ = new_n377_ & new_n948_;
  assign new_n1328_ = ~new_n751_ & ~new_n1327_;
  assign new_n1329_ = ~new_n911_ & new_n1328_;
  assign new_n1330_ = ~new_n583_ & ~new_n596_;
  assign new_n1331_ = ~new_n747_ & new_n1330_;
  assign new_n1332_ = ~new_n323_ & new_n760_;
  assign new_n1333_ = new_n1329_ & new_n1331_;
  assign new_n1334_ = new_n1332_ & new_n1333_;
  assign new_n1335_ = ~new_n375_ & ~o_42_;
  assign new_n1336_ = ~o_43_ & new_n1335_;
  assign new_n1337_ = ~new_n793_ & ~new_n1187_;
  assign new_n1338_ = ~new_n378_ & new_n1337_;
  assign new_n1339_ = ~o_33_ & ~new_n627_;
  assign new_n1340_ = ~new_n397_ & new_n1339_;
  assign new_n1341_ = new_n1336_ & new_n1338_;
  assign new_n1342_ = new_n1340_ & new_n1341_;
  assign new_n1343_ = new_n1326_ & new_n1334_;
  assign new_n1344_ = new_n1342_ & new_n1343_;
  assign new_n1345_ = new_n1288_ & new_n1320_;
  assign new_n1346_ = new_n1344_ & new_n1345_;
  assign o_5_ = ~new_n1262_ | ~new_n1346_;
  assign new_n1348_ = ~new_n271_ & ~new_n705_;
  assign new_n1349_ = ~new_n714_ & new_n1348_;
  assign new_n1350_ = ~new_n709_ & ~new_n1215_;
  assign new_n1351_ = ~new_n700_ & new_n1350_;
  assign new_n1352_ = i_53_ & ~i_51_;
  assign new_n1353_ = ~i_15_ & new_n263_;
  assign new_n1354_ = new_n145_ & new_n1352_;
  assign new_n1355_ = new_n1353_ & new_n1354_;
  assign new_n1356_ = ~new_n878_ & ~new_n1355_;
  assign new_n1357_ = ~new_n1002_ & new_n1356_;
  assign new_n1358_ = new_n1349_ & new_n1351_;
  assign new_n1359_ = new_n1357_ & new_n1358_;
  assign new_n1360_ = ~new_n262_ & ~new_n964_;
  assign new_n1361_ = ~new_n1009_ & new_n1360_;
  assign new_n1362_ = new_n727_ & new_n1361_;
  assign new_n1363_ = ~i_48_ & new_n379_;
  assign new_n1364_ = new_n162_ & new_n1363_;
  assign new_n1365_ = new_n872_ & new_n1364_;
  assign new_n1366_ = ~new_n548_ & ~new_n1365_;
  assign new_n1367_ = ~new_n1014_ & new_n1366_;
  assign new_n1368_ = ~i_48_ & new_n200_;
  assign new_n1369_ = i_36_ & new_n108_;
  assign new_n1370_ = ~i_53_ & new_n1368_;
  assign new_n1371_ = new_n1369_ & new_n1370_;
  assign new_n1372_ = ~new_n297_ & ~new_n543_;
  assign new_n1373_ = ~new_n1371_ & new_n1372_;
  assign new_n1374_ = i_49_ & ~i_52_;
  assign new_n1375_ = i_48_ & new_n1374_;
  assign new_n1376_ = i_53_ & new_n1375_;
  assign new_n1377_ = new_n147_ & new_n1376_;
  assign new_n1378_ = ~new_n730_ & ~new_n1026_;
  assign new_n1379_ = ~new_n1377_ & new_n1378_;
  assign new_n1380_ = new_n1367_ & new_n1373_;
  assign new_n1381_ = new_n1379_ & new_n1380_;
  assign new_n1382_ = new_n1359_ & new_n1362_;
  assign new_n1383_ = new_n1381_ & new_n1382_;
  assign new_n1384_ = ~new_n502_ & ~new_n943_;
  assign new_n1385_ = ~new_n678_ & new_n1384_;
  assign new_n1386_ = ~new_n831_ & ~new_n981_;
  assign new_n1387_ = ~new_n238_ & new_n1386_;
  assign new_n1388_ = ~new_n351_ & ~new_n357_;
  assign new_n1389_ = ~new_n691_ & new_n1388_;
  assign new_n1390_ = new_n1385_ & new_n1387_;
  assign new_n1391_ = new_n1389_ & new_n1390_;
  assign new_n1392_ = ~new_n459_ & ~new_n649_;
  assign new_n1393_ = ~new_n228_ & new_n1392_;
  assign new_n1394_ = ~new_n124_ & ~new_n471_;
  assign new_n1395_ = ~new_n1292_ & new_n1394_;
  assign new_n1396_ = ~new_n217_ & ~new_n1146_;
  assign new_n1397_ = ~new_n465_ & new_n1396_;
  assign new_n1398_ = new_n1393_ & new_n1395_;
  assign new_n1399_ = new_n1397_ & new_n1398_;
  assign new_n1400_ = ~new_n773_ & ~new_n1123_;
  assign new_n1401_ = ~new_n608_ & new_n1400_;
  assign new_n1402_ = ~new_n493_ & ~new_n1121_;
  assign new_n1403_ = ~new_n507_ & new_n1402_;
  assign new_n1404_ = ~new_n609_ & ~new_n772_;
  assign new_n1405_ = ~new_n366_ & new_n1404_;
  assign new_n1406_ = new_n1401_ & new_n1403_;
  assign new_n1407_ = new_n1405_ & new_n1406_;
  assign new_n1408_ = new_n1391_ & new_n1399_;
  assign new_n1409_ = new_n1407_ & new_n1408_;
  assign new_n1410_ = ~new_n554_ & ~new_n557_;
  assign new_n1411_ = ~new_n1089_ & new_n1410_;
  assign new_n1412_ = ~new_n556_ & ~new_n829_;
  assign new_n1413_ = ~new_n874_ & new_n1412_;
  assign new_n1414_ = ~new_n571_ & ~new_n668_;
  assign new_n1415_ = ~new_n568_ & new_n1414_;
  assign new_n1416_ = new_n1411_ & new_n1413_;
  assign new_n1417_ = new_n1415_ & new_n1416_;
  assign new_n1418_ = ~new_n662_ & ~new_n1228_;
  assign new_n1419_ = ~new_n199_ & new_n1418_;
  assign new_n1420_ = ~new_n188_ & ~new_n1073_;
  assign new_n1421_ = ~new_n1078_ & new_n1420_;
  assign new_n1422_ = i_25_ & new_n674_;
  assign new_n1423_ = new_n894_ & new_n1422_;
  assign new_n1424_ = ~new_n195_ & ~new_n1423_;
  assign new_n1425_ = ~new_n564_ & new_n1424_;
  assign new_n1426_ = new_n1419_ & new_n1421_;
  assign new_n1427_ = new_n1425_ & new_n1426_;
  assign new_n1428_ = ~o_27_ & new_n1155_;
  assign new_n1429_ = ~new_n573_ & ~new_n1304_;
  assign new_n1430_ = ~new_n667_ & new_n1429_;
  assign new_n1431_ = ~new_n111_ & ~new_n474_;
  assign new_n1432_ = ~new_n645_ & new_n1431_;
  assign new_n1433_ = new_n1428_ & new_n1430_;
  assign new_n1434_ = new_n1432_ & new_n1433_;
  assign new_n1435_ = new_n1417_ & new_n1427_;
  assign new_n1436_ = new_n1434_ & new_n1435_;
  assign new_n1437_ = ~new_n320_ & ~new_n596_;
  assign new_n1438_ = ~new_n316_ & new_n1437_;
  assign new_n1439_ = ~new_n582_ & ~new_n592_;
  assign new_n1440_ = ~new_n583_ & new_n1439_;
  assign new_n1441_ = ~new_n756_ & ~new_n911_;
  assign new_n1442_ = ~new_n759_ & new_n1441_;
  assign new_n1443_ = new_n1438_ & new_n1440_;
  assign new_n1444_ = new_n1442_ & new_n1443_;
  assign new_n1445_ = ~new_n329_ & ~new_n1202_;
  assign new_n1446_ = ~new_n336_ & new_n1445_;
  assign new_n1447_ = ~new_n364_ & ~new_n369_;
  assign new_n1448_ = ~new_n334_ & new_n1447_;
  assign new_n1449_ = ~new_n589_ & ~new_n1129_;
  assign new_n1450_ = ~new_n586_ & new_n1449_;
  assign new_n1451_ = new_n1446_ & new_n1448_;
  assign new_n1452_ = new_n1450_ & new_n1451_;
  assign new_n1453_ = new_n381_ & ~o_33_;
  assign new_n1454_ = ~new_n388_ & ~new_n620_;
  assign new_n1455_ = ~new_n390_ & new_n1454_;
  assign new_n1456_ = ~new_n393_ & ~new_n627_;
  assign new_n1457_ = ~new_n397_ & new_n1456_;
  assign new_n1458_ = new_n1453_ & new_n1455_;
  assign new_n1459_ = new_n1457_ & new_n1458_;
  assign new_n1460_ = new_n1444_ & new_n1452_;
  assign new_n1461_ = new_n1459_ & new_n1460_;
  assign new_n1462_ = new_n1409_ & new_n1436_;
  assign new_n1463_ = new_n1461_ & new_n1462_;
  assign o_6_ = ~new_n1383_ | ~new_n1463_;
  assign new_n1465_ = new_n197_ & new_n1303_;
  assign new_n1466_ = ~new_n293_ & ~new_n1465_;
  assign new_n1467_ = ~new_n808_ & new_n1466_;
  assign new_n1468_ = ~new_n878_ & ~new_n969_;
  assign new_n1469_ = ~new_n880_ & new_n1468_;
  assign new_n1470_ = new_n275_ & new_n1467_;
  assign new_n1471_ = new_n1469_ & new_n1470_;
  assign new_n1472_ = ~new_n412_ & new_n1471_;
  assign new_n1473_ = new_n176_ & ~new_n1228_;
  assign new_n1474_ = ~new_n188_ & new_n429_;
  assign new_n1475_ = ~new_n175_ & ~new_n657_;
  assign new_n1476_ = ~new_n199_ & new_n1475_;
  assign new_n1477_ = new_n1473_ & new_n1474_;
  assign new_n1478_ = new_n1476_ & new_n1477_;
  assign new_n1479_ = ~new_n521_ & ~new_n730_;
  assign new_n1480_ = ~new_n1026_ & new_n1479_;
  assign new_n1481_ = ~new_n283_ & ~new_n890_;
  assign new_n1482_ = ~new_n1014_ & new_n1481_;
  assign new_n1483_ = ~new_n823_ & ~new_n1073_;
  assign new_n1484_ = ~new_n415_ & new_n1483_;
  assign new_n1485_ = new_n1480_ & new_n1482_;
  assign new_n1486_ = new_n1484_ & new_n1485_;
  assign new_n1487_ = ~new_n556_ & ~o_13_;
  assign new_n1488_ = ~new_n136_ & new_n1487_;
  assign new_n1489_ = new_n107_ & new_n153_;
  assign new_n1490_ = new_n122_ & new_n1489_;
  assign new_n1491_ = ~new_n829_ & ~new_n1490_;
  assign new_n1492_ = ~new_n428_ & new_n1491_;
  assign new_n1493_ = ~new_n131_ & ~new_n668_;
  assign new_n1494_ = ~new_n484_ & new_n1493_;
  assign new_n1495_ = new_n1488_ & new_n1492_;
  assign new_n1496_ = new_n1494_ & new_n1495_;
  assign new_n1497_ = new_n1478_ & new_n1486_;
  assign new_n1498_ = new_n1496_ & new_n1497_;
  assign new_n1499_ = new_n1472_ & new_n1498_;
  assign new_n1500_ = ~new_n334_ & ~new_n369_;
  assign new_n1501_ = ~new_n1110_ & new_n1500_;
  assign new_n1502_ = ~new_n364_ & new_n1105_;
  assign new_n1503_ = new_n1501_ & new_n1502_;
  assign new_n1504_ = new_n771_ & new_n1503_;
  assign new_n1505_ = ~new_n351_ & ~new_n691_;
  assign new_n1506_ = ~new_n496_ & new_n1505_;
  assign new_n1507_ = ~o_36_ & ~new_n678_;
  assign new_n1508_ = ~new_n360_ & new_n1507_;
  assign new_n1509_ = ~o_37_ & ~new_n1123_;
  assign new_n1510_ = ~new_n353_ & new_n1509_;
  assign new_n1511_ = new_n1506_ & new_n1508_;
  assign new_n1512_ = new_n1510_ & new_n1511_;
  assign new_n1513_ = i_50_ & i_48_;
  assign new_n1514_ = ~i_46_ & new_n1513_;
  assign new_n1515_ = new_n209_ & new_n1514_;
  assign new_n1516_ = ~new_n336_ & ~new_n1129_;
  assign new_n1517_ = ~new_n1515_ & new_n1516_;
  assign new_n1518_ = ~new_n776_ & new_n1445_;
  assign new_n1519_ = ~new_n582_ & new_n1283_;
  assign new_n1520_ = new_n1517_ & new_n1518_;
  assign new_n1521_ = new_n1519_ & new_n1520_;
  assign new_n1522_ = new_n1504_ & new_n1512_;
  assign new_n1523_ = new_n1521_ & new_n1522_;
  assign new_n1524_ = ~i_30_ & new_n1058_;
  assign new_n1525_ = new_n626_ & new_n1524_;
  assign new_n1526_ = ~new_n232_ & ~new_n1525_;
  assign new_n1527_ = ~new_n217_ & new_n1526_;
  assign new_n1528_ = ~new_n228_ & ~new_n1296_;
  assign new_n1529_ = ~new_n1295_ & new_n1528_;
  assign new_n1530_ = ~new_n652_ & ~new_n1140_;
  assign new_n1531_ = ~new_n212_ & new_n1530_;
  assign new_n1532_ = new_n1527_ & new_n1529_;
  assign new_n1533_ = new_n1531_ & new_n1532_;
  assign new_n1534_ = ~new_n151_ & ~new_n646_;
  assign new_n1535_ = ~new_n149_ & new_n1534_;
  assign new_n1536_ = ~new_n117_ & ~new_n669_;
  assign new_n1537_ = ~new_n111_ & new_n1536_;
  assign new_n1538_ = ~new_n640_ & ~new_n1292_;
  assign new_n1539_ = ~new_n639_ & new_n1538_;
  assign new_n1540_ = new_n1535_ & new_n1537_;
  assign new_n1541_ = new_n1539_ & new_n1540_;
  assign new_n1542_ = i_48_ & new_n317_;
  assign new_n1543_ = ~i_8_ & new_n263_;
  assign new_n1544_ = ~i_53_ & new_n1542_;
  assign new_n1545_ = new_n1543_ & new_n1544_;
  assign new_n1546_ = ~new_n502_ & ~new_n1545_;
  assign new_n1547_ = ~new_n688_ & new_n1546_;
  assign new_n1548_ = i_53_ & new_n1542_;
  assign new_n1549_ = new_n475_ & new_n1548_;
  assign new_n1550_ = ~new_n242_ & ~new_n955_;
  assign new_n1551_ = ~new_n1549_ & new_n1550_;
  assign new_n1552_ = ~i_52_ & new_n301_;
  assign new_n1553_ = new_n377_ & new_n1552_;
  assign new_n1554_ = ~i_46_ & new_n892_;
  assign new_n1555_ = i_53_ & new_n624_;
  assign new_n1556_ = new_n1554_ & new_n1555_;
  assign new_n1557_ = ~new_n1553_ & ~new_n1556_;
  assign new_n1558_ = ~new_n677_ & new_n1557_;
  assign new_n1559_ = new_n1547_ & new_n1551_;
  assign new_n1560_ = new_n1558_ & new_n1559_;
  assign new_n1561_ = new_n1533_ & new_n1541_;
  assign new_n1562_ = new_n1560_ & new_n1561_;
  assign new_n1563_ = ~new_n345_ & new_n1169_;
  assign new_n1564_ = new_n1324_ & new_n1563_;
  assign new_n1565_ = new_n785_ & new_n1564_;
  assign new_n1566_ = ~new_n911_ & ~new_n1327_;
  assign new_n1567_ = ~new_n758_ & new_n1566_;
  assign new_n1568_ = ~new_n756_ & ~new_n957_;
  assign new_n1569_ = ~new_n323_ & new_n1568_;
  assign new_n1570_ = new_n1178_ & new_n1567_;
  assign new_n1571_ = new_n1569_ & new_n1570_;
  assign new_n1572_ = ~i_46_ & new_n171_;
  assign new_n1573_ = new_n114_ & new_n1572_;
  assign new_n1574_ = ~new_n390_ & ~new_n1573_;
  assign new_n1575_ = ~new_n378_ & new_n1574_;
  assign new_n1576_ = new_n1336_ & new_n1575_;
  assign new_n1577_ = new_n399_ & new_n1576_;
  assign new_n1578_ = new_n1565_ & new_n1571_;
  assign new_n1579_ = new_n1577_ & new_n1578_;
  assign new_n1580_ = new_n1523_ & new_n1562_;
  assign new_n1581_ = new_n1579_ & new_n1580_;
  assign o_3_ = ~new_n1499_ | ~new_n1581_;
  assign new_n1583_ = new_n107_ & new_n1363_;
  assign new_n1584_ = new_n236_ & new_n1583_;
  assign new_n1585_ = ~new_n717_ & ~new_n1584_;
  assign new_n1586_ = ~new_n969_ & new_n1585_;
  assign new_n1587_ = ~new_n271_ & ~new_n539_;
  assign new_n1588_ = ~new_n808_ & new_n1587_;
  assign new_n1589_ = ~new_n735_ & ~new_n890_;
  assign new_n1590_ = ~new_n548_ & new_n1589_;
  assign new_n1591_ = new_n1586_ & new_n1588_;
  assign new_n1592_ = new_n1590_ & new_n1591_;
  assign new_n1593_ = new_n727_ & ~new_n932_;
  assign new_n1594_ = new_n288_ & ~new_n521_;
  assign new_n1595_ = ~new_n424_ & ~new_n563_;
  assign new_n1596_ = ~new_n662_ & new_n1595_;
  assign new_n1597_ = new_n740_ & new_n1594_;
  assign new_n1598_ = new_n1596_ & new_n1597_;
  assign new_n1599_ = new_n1592_ & new_n1593_;
  assign new_n1600_ = new_n1598_ & new_n1599_;
  assign new_n1601_ = i_14_ & new_n674_;
  assign new_n1602_ = new_n956_ & new_n1601_;
  assign new_n1603_ = ~new_n141_ & ~new_n1602_;
  assign new_n1604_ = ~new_n573_ & new_n1603_;
  assign new_n1605_ = ~new_n557_ & ~new_n839_;
  assign new_n1606_ = ~new_n883_ & new_n1605_;
  assign new_n1607_ = ~new_n667_ & ~new_n1304_;
  assign new_n1608_ = ~new_n474_ & new_n1607_;
  assign new_n1609_ = new_n1604_ & new_n1606_;
  assign new_n1610_ = new_n1608_ & new_n1609_;
  assign new_n1611_ = ~i_27_ & new_n133_;
  assign new_n1612_ = i_52_ & new_n106_;
  assign new_n1613_ = new_n1611_ & new_n1612_;
  assign new_n1614_ = ~new_n175_ & ~new_n1613_;
  assign new_n1615_ = ~new_n199_ & new_n1614_;
  assign new_n1616_ = ~i_21_ & new_n133_;
  assign new_n1617_ = i_53_ & new_n1086_;
  assign new_n1618_ = new_n1616_ & new_n1617_;
  assign new_n1619_ = ~new_n561_ & ~new_n1618_;
  assign new_n1620_ = ~new_n1037_ & new_n1619_;
  assign new_n1621_ = ~new_n874_ & ~new_n1490_;
  assign new_n1622_ = ~new_n554_ & new_n1621_;
  assign new_n1623_ = new_n1615_ & new_n1620_;
  assign new_n1624_ = new_n1622_ & new_n1623_;
  assign new_n1625_ = ~new_n124_ & ~new_n418_;
  assign new_n1626_ = ~new_n646_ & new_n1625_;
  assign new_n1627_ = ~new_n111_ & ~new_n645_;
  assign new_n1628_ = ~new_n471_ & new_n1627_;
  assign new_n1629_ = ~new_n462_ & ~new_n477_;
  assign new_n1630_ = ~new_n640_ & new_n1629_;
  assign new_n1631_ = new_n1626_ & new_n1628_;
  assign new_n1632_ = new_n1630_ & new_n1631_;
  assign new_n1633_ = new_n1610_ & new_n1624_;
  assign new_n1634_ = new_n1632_ & new_n1633_;
  assign new_n1635_ = new_n1600_ & new_n1634_;
  assign new_n1636_ = ~new_n769_ & ~new_n1202_;
  assign new_n1637_ = ~new_n776_ & new_n1636_;
  assign new_n1638_ = ~new_n767_ & ~new_n1110_;
  assign new_n1639_ = ~new_n766_ & new_n1638_;
  assign new_n1640_ = ~new_n613_ & ~new_n777_;
  assign new_n1641_ = ~new_n589_ & new_n1640_;
  assign new_n1642_ = new_n1637_ & new_n1639_;
  assign new_n1643_ = new_n1641_ & new_n1642_;
  assign new_n1644_ = new_n113_ & new_n482_;
  assign new_n1645_ = ~new_n1123_ & ~new_n1644_;
  assign new_n1646_ = ~new_n603_ & new_n1645_;
  assign new_n1647_ = ~new_n507_ & ~new_n1121_;
  assign new_n1648_ = ~new_n350_ & new_n1647_;
  assign new_n1649_ = ~new_n366_ & ~new_n612_;
  assign new_n1650_ = ~new_n369_ & new_n1649_;
  assign new_n1651_ = new_n1646_ & new_n1648_;
  assign new_n1652_ = new_n1650_ & new_n1651_;
  assign new_n1653_ = ~new_n747_ & new_n1437_;
  assign new_n1654_ = ~new_n586_ & ~new_n592_;
  assign new_n1655_ = ~new_n583_ & new_n1654_;
  assign new_n1656_ = ~new_n316_ & ~new_n751_;
  assign new_n1657_ = ~new_n1327_ & new_n1656_;
  assign new_n1658_ = new_n1653_ & new_n1655_;
  assign new_n1659_ = new_n1657_ & new_n1658_;
  assign new_n1660_ = new_n1643_ & new_n1652_;
  assign new_n1661_ = new_n1659_ & new_n1660_;
  assign new_n1662_ = ~new_n955_ & ~new_n1549_;
  assign new_n1663_ = ~new_n1545_ & new_n1662_;
  assign new_n1664_ = ~new_n212_ & ~new_n831_;
  assign new_n1665_ = ~new_n242_ & new_n1664_;
  assign new_n1666_ = ~new_n244_ & ~new_n943_;
  assign new_n1667_ = ~new_n688_ & new_n1666_;
  assign new_n1668_ = new_n1663_ & new_n1665_;
  assign new_n1669_ = new_n1667_ & new_n1668_;
  assign new_n1670_ = ~new_n230_ & ~new_n1296_;
  assign new_n1671_ = ~new_n232_ & new_n1670_;
  assign new_n1672_ = ~new_n639_ & ~new_n1292_;
  assign new_n1673_ = ~new_n649_ & new_n1672_;
  assign new_n1674_ = ~new_n453_ & ~new_n1525_;
  assign new_n1675_ = ~new_n217_ & new_n1674_;
  assign new_n1676_ = new_n1671_ & new_n1673_;
  assign new_n1677_ = new_n1675_ & new_n1676_;
  assign new_n1678_ = ~new_n504_ & ~new_n676_;
  assign new_n1679_ = ~new_n360_ & new_n1678_;
  assign new_n1680_ = ~new_n359_ & ~new_n825_;
  assign new_n1681_ = ~new_n1553_ & new_n1680_;
  assign new_n1682_ = ~new_n493_ & ~new_n691_;
  assign new_n1683_ = ~new_n496_ & new_n1682_;
  assign new_n1684_ = new_n1679_ & new_n1681_;
  assign new_n1685_ = new_n1683_ & new_n1684_;
  assign new_n1686_ = new_n1669_ & new_n1677_;
  assign new_n1687_ = new_n1685_ & new_n1686_;
  assign new_n1688_ = new_n1188_ & ~new_n1573_;
  assign new_n1689_ = new_n785_ & new_n1563_;
  assign new_n1690_ = new_n1688_ & new_n1689_;
  assign new_n1691_ = ~new_n323_ & ~new_n957_;
  assign new_n1692_ = ~new_n597_ & new_n1691_;
  assign new_n1693_ = ~new_n758_ & ~new_n911_;
  assign new_n1694_ = ~new_n756_ & new_n1693_;
  assign new_n1695_ = ~new_n786_ & ~new_n949_;
  assign new_n1696_ = ~new_n342_ & new_n1695_;
  assign new_n1697_ = new_n1692_ & new_n1694_;
  assign new_n1698_ = new_n1696_ & new_n1697_;
  assign new_n1699_ = ~o_42_ & ~o_43_;
  assign new_n1700_ = ~o_33_ & new_n1699_;
  assign new_n1701_ = new_n1338_ & new_n1700_;
  assign new_n1702_ = new_n1457_ & new_n1701_;
  assign new_n1703_ = new_n1690_ & new_n1698_;
  assign new_n1704_ = new_n1702_ & new_n1703_;
  assign new_n1705_ = new_n1661_ & new_n1687_;
  assign new_n1706_ = new_n1704_ & new_n1705_;
  assign o_4_ = ~new_n1635_ | ~new_n1706_;
  assign o_45_ = o_31_;
endmodule

