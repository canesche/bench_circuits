// Benchmark "top" written by ABC on Thu Oct  8 22:51:57 2020

module top ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \b[0] ,
    \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] , \b[17] ,
    \b[18] , \b[19] , \b[20] , \b[21] , \b[22] , \b[23] , \b[24] , \b[25] ,
    \b[26] , \b[27] , \b[28] , \b[29] , \b[30] , \b[31] , \b[32] , \b[33] ,
    \b[34] , \b[35] , \b[36] , \b[37] , \b[38] , \b[39] , \b[40] , \b[41] ,
    \b[42] , \b[43] , \b[44] , \b[45] , \b[46] , \b[47] , \b[48] , \b[49] ,
    \b[50] , \b[51] , \b[52] , \b[53] , \b[54] , \b[55] , \b[56] , \b[57] ,
    \b[58] , \b[59] , \b[60] , \b[61] , \b[62] , \b[63] ,
    \quotient[0] , \quotient[1] , \quotient[2] , \quotient[3] ,
    \quotient[4] , \quotient[5] , \quotient[6] , \quotient[7] ,
    \quotient[8] , \quotient[9] , \quotient[10] , \quotient[11] ,
    \quotient[12] , \quotient[13] , \quotient[14] , \quotient[15] ,
    \quotient[16] , \quotient[17] , \quotient[18] , \quotient[19] ,
    \quotient[20] , \quotient[21] , \quotient[22] , \quotient[23] ,
    \quotient[24] , \quotient[25] , \quotient[26] , \quotient[27] ,
    \quotient[28] , \quotient[29] , \quotient[30] , \quotient[31] ,
    \quotient[32] , \quotient[33] , \quotient[34] , \quotient[35] ,
    \quotient[36] , \quotient[37] , \quotient[38] , \quotient[39] ,
    \quotient[40] , \quotient[41] , \quotient[42] , \quotient[43] ,
    \quotient[44] , \quotient[45] , \quotient[46] , \quotient[47] ,
    \quotient[48] , \quotient[49] , \quotient[50] , \quotient[51] ,
    \quotient[52] , \quotient[53] , \quotient[54] , \quotient[55] ,
    \quotient[56] , \quotient[57] , \quotient[58] , \quotient[59] ,
    \quotient[60] , \quotient[61] , \quotient[62] , \quotient[63] ,
    \remainder[0] , \remainder[1] , \remainder[2] , \remainder[3] ,
    \remainder[4] , \remainder[5] , \remainder[6] , \remainder[7] ,
    \remainder[8] , \remainder[9] , \remainder[10] , \remainder[11] ,
    \remainder[12] , \remainder[13] , \remainder[14] , \remainder[15] ,
    \remainder[16] , \remainder[17] , \remainder[18] , \remainder[19] ,
    \remainder[20] , \remainder[21] , \remainder[22] , \remainder[23] ,
    \remainder[24] , \remainder[25] , \remainder[26] , \remainder[27] ,
    \remainder[28] , \remainder[29] , \remainder[30] , \remainder[31] ,
    \remainder[32] , \remainder[33] , \remainder[34] , \remainder[35] ,
    \remainder[36] , \remainder[37] , \remainder[38] , \remainder[39] ,
    \remainder[40] , \remainder[41] , \remainder[42] , \remainder[43] ,
    \remainder[44] , \remainder[45] , \remainder[46] , \remainder[47] ,
    \remainder[48] , \remainder[49] , \remainder[50] , \remainder[51] ,
    \remainder[52] , \remainder[53] , \remainder[54] , \remainder[55] ,
    \remainder[56] , \remainder[57] , \remainder[58] , \remainder[59] ,
    \remainder[60] , \remainder[61] , \remainder[62] , \remainder[63]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \b[0] , \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] ,
    \b[9] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[20] , \b[21] , \b[22] , \b[23] , \b[24] ,
    \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[30] , \b[31] , \b[32] ,
    \b[33] , \b[34] , \b[35] , \b[36] , \b[37] , \b[38] , \b[39] , \b[40] ,
    \b[41] , \b[42] , \b[43] , \b[44] , \b[45] , \b[46] , \b[47] , \b[48] ,
    \b[49] , \b[50] , \b[51] , \b[52] , \b[53] , \b[54] , \b[55] , \b[56] ,
    \b[57] , \b[58] , \b[59] , \b[60] , \b[61] , \b[62] , \b[63] ;
  output \quotient[0] , \quotient[1] , \quotient[2] , \quotient[3] ,
    \quotient[4] , \quotient[5] , \quotient[6] , \quotient[7] ,
    \quotient[8] , \quotient[9] , \quotient[10] , \quotient[11] ,
    \quotient[12] , \quotient[13] , \quotient[14] , \quotient[15] ,
    \quotient[16] , \quotient[17] , \quotient[18] , \quotient[19] ,
    \quotient[20] , \quotient[21] , \quotient[22] , \quotient[23] ,
    \quotient[24] , \quotient[25] , \quotient[26] , \quotient[27] ,
    \quotient[28] , \quotient[29] , \quotient[30] , \quotient[31] ,
    \quotient[32] , \quotient[33] , \quotient[34] , \quotient[35] ,
    \quotient[36] , \quotient[37] , \quotient[38] , \quotient[39] ,
    \quotient[40] , \quotient[41] , \quotient[42] , \quotient[43] ,
    \quotient[44] , \quotient[45] , \quotient[46] , \quotient[47] ,
    \quotient[48] , \quotient[49] , \quotient[50] , \quotient[51] ,
    \quotient[52] , \quotient[53] , \quotient[54] , \quotient[55] ,
    \quotient[56] , \quotient[57] , \quotient[58] , \quotient[59] ,
    \quotient[60] , \quotient[61] , \quotient[62] , \quotient[63] ,
    \remainder[0] , \remainder[1] , \remainder[2] , \remainder[3] ,
    \remainder[4] , \remainder[5] , \remainder[6] , \remainder[7] ,
    \remainder[8] , \remainder[9] , \remainder[10] , \remainder[11] ,
    \remainder[12] , \remainder[13] , \remainder[14] , \remainder[15] ,
    \remainder[16] , \remainder[17] , \remainder[18] , \remainder[19] ,
    \remainder[20] , \remainder[21] , \remainder[22] , \remainder[23] ,
    \remainder[24] , \remainder[25] , \remainder[26] , \remainder[27] ,
    \remainder[28] , \remainder[29] , \remainder[30] , \remainder[31] ,
    \remainder[32] , \remainder[33] , \remainder[34] , \remainder[35] ,
    \remainder[36] , \remainder[37] , \remainder[38] , \remainder[39] ,
    \remainder[40] , \remainder[41] , \remainder[42] , \remainder[43] ,
    \remainder[44] , \remainder[45] , \remainder[46] , \remainder[47] ,
    \remainder[48] , \remainder[49] , \remainder[50] , \remainder[51] ,
    \remainder[52] , \remainder[53] , \remainder[54] , \remainder[55] ,
    \remainder[56] , \remainder[57] , \remainder[58] , \remainder[59] ,
    \remainder[60] , \remainder[61] , \remainder[62] , \remainder[63] ;
  wire new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_,
    new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_,
    new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_,
    new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_,
    new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_,
    new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_,
    new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_,
    new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_,
    new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_,
    new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_,
    new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_,
    new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_,
    new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_,
    new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_,
    new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_,
    new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_,
    new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_,
    new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_,
    new_n449_, new_n450_, new_n452_, new_n453_, new_n454_, new_n455_,
    new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_,
    new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_,
    new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_,
    new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_,
    new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_,
    new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_,
    new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_,
    new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_,
    new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_,
    new_n510_, new_n511_, new_n512_, new_n513_, new_n514_, new_n515_,
    new_n516_, new_n517_, new_n519_, new_n520_, new_n521_, new_n522_,
    new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_,
    new_n529_, new_n530_, new_n531_, new_n532_, new_n533_, new_n534_,
    new_n535_, new_n536_, new_n537_, new_n538_, new_n539_, new_n540_,
    new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_,
    new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_,
    new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_,
    new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_,
    new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_,
    new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_,
    new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_,
    new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_,
    new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_,
    new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_,
    new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_,
    new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1018_,
    new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_,
    new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_,
    new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_,
    new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_,
    new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_,
    new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_,
    new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_,
    new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_,
    new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_,
    new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_,
    new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_,
    new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_,
    new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_,
    new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_,
    new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_,
    new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_,
    new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_,
    new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_,
    new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_,
    new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_,
    new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_,
    new_n1145_, new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_,
    new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_,
    new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_,
    new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_,
    new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_,
    new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_,
    new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_,
    new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_,
    new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_,
    new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_,
    new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_,
    new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_,
    new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_,
    new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_,
    new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_,
    new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_,
    new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_,
    new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_,
    new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_,
    new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_,
    new_n1266_, new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_,
    new_n1272_, new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_,
    new_n1278_, new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_,
    new_n1284_, new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_,
    new_n1290_, new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1296_,
    new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_,
    new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1308_,
    new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_,
    new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1320_,
    new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_,
    new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_,
    new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_,
    new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_,
    new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_,
    new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_,
    new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_,
    new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_,
    new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_,
    new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_,
    new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_,
    new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_,
    new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_, new_n1398_,
    new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_,
    new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_,
    new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_,
    new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_,
    new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_,
    new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_,
    new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_,
    new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_, new_n1446_,
    new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_, new_n1452_,
    new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1458_, new_n1459_,
    new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1464_, new_n1465_,
    new_n1466_, new_n1467_, new_n1468_, new_n1469_, new_n1470_, new_n1471_,
    new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_, new_n1477_,
    new_n1478_, new_n1479_, new_n1480_, new_n1481_, new_n1482_, new_n1483_,
    new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_, new_n1489_,
    new_n1490_, new_n1491_, new_n1492_, new_n1493_, new_n1494_, new_n1495_,
    new_n1496_, new_n1497_, new_n1498_, new_n1499_, new_n1500_, new_n1501_,
    new_n1502_, new_n1503_, new_n1504_, new_n1505_, new_n1506_, new_n1507_,
    new_n1508_, new_n1509_, new_n1510_, new_n1511_, new_n1512_, new_n1513_,
    new_n1514_, new_n1515_, new_n1516_, new_n1517_, new_n1518_, new_n1519_,
    new_n1520_, new_n1521_, new_n1522_, new_n1523_, new_n1524_, new_n1525_,
    new_n1526_, new_n1527_, new_n1528_, new_n1529_, new_n1530_, new_n1531_,
    new_n1532_, new_n1533_, new_n1534_, new_n1535_, new_n1536_, new_n1537_,
    new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1542_, new_n1543_,
    new_n1544_, new_n1545_, new_n1546_, new_n1547_, new_n1548_, new_n1549_,
    new_n1550_, new_n1551_, new_n1552_, new_n1553_, new_n1554_, new_n1555_,
    new_n1556_, new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1561_,
    new_n1562_, new_n1563_, new_n1564_, new_n1565_, new_n1566_, new_n1567_,
    new_n1568_, new_n1569_, new_n1570_, new_n1571_, new_n1572_, new_n1573_,
    new_n1574_, new_n1575_, new_n1576_, new_n1577_, new_n1578_, new_n1579_,
    new_n1580_, new_n1581_, new_n1582_, new_n1583_, new_n1584_, new_n1585_,
    new_n1586_, new_n1587_, new_n1588_, new_n1589_, new_n1590_, new_n1591_,
    new_n1592_, new_n1593_, new_n1594_, new_n1595_, new_n1596_, new_n1597_,
    new_n1598_, new_n1599_, new_n1600_, new_n1601_, new_n1602_, new_n1603_,
    new_n1604_, new_n1605_, new_n1606_, new_n1607_, new_n1608_, new_n1609_,
    new_n1610_, new_n1611_, new_n1612_, new_n1613_, new_n1614_, new_n1615_,
    new_n1616_, new_n1617_, new_n1618_, new_n1619_, new_n1620_, new_n1621_,
    new_n1622_, new_n1623_, new_n1624_, new_n1625_, new_n1626_, new_n1628_,
    new_n1629_, new_n1630_, new_n1631_, new_n1632_, new_n1633_, new_n1634_,
    new_n1635_, new_n1636_, new_n1637_, new_n1638_, new_n1639_, new_n1640_,
    new_n1641_, new_n1642_, new_n1643_, new_n1644_, new_n1645_, new_n1646_,
    new_n1647_, new_n1648_, new_n1649_, new_n1650_, new_n1651_, new_n1652_,
    new_n1653_, new_n1654_, new_n1655_, new_n1656_, new_n1657_, new_n1658_,
    new_n1659_, new_n1660_, new_n1661_, new_n1662_, new_n1663_, new_n1664_,
    new_n1665_, new_n1666_, new_n1667_, new_n1668_, new_n1669_, new_n1670_,
    new_n1671_, new_n1672_, new_n1673_, new_n1674_, new_n1675_, new_n1676_,
    new_n1677_, new_n1678_, new_n1679_, new_n1680_, new_n1681_, new_n1682_,
    new_n1683_, new_n1684_, new_n1685_, new_n1686_, new_n1687_, new_n1688_,
    new_n1689_, new_n1690_, new_n1691_, new_n1692_, new_n1693_, new_n1694_,
    new_n1695_, new_n1696_, new_n1697_, new_n1698_, new_n1699_, new_n1700_,
    new_n1701_, new_n1702_, new_n1703_, new_n1704_, new_n1705_, new_n1706_,
    new_n1707_, new_n1708_, new_n1709_, new_n1710_, new_n1711_, new_n1712_,
    new_n1713_, new_n1714_, new_n1715_, new_n1716_, new_n1717_, new_n1718_,
    new_n1719_, new_n1720_, new_n1721_, new_n1722_, new_n1723_, new_n1724_,
    new_n1725_, new_n1726_, new_n1727_, new_n1728_, new_n1729_, new_n1730_,
    new_n1731_, new_n1732_, new_n1733_, new_n1734_, new_n1735_, new_n1736_,
    new_n1737_, new_n1738_, new_n1739_, new_n1740_, new_n1741_, new_n1742_,
    new_n1743_, new_n1744_, new_n1745_, new_n1746_, new_n1747_, new_n1748_,
    new_n1749_, new_n1750_, new_n1751_, new_n1752_, new_n1753_, new_n1754_,
    new_n1755_, new_n1756_, new_n1757_, new_n1758_, new_n1759_, new_n1760_,
    new_n1761_, new_n1762_, new_n1763_, new_n1764_, new_n1765_, new_n1766_,
    new_n1767_, new_n1768_, new_n1769_, new_n1770_, new_n1771_, new_n1772_,
    new_n1773_, new_n1774_, new_n1775_, new_n1776_, new_n1777_, new_n1778_,
    new_n1779_, new_n1780_, new_n1781_, new_n1782_, new_n1783_, new_n1784_,
    new_n1785_, new_n1786_, new_n1787_, new_n1788_, new_n1789_, new_n1790_,
    new_n1791_, new_n1792_, new_n1793_, new_n1794_, new_n1795_, new_n1796_,
    new_n1797_, new_n1798_, new_n1799_, new_n1800_, new_n1801_, new_n1802_,
    new_n1803_, new_n1804_, new_n1805_, new_n1806_, new_n1807_, new_n1808_,
    new_n1809_, new_n1810_, new_n1811_, new_n1812_, new_n1813_, new_n1814_,
    new_n1815_, new_n1816_, new_n1818_, new_n1819_, new_n1820_, new_n1821_,
    new_n1822_, new_n1823_, new_n1824_, new_n1825_, new_n1826_, new_n1827_,
    new_n1828_, new_n1829_, new_n1830_, new_n1831_, new_n1832_, new_n1833_,
    new_n1834_, new_n1835_, new_n1836_, new_n1837_, new_n1838_, new_n1839_,
    new_n1840_, new_n1841_, new_n1842_, new_n1843_, new_n1844_, new_n1845_,
    new_n1846_, new_n1847_, new_n1848_, new_n1849_, new_n1850_, new_n1851_,
    new_n1852_, new_n1853_, new_n1854_, new_n1855_, new_n1856_, new_n1857_,
    new_n1858_, new_n1859_, new_n1860_, new_n1861_, new_n1862_, new_n1863_,
    new_n1864_, new_n1865_, new_n1866_, new_n1867_, new_n1868_, new_n1869_,
    new_n1870_, new_n1871_, new_n1872_, new_n1873_, new_n1874_, new_n1875_,
    new_n1876_, new_n1877_, new_n1878_, new_n1879_, new_n1880_, new_n1881_,
    new_n1882_, new_n1883_, new_n1884_, new_n1885_, new_n1886_, new_n1887_,
    new_n1888_, new_n1889_, new_n1890_, new_n1891_, new_n1892_, new_n1893_,
    new_n1894_, new_n1895_, new_n1896_, new_n1897_, new_n1898_, new_n1899_,
    new_n1900_, new_n1901_, new_n1902_, new_n1903_, new_n1904_, new_n1905_,
    new_n1906_, new_n1907_, new_n1908_, new_n1909_, new_n1910_, new_n1911_,
    new_n1912_, new_n1913_, new_n1914_, new_n1915_, new_n1916_, new_n1917_,
    new_n1918_, new_n1919_, new_n1920_, new_n1921_, new_n1922_, new_n1923_,
    new_n1924_, new_n1925_, new_n1926_, new_n1927_, new_n1928_, new_n1929_,
    new_n1930_, new_n1931_, new_n1932_, new_n1933_, new_n1934_, new_n1935_,
    new_n1936_, new_n1937_, new_n1938_, new_n1939_, new_n1940_, new_n1941_,
    new_n1942_, new_n1943_, new_n1944_, new_n1945_, new_n1946_, new_n1947_,
    new_n1948_, new_n1949_, new_n1950_, new_n1951_, new_n1952_, new_n1953_,
    new_n1954_, new_n1955_, new_n1956_, new_n1957_, new_n1958_, new_n1959_,
    new_n1960_, new_n1961_, new_n1962_, new_n1963_, new_n1964_, new_n1965_,
    new_n1966_, new_n1967_, new_n1968_, new_n1969_, new_n1970_, new_n1971_,
    new_n1972_, new_n1973_, new_n1974_, new_n1975_, new_n1976_, new_n1977_,
    new_n1978_, new_n1979_, new_n1980_, new_n1981_, new_n1982_, new_n1983_,
    new_n1984_, new_n1985_, new_n1986_, new_n1987_, new_n1988_, new_n1989_,
    new_n1990_, new_n1991_, new_n1992_, new_n1993_, new_n1994_, new_n1995_,
    new_n1996_, new_n1997_, new_n1998_, new_n1999_, new_n2000_, new_n2001_,
    new_n2002_, new_n2003_, new_n2004_, new_n2005_, new_n2006_, new_n2007_,
    new_n2008_, new_n2009_, new_n2010_, new_n2011_, new_n2012_, new_n2013_,
    new_n2014_, new_n2015_, new_n2016_, new_n2017_, new_n2018_, new_n2019_,
    new_n2020_, new_n2021_, new_n2022_, new_n2024_, new_n2025_, new_n2026_,
    new_n2027_, new_n2028_, new_n2029_, new_n2030_, new_n2031_, new_n2032_,
    new_n2033_, new_n2034_, new_n2035_, new_n2036_, new_n2037_, new_n2038_,
    new_n2039_, new_n2040_, new_n2041_, new_n2042_, new_n2043_, new_n2044_,
    new_n2045_, new_n2046_, new_n2047_, new_n2048_, new_n2049_, new_n2050_,
    new_n2051_, new_n2052_, new_n2053_, new_n2054_, new_n2055_, new_n2056_,
    new_n2057_, new_n2058_, new_n2059_, new_n2060_, new_n2061_, new_n2062_,
    new_n2063_, new_n2064_, new_n2065_, new_n2066_, new_n2067_, new_n2068_,
    new_n2069_, new_n2070_, new_n2071_, new_n2072_, new_n2073_, new_n2074_,
    new_n2075_, new_n2076_, new_n2077_, new_n2078_, new_n2079_, new_n2080_,
    new_n2081_, new_n2082_, new_n2083_, new_n2084_, new_n2085_, new_n2086_,
    new_n2087_, new_n2088_, new_n2089_, new_n2090_, new_n2091_, new_n2092_,
    new_n2093_, new_n2094_, new_n2095_, new_n2096_, new_n2097_, new_n2098_,
    new_n2099_, new_n2100_, new_n2101_, new_n2102_, new_n2103_, new_n2104_,
    new_n2105_, new_n2106_, new_n2107_, new_n2108_, new_n2109_, new_n2110_,
    new_n2111_, new_n2112_, new_n2113_, new_n2114_, new_n2115_, new_n2116_,
    new_n2117_, new_n2118_, new_n2119_, new_n2120_, new_n2121_, new_n2122_,
    new_n2123_, new_n2124_, new_n2125_, new_n2126_, new_n2127_, new_n2128_,
    new_n2129_, new_n2130_, new_n2131_, new_n2132_, new_n2133_, new_n2134_,
    new_n2135_, new_n2136_, new_n2137_, new_n2138_, new_n2139_, new_n2140_,
    new_n2141_, new_n2142_, new_n2143_, new_n2144_, new_n2145_, new_n2146_,
    new_n2147_, new_n2148_, new_n2149_, new_n2150_, new_n2151_, new_n2152_,
    new_n2153_, new_n2154_, new_n2155_, new_n2156_, new_n2157_, new_n2158_,
    new_n2159_, new_n2160_, new_n2161_, new_n2162_, new_n2163_, new_n2164_,
    new_n2165_, new_n2166_, new_n2167_, new_n2168_, new_n2169_, new_n2170_,
    new_n2171_, new_n2172_, new_n2173_, new_n2174_, new_n2175_, new_n2176_,
    new_n2177_, new_n2178_, new_n2179_, new_n2180_, new_n2181_, new_n2182_,
    new_n2183_, new_n2184_, new_n2185_, new_n2186_, new_n2187_, new_n2188_,
    new_n2189_, new_n2190_, new_n2191_, new_n2192_, new_n2193_, new_n2194_,
    new_n2195_, new_n2196_, new_n2197_, new_n2198_, new_n2199_, new_n2200_,
    new_n2201_, new_n2202_, new_n2203_, new_n2204_, new_n2205_, new_n2206_,
    new_n2207_, new_n2208_, new_n2209_, new_n2210_, new_n2211_, new_n2212_,
    new_n2213_, new_n2214_, new_n2215_, new_n2216_, new_n2217_, new_n2218_,
    new_n2219_, new_n2220_, new_n2221_, new_n2222_, new_n2223_, new_n2224_,
    new_n2225_, new_n2226_, new_n2227_, new_n2228_, new_n2229_, new_n2230_,
    new_n2231_, new_n2232_, new_n2234_, new_n2235_, new_n2236_, new_n2237_,
    new_n2238_, new_n2239_, new_n2240_, new_n2241_, new_n2242_, new_n2243_,
    new_n2244_, new_n2245_, new_n2246_, new_n2247_, new_n2248_, new_n2249_,
    new_n2250_, new_n2251_, new_n2252_, new_n2253_, new_n2254_, new_n2255_,
    new_n2256_, new_n2257_, new_n2258_, new_n2259_, new_n2260_, new_n2261_,
    new_n2262_, new_n2263_, new_n2264_, new_n2265_, new_n2266_, new_n2267_,
    new_n2268_, new_n2269_, new_n2270_, new_n2271_, new_n2272_, new_n2273_,
    new_n2274_, new_n2275_, new_n2276_, new_n2277_, new_n2278_, new_n2279_,
    new_n2280_, new_n2281_, new_n2282_, new_n2283_, new_n2284_, new_n2285_,
    new_n2286_, new_n2287_, new_n2288_, new_n2289_, new_n2290_, new_n2291_,
    new_n2292_, new_n2293_, new_n2294_, new_n2295_, new_n2296_, new_n2297_,
    new_n2298_, new_n2299_, new_n2300_, new_n2301_, new_n2302_, new_n2303_,
    new_n2304_, new_n2305_, new_n2306_, new_n2307_, new_n2308_, new_n2309_,
    new_n2310_, new_n2311_, new_n2312_, new_n2313_, new_n2314_, new_n2315_,
    new_n2316_, new_n2317_, new_n2318_, new_n2319_, new_n2320_, new_n2321_,
    new_n2322_, new_n2323_, new_n2324_, new_n2325_, new_n2326_, new_n2327_,
    new_n2328_, new_n2329_, new_n2330_, new_n2331_, new_n2332_, new_n2333_,
    new_n2334_, new_n2335_, new_n2336_, new_n2337_, new_n2338_, new_n2339_,
    new_n2340_, new_n2341_, new_n2342_, new_n2343_, new_n2344_, new_n2345_,
    new_n2346_, new_n2347_, new_n2348_, new_n2349_, new_n2350_, new_n2351_,
    new_n2352_, new_n2353_, new_n2354_, new_n2355_, new_n2356_, new_n2357_,
    new_n2358_, new_n2359_, new_n2360_, new_n2361_, new_n2362_, new_n2363_,
    new_n2364_, new_n2365_, new_n2366_, new_n2367_, new_n2368_, new_n2369_,
    new_n2370_, new_n2371_, new_n2372_, new_n2373_, new_n2374_, new_n2375_,
    new_n2376_, new_n2377_, new_n2378_, new_n2379_, new_n2380_, new_n2381_,
    new_n2382_, new_n2383_, new_n2384_, new_n2385_, new_n2386_, new_n2387_,
    new_n2388_, new_n2389_, new_n2390_, new_n2391_, new_n2392_, new_n2393_,
    new_n2394_, new_n2395_, new_n2396_, new_n2397_, new_n2398_, new_n2399_,
    new_n2400_, new_n2401_, new_n2402_, new_n2403_, new_n2404_, new_n2405_,
    new_n2406_, new_n2407_, new_n2408_, new_n2409_, new_n2410_, new_n2411_,
    new_n2412_, new_n2413_, new_n2414_, new_n2415_, new_n2416_, new_n2417_,
    new_n2418_, new_n2419_, new_n2420_, new_n2421_, new_n2422_, new_n2423_,
    new_n2424_, new_n2425_, new_n2426_, new_n2427_, new_n2428_, new_n2429_,
    new_n2430_, new_n2431_, new_n2432_, new_n2433_, new_n2434_, new_n2435_,
    new_n2436_, new_n2437_, new_n2438_, new_n2439_, new_n2440_, new_n2441_,
    new_n2442_, new_n2443_, new_n2444_, new_n2445_, new_n2446_, new_n2447_,
    new_n2448_, new_n2449_, new_n2450_, new_n2451_, new_n2452_, new_n2453_,
    new_n2454_, new_n2455_, new_n2456_, new_n2457_, new_n2458_, new_n2459_,
    new_n2460_, new_n2462_, new_n2463_, new_n2464_, new_n2465_, new_n2466_,
    new_n2467_, new_n2468_, new_n2469_, new_n2470_, new_n2471_, new_n2472_,
    new_n2473_, new_n2474_, new_n2475_, new_n2476_, new_n2477_, new_n2478_,
    new_n2479_, new_n2480_, new_n2481_, new_n2482_, new_n2483_, new_n2484_,
    new_n2485_, new_n2486_, new_n2487_, new_n2488_, new_n2489_, new_n2490_,
    new_n2491_, new_n2492_, new_n2493_, new_n2494_, new_n2495_, new_n2496_,
    new_n2497_, new_n2498_, new_n2499_, new_n2500_, new_n2501_, new_n2502_,
    new_n2503_, new_n2504_, new_n2505_, new_n2506_, new_n2507_, new_n2508_,
    new_n2509_, new_n2510_, new_n2511_, new_n2512_, new_n2513_, new_n2514_,
    new_n2515_, new_n2516_, new_n2517_, new_n2518_, new_n2519_, new_n2520_,
    new_n2521_, new_n2522_, new_n2523_, new_n2524_, new_n2525_, new_n2526_,
    new_n2527_, new_n2528_, new_n2529_, new_n2530_, new_n2531_, new_n2532_,
    new_n2533_, new_n2534_, new_n2535_, new_n2536_, new_n2537_, new_n2538_,
    new_n2539_, new_n2540_, new_n2541_, new_n2542_, new_n2543_, new_n2544_,
    new_n2545_, new_n2546_, new_n2547_, new_n2548_, new_n2549_, new_n2550_,
    new_n2551_, new_n2552_, new_n2553_, new_n2554_, new_n2555_, new_n2556_,
    new_n2557_, new_n2558_, new_n2559_, new_n2560_, new_n2561_, new_n2562_,
    new_n2563_, new_n2564_, new_n2565_, new_n2566_, new_n2567_, new_n2568_,
    new_n2569_, new_n2570_, new_n2571_, new_n2572_, new_n2573_, new_n2574_,
    new_n2575_, new_n2576_, new_n2577_, new_n2578_, new_n2579_, new_n2580_,
    new_n2581_, new_n2582_, new_n2583_, new_n2584_, new_n2585_, new_n2586_,
    new_n2587_, new_n2588_, new_n2589_, new_n2590_, new_n2591_, new_n2592_,
    new_n2593_, new_n2594_, new_n2595_, new_n2596_, new_n2597_, new_n2598_,
    new_n2599_, new_n2600_, new_n2601_, new_n2602_, new_n2603_, new_n2604_,
    new_n2605_, new_n2606_, new_n2607_, new_n2608_, new_n2609_, new_n2610_,
    new_n2611_, new_n2612_, new_n2613_, new_n2614_, new_n2615_, new_n2616_,
    new_n2617_, new_n2618_, new_n2619_, new_n2620_, new_n2621_, new_n2622_,
    new_n2623_, new_n2624_, new_n2625_, new_n2626_, new_n2627_, new_n2628_,
    new_n2629_, new_n2630_, new_n2631_, new_n2632_, new_n2633_, new_n2634_,
    new_n2635_, new_n2636_, new_n2637_, new_n2638_, new_n2639_, new_n2640_,
    new_n2641_, new_n2642_, new_n2643_, new_n2644_, new_n2645_, new_n2646_,
    new_n2647_, new_n2648_, new_n2649_, new_n2650_, new_n2651_, new_n2652_,
    new_n2653_, new_n2654_, new_n2655_, new_n2656_, new_n2657_, new_n2658_,
    new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2663_, new_n2664_,
    new_n2665_, new_n2666_, new_n2667_, new_n2668_, new_n2669_, new_n2670_,
    new_n2671_, new_n2672_, new_n2673_, new_n2674_, new_n2675_, new_n2676_,
    new_n2677_, new_n2678_, new_n2679_, new_n2680_, new_n2681_, new_n2682_,
    new_n2683_, new_n2684_, new_n2685_, new_n2686_, new_n2687_, new_n2688_,
    new_n2689_, new_n2690_, new_n2691_, new_n2692_, new_n2693_, new_n2694_,
    new_n2695_, new_n2696_, new_n2697_, new_n2698_, new_n2699_, new_n2700_,
    new_n2701_, new_n2702_, new_n2703_, new_n2704_, new_n2705_, new_n2706_,
    new_n2707_, new_n2708_, new_n2709_, new_n2711_, new_n2712_, new_n2713_,
    new_n2714_, new_n2715_, new_n2716_, new_n2717_, new_n2718_, new_n2719_,
    new_n2720_, new_n2721_, new_n2722_, new_n2723_, new_n2724_, new_n2725_,
    new_n2726_, new_n2727_, new_n2728_, new_n2729_, new_n2730_, new_n2731_,
    new_n2732_, new_n2733_, new_n2734_, new_n2735_, new_n2736_, new_n2737_,
    new_n2738_, new_n2739_, new_n2740_, new_n2741_, new_n2742_, new_n2743_,
    new_n2744_, new_n2745_, new_n2746_, new_n2747_, new_n2748_, new_n2749_,
    new_n2750_, new_n2751_, new_n2752_, new_n2753_, new_n2754_, new_n2755_,
    new_n2756_, new_n2757_, new_n2758_, new_n2759_, new_n2760_, new_n2761_,
    new_n2762_, new_n2763_, new_n2764_, new_n2765_, new_n2766_, new_n2767_,
    new_n2768_, new_n2769_, new_n2770_, new_n2771_, new_n2772_, new_n2773_,
    new_n2774_, new_n2775_, new_n2776_, new_n2777_, new_n2778_, new_n2779_,
    new_n2780_, new_n2781_, new_n2782_, new_n2783_, new_n2784_, new_n2785_,
    new_n2786_, new_n2787_, new_n2788_, new_n2789_, new_n2790_, new_n2791_,
    new_n2792_, new_n2793_, new_n2794_, new_n2795_, new_n2796_, new_n2797_,
    new_n2798_, new_n2799_, new_n2800_, new_n2801_, new_n2802_, new_n2803_,
    new_n2804_, new_n2805_, new_n2806_, new_n2807_, new_n2808_, new_n2809_,
    new_n2810_, new_n2811_, new_n2812_, new_n2813_, new_n2814_, new_n2815_,
    new_n2816_, new_n2817_, new_n2818_, new_n2819_, new_n2820_, new_n2821_,
    new_n2822_, new_n2823_, new_n2824_, new_n2825_, new_n2826_, new_n2827_,
    new_n2828_, new_n2829_, new_n2830_, new_n2831_, new_n2832_, new_n2833_,
    new_n2834_, new_n2835_, new_n2836_, new_n2837_, new_n2838_, new_n2839_,
    new_n2840_, new_n2841_, new_n2842_, new_n2843_, new_n2844_, new_n2845_,
    new_n2846_, new_n2847_, new_n2848_, new_n2849_, new_n2850_, new_n2851_,
    new_n2852_, new_n2853_, new_n2854_, new_n2855_, new_n2856_, new_n2857_,
    new_n2858_, new_n2859_, new_n2860_, new_n2861_, new_n2862_, new_n2863_,
    new_n2864_, new_n2865_, new_n2866_, new_n2867_, new_n2868_, new_n2869_,
    new_n2870_, new_n2871_, new_n2872_, new_n2873_, new_n2874_, new_n2875_,
    new_n2876_, new_n2877_, new_n2878_, new_n2879_, new_n2880_, new_n2881_,
    new_n2882_, new_n2883_, new_n2884_, new_n2885_, new_n2886_, new_n2887_,
    new_n2888_, new_n2889_, new_n2890_, new_n2891_, new_n2892_, new_n2893_,
    new_n2894_, new_n2895_, new_n2896_, new_n2897_, new_n2898_, new_n2899_,
    new_n2900_, new_n2901_, new_n2902_, new_n2903_, new_n2904_, new_n2905_,
    new_n2906_, new_n2907_, new_n2908_, new_n2909_, new_n2910_, new_n2911_,
    new_n2912_, new_n2913_, new_n2914_, new_n2915_, new_n2916_, new_n2917_,
    new_n2918_, new_n2919_, new_n2920_, new_n2921_, new_n2922_, new_n2923_,
    new_n2924_, new_n2925_, new_n2926_, new_n2927_, new_n2928_, new_n2929_,
    new_n2930_, new_n2931_, new_n2932_, new_n2933_, new_n2934_, new_n2935_,
    new_n2936_, new_n2937_, new_n2938_, new_n2939_, new_n2940_, new_n2941_,
    new_n2942_, new_n2943_, new_n2944_, new_n2945_, new_n2946_, new_n2947_,
    new_n2948_, new_n2949_, new_n2950_, new_n2951_, new_n2952_, new_n2953_,
    new_n2954_, new_n2955_, new_n2956_, new_n2957_, new_n2958_, new_n2959_,
    new_n2960_, new_n2961_, new_n2962_, new_n2963_, new_n2964_, new_n2965_,
    new_n2967_, new_n2968_, new_n2969_, new_n2970_, new_n2971_, new_n2972_,
    new_n2973_, new_n2974_, new_n2975_, new_n2976_, new_n2977_, new_n2978_,
    new_n2979_, new_n2980_, new_n2981_, new_n2982_, new_n2983_, new_n2984_,
    new_n2985_, new_n2986_, new_n2987_, new_n2988_, new_n2989_, new_n2990_,
    new_n2991_, new_n2992_, new_n2993_, new_n2994_, new_n2995_, new_n2996_,
    new_n2997_, new_n2998_, new_n2999_, new_n3000_, new_n3001_, new_n3002_,
    new_n3003_, new_n3004_, new_n3005_, new_n3006_, new_n3007_, new_n3008_,
    new_n3009_, new_n3010_, new_n3011_, new_n3012_, new_n3013_, new_n3014_,
    new_n3015_, new_n3016_, new_n3017_, new_n3018_, new_n3019_, new_n3020_,
    new_n3021_, new_n3022_, new_n3023_, new_n3024_, new_n3025_, new_n3026_,
    new_n3027_, new_n3028_, new_n3029_, new_n3030_, new_n3031_, new_n3032_,
    new_n3033_, new_n3034_, new_n3035_, new_n3036_, new_n3037_, new_n3038_,
    new_n3039_, new_n3040_, new_n3041_, new_n3042_, new_n3043_, new_n3044_,
    new_n3045_, new_n3046_, new_n3047_, new_n3048_, new_n3049_, new_n3050_,
    new_n3051_, new_n3052_, new_n3053_, new_n3054_, new_n3055_, new_n3056_,
    new_n3057_, new_n3058_, new_n3059_, new_n3060_, new_n3061_, new_n3062_,
    new_n3063_, new_n3064_, new_n3065_, new_n3066_, new_n3067_, new_n3068_,
    new_n3069_, new_n3070_, new_n3071_, new_n3072_, new_n3073_, new_n3074_,
    new_n3075_, new_n3076_, new_n3077_, new_n3078_, new_n3079_, new_n3080_,
    new_n3081_, new_n3082_, new_n3083_, new_n3084_, new_n3085_, new_n3086_,
    new_n3087_, new_n3088_, new_n3089_, new_n3090_, new_n3091_, new_n3092_,
    new_n3093_, new_n3094_, new_n3095_, new_n3096_, new_n3097_, new_n3098_,
    new_n3099_, new_n3100_, new_n3101_, new_n3102_, new_n3103_, new_n3104_,
    new_n3105_, new_n3106_, new_n3107_, new_n3108_, new_n3109_, new_n3110_,
    new_n3111_, new_n3112_, new_n3113_, new_n3114_, new_n3115_, new_n3116_,
    new_n3117_, new_n3118_, new_n3119_, new_n3120_, new_n3121_, new_n3122_,
    new_n3123_, new_n3124_, new_n3125_, new_n3126_, new_n3127_, new_n3128_,
    new_n3129_, new_n3130_, new_n3131_, new_n3132_, new_n3133_, new_n3134_,
    new_n3135_, new_n3136_, new_n3137_, new_n3138_, new_n3139_, new_n3140_,
    new_n3141_, new_n3142_, new_n3143_, new_n3144_, new_n3145_, new_n3146_,
    new_n3147_, new_n3148_, new_n3149_, new_n3150_, new_n3151_, new_n3152_,
    new_n3153_, new_n3154_, new_n3155_, new_n3156_, new_n3157_, new_n3158_,
    new_n3159_, new_n3160_, new_n3161_, new_n3162_, new_n3163_, new_n3164_,
    new_n3165_, new_n3166_, new_n3167_, new_n3168_, new_n3169_, new_n3170_,
    new_n3171_, new_n3172_, new_n3173_, new_n3174_, new_n3175_, new_n3176_,
    new_n3177_, new_n3178_, new_n3179_, new_n3180_, new_n3181_, new_n3182_,
    new_n3183_, new_n3184_, new_n3185_, new_n3186_, new_n3187_, new_n3188_,
    new_n3189_, new_n3190_, new_n3191_, new_n3192_, new_n3193_, new_n3194_,
    new_n3195_, new_n3196_, new_n3197_, new_n3198_, new_n3199_, new_n3200_,
    new_n3201_, new_n3202_, new_n3203_, new_n3204_, new_n3205_, new_n3206_,
    new_n3207_, new_n3208_, new_n3209_, new_n3210_, new_n3211_, new_n3212_,
    new_n3213_, new_n3214_, new_n3215_, new_n3216_, new_n3217_, new_n3218_,
    new_n3219_, new_n3220_, new_n3221_, new_n3222_, new_n3223_, new_n3224_,
    new_n3225_, new_n3226_, new_n3227_, new_n3228_, new_n3229_, new_n3230_,
    new_n3231_, new_n3232_, new_n3233_, new_n3234_, new_n3235_, new_n3236_,
    new_n3237_, new_n3238_, new_n3240_, new_n3241_, new_n3242_, new_n3243_,
    new_n3244_, new_n3245_, new_n3246_, new_n3247_, new_n3248_, new_n3249_,
    new_n3250_, new_n3251_, new_n3252_, new_n3253_, new_n3254_, new_n3255_,
    new_n3256_, new_n3257_, new_n3258_, new_n3259_, new_n3260_, new_n3261_,
    new_n3262_, new_n3263_, new_n3264_, new_n3265_, new_n3266_, new_n3267_,
    new_n3268_, new_n3269_, new_n3270_, new_n3271_, new_n3272_, new_n3273_,
    new_n3274_, new_n3275_, new_n3276_, new_n3277_, new_n3278_, new_n3279_,
    new_n3280_, new_n3281_, new_n3282_, new_n3283_, new_n3284_, new_n3285_,
    new_n3286_, new_n3287_, new_n3288_, new_n3289_, new_n3290_, new_n3291_,
    new_n3292_, new_n3293_, new_n3294_, new_n3295_, new_n3296_, new_n3297_,
    new_n3298_, new_n3299_, new_n3300_, new_n3301_, new_n3302_, new_n3303_,
    new_n3304_, new_n3305_, new_n3306_, new_n3307_, new_n3308_, new_n3309_,
    new_n3310_, new_n3311_, new_n3312_, new_n3313_, new_n3314_, new_n3315_,
    new_n3316_, new_n3317_, new_n3318_, new_n3319_, new_n3320_, new_n3321_,
    new_n3322_, new_n3323_, new_n3324_, new_n3325_, new_n3326_, new_n3327_,
    new_n3328_, new_n3329_, new_n3330_, new_n3331_, new_n3332_, new_n3333_,
    new_n3334_, new_n3335_, new_n3336_, new_n3337_, new_n3338_, new_n3339_,
    new_n3340_, new_n3341_, new_n3342_, new_n3343_, new_n3344_, new_n3345_,
    new_n3346_, new_n3347_, new_n3348_, new_n3349_, new_n3350_, new_n3351_,
    new_n3352_, new_n3353_, new_n3354_, new_n3355_, new_n3356_, new_n3357_,
    new_n3358_, new_n3359_, new_n3360_, new_n3361_, new_n3362_, new_n3363_,
    new_n3364_, new_n3365_, new_n3366_, new_n3367_, new_n3368_, new_n3369_,
    new_n3370_, new_n3371_, new_n3372_, new_n3373_, new_n3374_, new_n3375_,
    new_n3376_, new_n3377_, new_n3378_, new_n3379_, new_n3380_, new_n3381_,
    new_n3382_, new_n3383_, new_n3384_, new_n3385_, new_n3386_, new_n3387_,
    new_n3388_, new_n3389_, new_n3390_, new_n3391_, new_n3392_, new_n3393_,
    new_n3394_, new_n3395_, new_n3396_, new_n3397_, new_n3398_, new_n3399_,
    new_n3400_, new_n3401_, new_n3402_, new_n3403_, new_n3404_, new_n3405_,
    new_n3406_, new_n3407_, new_n3408_, new_n3409_, new_n3410_, new_n3411_,
    new_n3412_, new_n3413_, new_n3414_, new_n3415_, new_n3416_, new_n3417_,
    new_n3418_, new_n3419_, new_n3420_, new_n3421_, new_n3422_, new_n3423_,
    new_n3424_, new_n3425_, new_n3426_, new_n3427_, new_n3428_, new_n3429_,
    new_n3430_, new_n3431_, new_n3432_, new_n3433_, new_n3434_, new_n3435_,
    new_n3436_, new_n3437_, new_n3438_, new_n3439_, new_n3440_, new_n3441_,
    new_n3442_, new_n3443_, new_n3444_, new_n3445_, new_n3446_, new_n3447_,
    new_n3448_, new_n3449_, new_n3450_, new_n3451_, new_n3452_, new_n3453_,
    new_n3454_, new_n3455_, new_n3456_, new_n3457_, new_n3458_, new_n3459_,
    new_n3460_, new_n3461_, new_n3462_, new_n3463_, new_n3464_, new_n3465_,
    new_n3466_, new_n3467_, new_n3468_, new_n3469_, new_n3470_, new_n3471_,
    new_n3472_, new_n3473_, new_n3474_, new_n3475_, new_n3476_, new_n3477_,
    new_n3478_, new_n3479_, new_n3480_, new_n3481_, new_n3482_, new_n3483_,
    new_n3484_, new_n3485_, new_n3486_, new_n3487_, new_n3488_, new_n3489_,
    new_n3490_, new_n3491_, new_n3492_, new_n3493_, new_n3494_, new_n3495_,
    new_n3496_, new_n3497_, new_n3498_, new_n3499_, new_n3500_, new_n3501_,
    new_n3502_, new_n3503_, new_n3504_, new_n3505_, new_n3506_, new_n3507_,
    new_n3508_, new_n3509_, new_n3510_, new_n3511_, new_n3512_, new_n3513_,
    new_n3514_, new_n3515_, new_n3516_, new_n3517_, new_n3518_, new_n3519_,
    new_n3520_, new_n3521_, new_n3522_, new_n3523_, new_n3524_, new_n3525_,
    new_n3527_, new_n3528_, new_n3529_, new_n3530_, new_n3531_, new_n3532_,
    new_n3533_, new_n3534_, new_n3535_, new_n3536_, new_n3537_, new_n3538_,
    new_n3539_, new_n3540_, new_n3541_, new_n3542_, new_n3543_, new_n3544_,
    new_n3545_, new_n3546_, new_n3547_, new_n3548_, new_n3549_, new_n3550_,
    new_n3551_, new_n3552_, new_n3553_, new_n3554_, new_n3555_, new_n3556_,
    new_n3557_, new_n3558_, new_n3559_, new_n3560_, new_n3561_, new_n3562_,
    new_n3563_, new_n3564_, new_n3565_, new_n3566_, new_n3567_, new_n3568_,
    new_n3569_, new_n3570_, new_n3571_, new_n3572_, new_n3573_, new_n3574_,
    new_n3575_, new_n3576_, new_n3577_, new_n3578_, new_n3579_, new_n3580_,
    new_n3581_, new_n3582_, new_n3583_, new_n3584_, new_n3585_, new_n3586_,
    new_n3587_, new_n3588_, new_n3589_, new_n3590_, new_n3591_, new_n3592_,
    new_n3593_, new_n3594_, new_n3595_, new_n3596_, new_n3597_, new_n3598_,
    new_n3599_, new_n3600_, new_n3601_, new_n3602_, new_n3603_, new_n3604_,
    new_n3605_, new_n3606_, new_n3607_, new_n3608_, new_n3609_, new_n3610_,
    new_n3611_, new_n3612_, new_n3613_, new_n3614_, new_n3615_, new_n3616_,
    new_n3617_, new_n3618_, new_n3619_, new_n3620_, new_n3621_, new_n3622_,
    new_n3623_, new_n3624_, new_n3625_, new_n3626_, new_n3627_, new_n3628_,
    new_n3629_, new_n3630_, new_n3631_, new_n3632_, new_n3633_, new_n3634_,
    new_n3635_, new_n3636_, new_n3637_, new_n3638_, new_n3639_, new_n3640_,
    new_n3641_, new_n3642_, new_n3643_, new_n3644_, new_n3645_, new_n3646_,
    new_n3647_, new_n3648_, new_n3649_, new_n3650_, new_n3651_, new_n3652_,
    new_n3653_, new_n3654_, new_n3655_, new_n3656_, new_n3657_, new_n3658_,
    new_n3659_, new_n3660_, new_n3661_, new_n3662_, new_n3663_, new_n3664_,
    new_n3665_, new_n3666_, new_n3667_, new_n3668_, new_n3669_, new_n3670_,
    new_n3671_, new_n3672_, new_n3673_, new_n3674_, new_n3675_, new_n3676_,
    new_n3677_, new_n3678_, new_n3679_, new_n3680_, new_n3681_, new_n3682_,
    new_n3683_, new_n3684_, new_n3685_, new_n3686_, new_n3687_, new_n3688_,
    new_n3689_, new_n3690_, new_n3691_, new_n3692_, new_n3693_, new_n3694_,
    new_n3695_, new_n3696_, new_n3697_, new_n3698_, new_n3699_, new_n3700_,
    new_n3701_, new_n3702_, new_n3703_, new_n3704_, new_n3705_, new_n3706_,
    new_n3707_, new_n3708_, new_n3709_, new_n3710_, new_n3711_, new_n3712_,
    new_n3713_, new_n3714_, new_n3715_, new_n3716_, new_n3717_, new_n3718_,
    new_n3719_, new_n3720_, new_n3721_, new_n3722_, new_n3723_, new_n3724_,
    new_n3725_, new_n3726_, new_n3727_, new_n3728_, new_n3729_, new_n3730_,
    new_n3731_, new_n3732_, new_n3733_, new_n3734_, new_n3735_, new_n3736_,
    new_n3737_, new_n3738_, new_n3739_, new_n3740_, new_n3741_, new_n3742_,
    new_n3743_, new_n3744_, new_n3745_, new_n3746_, new_n3747_, new_n3748_,
    new_n3749_, new_n3750_, new_n3751_, new_n3752_, new_n3753_, new_n3754_,
    new_n3755_, new_n3756_, new_n3757_, new_n3758_, new_n3759_, new_n3760_,
    new_n3761_, new_n3762_, new_n3763_, new_n3764_, new_n3765_, new_n3766_,
    new_n3767_, new_n3768_, new_n3769_, new_n3770_, new_n3771_, new_n3772_,
    new_n3773_, new_n3774_, new_n3775_, new_n3776_, new_n3777_, new_n3778_,
    new_n3779_, new_n3780_, new_n3781_, new_n3782_, new_n3783_, new_n3784_,
    new_n3785_, new_n3786_, new_n3787_, new_n3788_, new_n3789_, new_n3790_,
    new_n3791_, new_n3792_, new_n3793_, new_n3794_, new_n3795_, new_n3796_,
    new_n3797_, new_n3798_, new_n3799_, new_n3800_, new_n3801_, new_n3802_,
    new_n3803_, new_n3804_, new_n3805_, new_n3806_, new_n3807_, new_n3808_,
    new_n3809_, new_n3810_, new_n3811_, new_n3812_, new_n3813_, new_n3814_,
    new_n3815_, new_n3816_, new_n3817_, new_n3818_, new_n3819_, new_n3820_,
    new_n3821_, new_n3822_, new_n3823_, new_n3825_, new_n3826_, new_n3827_,
    new_n3828_, new_n3829_, new_n3830_, new_n3831_, new_n3832_, new_n3833_,
    new_n3834_, new_n3835_, new_n3836_, new_n3837_, new_n3838_, new_n3839_,
    new_n3840_, new_n3841_, new_n3842_, new_n3843_, new_n3844_, new_n3845_,
    new_n3846_, new_n3847_, new_n3848_, new_n3849_, new_n3850_, new_n3851_,
    new_n3852_, new_n3853_, new_n3854_, new_n3855_, new_n3856_, new_n3857_,
    new_n3858_, new_n3859_, new_n3860_, new_n3861_, new_n3862_, new_n3863_,
    new_n3864_, new_n3865_, new_n3866_, new_n3867_, new_n3868_, new_n3869_,
    new_n3870_, new_n3871_, new_n3872_, new_n3873_, new_n3874_, new_n3875_,
    new_n3876_, new_n3877_, new_n3878_, new_n3879_, new_n3880_, new_n3881_,
    new_n3882_, new_n3883_, new_n3884_, new_n3885_, new_n3886_, new_n3887_,
    new_n3888_, new_n3889_, new_n3890_, new_n3891_, new_n3892_, new_n3893_,
    new_n3894_, new_n3895_, new_n3896_, new_n3897_, new_n3898_, new_n3899_,
    new_n3900_, new_n3901_, new_n3902_, new_n3903_, new_n3904_, new_n3905_,
    new_n3906_, new_n3907_, new_n3908_, new_n3909_, new_n3910_, new_n3911_,
    new_n3912_, new_n3913_, new_n3914_, new_n3915_, new_n3916_, new_n3917_,
    new_n3918_, new_n3919_, new_n3920_, new_n3921_, new_n3922_, new_n3923_,
    new_n3924_, new_n3925_, new_n3926_, new_n3927_, new_n3928_, new_n3929_,
    new_n3930_, new_n3931_, new_n3932_, new_n3933_, new_n3934_, new_n3935_,
    new_n3936_, new_n3937_, new_n3938_, new_n3939_, new_n3940_, new_n3941_,
    new_n3942_, new_n3943_, new_n3944_, new_n3945_, new_n3946_, new_n3947_,
    new_n3948_, new_n3949_, new_n3950_, new_n3951_, new_n3952_, new_n3953_,
    new_n3954_, new_n3955_, new_n3956_, new_n3957_, new_n3958_, new_n3959_,
    new_n3960_, new_n3961_, new_n3962_, new_n3963_, new_n3964_, new_n3965_,
    new_n3966_, new_n3967_, new_n3968_, new_n3969_, new_n3970_, new_n3971_,
    new_n3972_, new_n3973_, new_n3974_, new_n3975_, new_n3976_, new_n3977_,
    new_n3978_, new_n3979_, new_n3980_, new_n3981_, new_n3982_, new_n3983_,
    new_n3984_, new_n3985_, new_n3986_, new_n3987_, new_n3988_, new_n3989_,
    new_n3990_, new_n3991_, new_n3992_, new_n3993_, new_n3994_, new_n3995_,
    new_n3996_, new_n3997_, new_n3998_, new_n3999_, new_n4000_, new_n4001_,
    new_n4002_, new_n4003_, new_n4004_, new_n4005_, new_n4006_, new_n4007_,
    new_n4008_, new_n4009_, new_n4010_, new_n4011_, new_n4012_, new_n4013_,
    new_n4014_, new_n4015_, new_n4016_, new_n4017_, new_n4018_, new_n4019_,
    new_n4020_, new_n4021_, new_n4022_, new_n4023_, new_n4024_, new_n4025_,
    new_n4026_, new_n4027_, new_n4028_, new_n4029_, new_n4030_, new_n4031_,
    new_n4032_, new_n4033_, new_n4034_, new_n4035_, new_n4036_, new_n4037_,
    new_n4038_, new_n4039_, new_n4040_, new_n4041_, new_n4042_, new_n4043_,
    new_n4044_, new_n4045_, new_n4046_, new_n4047_, new_n4048_, new_n4049_,
    new_n4050_, new_n4051_, new_n4052_, new_n4053_, new_n4054_, new_n4055_,
    new_n4056_, new_n4057_, new_n4058_, new_n4059_, new_n4060_, new_n4061_,
    new_n4062_, new_n4063_, new_n4064_, new_n4065_, new_n4066_, new_n4067_,
    new_n4068_, new_n4069_, new_n4070_, new_n4071_, new_n4072_, new_n4073_,
    new_n4074_, new_n4075_, new_n4076_, new_n4077_, new_n4078_, new_n4079_,
    new_n4080_, new_n4081_, new_n4082_, new_n4083_, new_n4084_, new_n4085_,
    new_n4086_, new_n4087_, new_n4088_, new_n4089_, new_n4090_, new_n4091_,
    new_n4092_, new_n4093_, new_n4094_, new_n4095_, new_n4096_, new_n4097_,
    new_n4098_, new_n4099_, new_n4100_, new_n4101_, new_n4102_, new_n4103_,
    new_n4104_, new_n4105_, new_n4106_, new_n4107_, new_n4108_, new_n4109_,
    new_n4110_, new_n4111_, new_n4112_, new_n4113_, new_n4114_, new_n4115_,
    new_n4116_, new_n4117_, new_n4118_, new_n4119_, new_n4120_, new_n4121_,
    new_n4122_, new_n4123_, new_n4124_, new_n4125_, new_n4126_, new_n4127_,
    new_n4128_, new_n4129_, new_n4130_, new_n4131_, new_n4132_, new_n4133_,
    new_n4134_, new_n4135_, new_n4136_, new_n4137_, new_n4138_, new_n4139_,
    new_n4140_, new_n4141_, new_n4142_, new_n4143_, new_n4145_, new_n4146_,
    new_n4147_, new_n4148_, new_n4149_, new_n4150_, new_n4151_, new_n4152_,
    new_n4153_, new_n4154_, new_n4155_, new_n4156_, new_n4157_, new_n4158_,
    new_n4159_, new_n4160_, new_n4161_, new_n4162_, new_n4163_, new_n4164_,
    new_n4165_, new_n4166_, new_n4167_, new_n4168_, new_n4169_, new_n4170_,
    new_n4171_, new_n4172_, new_n4173_, new_n4174_, new_n4175_, new_n4176_,
    new_n4177_, new_n4178_, new_n4179_, new_n4180_, new_n4181_, new_n4182_,
    new_n4183_, new_n4184_, new_n4185_, new_n4186_, new_n4187_, new_n4188_,
    new_n4189_, new_n4190_, new_n4191_, new_n4192_, new_n4193_, new_n4194_,
    new_n4195_, new_n4196_, new_n4197_, new_n4198_, new_n4199_, new_n4200_,
    new_n4201_, new_n4202_, new_n4203_, new_n4204_, new_n4205_, new_n4206_,
    new_n4207_, new_n4208_, new_n4209_, new_n4210_, new_n4211_, new_n4212_,
    new_n4213_, new_n4214_, new_n4215_, new_n4216_, new_n4217_, new_n4218_,
    new_n4219_, new_n4220_, new_n4221_, new_n4222_, new_n4223_, new_n4224_,
    new_n4225_, new_n4226_, new_n4227_, new_n4228_, new_n4229_, new_n4230_,
    new_n4231_, new_n4232_, new_n4233_, new_n4234_, new_n4235_, new_n4236_,
    new_n4237_, new_n4238_, new_n4239_, new_n4240_, new_n4241_, new_n4242_,
    new_n4243_, new_n4244_, new_n4245_, new_n4246_, new_n4247_, new_n4248_,
    new_n4249_, new_n4250_, new_n4251_, new_n4252_, new_n4253_, new_n4254_,
    new_n4255_, new_n4256_, new_n4257_, new_n4258_, new_n4259_, new_n4260_,
    new_n4261_, new_n4262_, new_n4263_, new_n4264_, new_n4265_, new_n4266_,
    new_n4267_, new_n4268_, new_n4269_, new_n4270_, new_n4271_, new_n4272_,
    new_n4273_, new_n4274_, new_n4275_, new_n4276_, new_n4277_, new_n4278_,
    new_n4279_, new_n4280_, new_n4281_, new_n4282_, new_n4283_, new_n4284_,
    new_n4285_, new_n4286_, new_n4287_, new_n4288_, new_n4289_, new_n4290_,
    new_n4291_, new_n4292_, new_n4293_, new_n4294_, new_n4295_, new_n4296_,
    new_n4297_, new_n4298_, new_n4299_, new_n4300_, new_n4301_, new_n4302_,
    new_n4303_, new_n4304_, new_n4305_, new_n4306_, new_n4307_, new_n4308_,
    new_n4309_, new_n4310_, new_n4311_, new_n4312_, new_n4313_, new_n4314_,
    new_n4315_, new_n4316_, new_n4317_, new_n4318_, new_n4319_, new_n4320_,
    new_n4321_, new_n4322_, new_n4323_, new_n4324_, new_n4325_, new_n4326_,
    new_n4327_, new_n4328_, new_n4329_, new_n4330_, new_n4331_, new_n4332_,
    new_n4333_, new_n4334_, new_n4335_, new_n4336_, new_n4337_, new_n4338_,
    new_n4339_, new_n4340_, new_n4341_, new_n4342_, new_n4343_, new_n4344_,
    new_n4345_, new_n4346_, new_n4347_, new_n4348_, new_n4349_, new_n4350_,
    new_n4351_, new_n4352_, new_n4353_, new_n4354_, new_n4355_, new_n4356_,
    new_n4357_, new_n4358_, new_n4359_, new_n4360_, new_n4361_, new_n4362_,
    new_n4363_, new_n4364_, new_n4365_, new_n4366_, new_n4367_, new_n4368_,
    new_n4369_, new_n4370_, new_n4371_, new_n4372_, new_n4373_, new_n4374_,
    new_n4375_, new_n4376_, new_n4377_, new_n4378_, new_n4379_, new_n4380_,
    new_n4381_, new_n4382_, new_n4383_, new_n4384_, new_n4385_, new_n4386_,
    new_n4387_, new_n4388_, new_n4389_, new_n4390_, new_n4391_, new_n4392_,
    new_n4393_, new_n4394_, new_n4395_, new_n4396_, new_n4397_, new_n4398_,
    new_n4399_, new_n4400_, new_n4401_, new_n4402_, new_n4403_, new_n4404_,
    new_n4405_, new_n4406_, new_n4407_, new_n4408_, new_n4409_, new_n4410_,
    new_n4411_, new_n4412_, new_n4413_, new_n4414_, new_n4415_, new_n4416_,
    new_n4417_, new_n4418_, new_n4419_, new_n4420_, new_n4421_, new_n4422_,
    new_n4423_, new_n4424_, new_n4425_, new_n4426_, new_n4427_, new_n4428_,
    new_n4429_, new_n4430_, new_n4431_, new_n4432_, new_n4433_, new_n4434_,
    new_n4435_, new_n4436_, new_n4437_, new_n4438_, new_n4439_, new_n4440_,
    new_n4441_, new_n4442_, new_n4443_, new_n4444_, new_n4445_, new_n4446_,
    new_n4447_, new_n4448_, new_n4449_, new_n4450_, new_n4451_, new_n4452_,
    new_n4453_, new_n4454_, new_n4455_, new_n4456_, new_n4457_, new_n4458_,
    new_n4459_, new_n4460_, new_n4461_, new_n4462_, new_n4463_, new_n4464_,
    new_n4465_, new_n4466_, new_n4467_, new_n4468_, new_n4469_, new_n4470_,
    new_n4471_, new_n4472_, new_n4473_, new_n4474_, new_n4475_, new_n4477_,
    new_n4478_, new_n4479_, new_n4480_, new_n4481_, new_n4482_, new_n4483_,
    new_n4484_, new_n4485_, new_n4486_, new_n4487_, new_n4488_, new_n4489_,
    new_n4490_, new_n4491_, new_n4492_, new_n4493_, new_n4494_, new_n4495_,
    new_n4496_, new_n4497_, new_n4498_, new_n4499_, new_n4500_, new_n4501_,
    new_n4502_, new_n4503_, new_n4504_, new_n4505_, new_n4506_, new_n4507_,
    new_n4508_, new_n4509_, new_n4510_, new_n4511_, new_n4512_, new_n4513_,
    new_n4514_, new_n4515_, new_n4516_, new_n4517_, new_n4518_, new_n4519_,
    new_n4520_, new_n4521_, new_n4522_, new_n4523_, new_n4524_, new_n4525_,
    new_n4526_, new_n4527_, new_n4528_, new_n4529_, new_n4530_, new_n4531_,
    new_n4532_, new_n4533_, new_n4534_, new_n4535_, new_n4536_, new_n4537_,
    new_n4538_, new_n4539_, new_n4540_, new_n4541_, new_n4542_, new_n4543_,
    new_n4544_, new_n4545_, new_n4546_, new_n4547_, new_n4548_, new_n4549_,
    new_n4550_, new_n4551_, new_n4552_, new_n4553_, new_n4554_, new_n4555_,
    new_n4556_, new_n4557_, new_n4558_, new_n4559_, new_n4560_, new_n4561_,
    new_n4562_, new_n4563_, new_n4564_, new_n4565_, new_n4566_, new_n4567_,
    new_n4568_, new_n4569_, new_n4570_, new_n4571_, new_n4572_, new_n4573_,
    new_n4574_, new_n4575_, new_n4576_, new_n4577_, new_n4578_, new_n4579_,
    new_n4580_, new_n4581_, new_n4582_, new_n4583_, new_n4584_, new_n4585_,
    new_n4586_, new_n4587_, new_n4588_, new_n4589_, new_n4590_, new_n4591_,
    new_n4592_, new_n4593_, new_n4594_, new_n4595_, new_n4596_, new_n4597_,
    new_n4598_, new_n4599_, new_n4600_, new_n4601_, new_n4602_, new_n4603_,
    new_n4604_, new_n4605_, new_n4606_, new_n4607_, new_n4608_, new_n4609_,
    new_n4610_, new_n4611_, new_n4612_, new_n4613_, new_n4614_, new_n4615_,
    new_n4616_, new_n4617_, new_n4618_, new_n4619_, new_n4620_, new_n4621_,
    new_n4622_, new_n4623_, new_n4624_, new_n4625_, new_n4626_, new_n4627_,
    new_n4628_, new_n4629_, new_n4630_, new_n4631_, new_n4632_, new_n4633_,
    new_n4634_, new_n4635_, new_n4636_, new_n4637_, new_n4638_, new_n4639_,
    new_n4640_, new_n4641_, new_n4642_, new_n4643_, new_n4644_, new_n4645_,
    new_n4646_, new_n4647_, new_n4648_, new_n4649_, new_n4650_, new_n4651_,
    new_n4652_, new_n4653_, new_n4654_, new_n4655_, new_n4656_, new_n4657_,
    new_n4658_, new_n4659_, new_n4660_, new_n4661_, new_n4662_, new_n4663_,
    new_n4664_, new_n4665_, new_n4666_, new_n4667_, new_n4668_, new_n4669_,
    new_n4670_, new_n4671_, new_n4672_, new_n4673_, new_n4674_, new_n4675_,
    new_n4676_, new_n4677_, new_n4678_, new_n4679_, new_n4680_, new_n4681_,
    new_n4682_, new_n4683_, new_n4684_, new_n4685_, new_n4686_, new_n4687_,
    new_n4688_, new_n4689_, new_n4690_, new_n4691_, new_n4692_, new_n4693_,
    new_n4694_, new_n4695_, new_n4696_, new_n4697_, new_n4698_, new_n4699_,
    new_n4700_, new_n4701_, new_n4702_, new_n4703_, new_n4704_, new_n4705_,
    new_n4706_, new_n4707_, new_n4708_, new_n4709_, new_n4710_, new_n4711_,
    new_n4712_, new_n4713_, new_n4714_, new_n4715_, new_n4716_, new_n4717_,
    new_n4718_, new_n4719_, new_n4720_, new_n4721_, new_n4722_, new_n4723_,
    new_n4724_, new_n4725_, new_n4726_, new_n4727_, new_n4728_, new_n4729_,
    new_n4730_, new_n4731_, new_n4732_, new_n4733_, new_n4734_, new_n4735_,
    new_n4736_, new_n4737_, new_n4738_, new_n4739_, new_n4740_, new_n4741_,
    new_n4742_, new_n4743_, new_n4744_, new_n4745_, new_n4746_, new_n4747_,
    new_n4748_, new_n4749_, new_n4750_, new_n4751_, new_n4752_, new_n4753_,
    new_n4754_, new_n4755_, new_n4756_, new_n4757_, new_n4758_, new_n4759_,
    new_n4760_, new_n4761_, new_n4762_, new_n4763_, new_n4764_, new_n4765_,
    new_n4766_, new_n4767_, new_n4768_, new_n4769_, new_n4770_, new_n4771_,
    new_n4772_, new_n4773_, new_n4774_, new_n4775_, new_n4776_, new_n4777_,
    new_n4778_, new_n4779_, new_n4780_, new_n4781_, new_n4782_, new_n4783_,
    new_n4784_, new_n4785_, new_n4786_, new_n4787_, new_n4788_, new_n4789_,
    new_n4790_, new_n4791_, new_n4792_, new_n4793_, new_n4794_, new_n4795_,
    new_n4796_, new_n4797_, new_n4798_, new_n4799_, new_n4800_, new_n4801_,
    new_n4802_, new_n4803_, new_n4804_, new_n4805_, new_n4806_, new_n4807_,
    new_n4808_, new_n4809_, new_n4810_, new_n4811_, new_n4812_, new_n4813_,
    new_n4815_, new_n4816_, new_n4817_, new_n4818_, new_n4819_, new_n4820_,
    new_n4821_, new_n4822_, new_n4823_, new_n4824_, new_n4825_, new_n4826_,
    new_n4827_, new_n4828_, new_n4829_, new_n4830_, new_n4831_, new_n4832_,
    new_n4833_, new_n4834_, new_n4835_, new_n4836_, new_n4837_, new_n4838_,
    new_n4839_, new_n4840_, new_n4841_, new_n4842_, new_n4843_, new_n4844_,
    new_n4845_, new_n4846_, new_n4847_, new_n4848_, new_n4849_, new_n4850_,
    new_n4851_, new_n4852_, new_n4853_, new_n4854_, new_n4855_, new_n4856_,
    new_n4857_, new_n4858_, new_n4859_, new_n4860_, new_n4861_, new_n4862_,
    new_n4863_, new_n4864_, new_n4865_, new_n4866_, new_n4867_, new_n4868_,
    new_n4869_, new_n4870_, new_n4871_, new_n4872_, new_n4873_, new_n4874_,
    new_n4875_, new_n4876_, new_n4877_, new_n4878_, new_n4879_, new_n4880_,
    new_n4881_, new_n4882_, new_n4883_, new_n4884_, new_n4885_, new_n4886_,
    new_n4887_, new_n4888_, new_n4889_, new_n4890_, new_n4891_, new_n4892_,
    new_n4893_, new_n4894_, new_n4895_, new_n4896_, new_n4897_, new_n4898_,
    new_n4899_, new_n4900_, new_n4901_, new_n4902_, new_n4903_, new_n4904_,
    new_n4905_, new_n4906_, new_n4907_, new_n4908_, new_n4909_, new_n4910_,
    new_n4911_, new_n4912_, new_n4913_, new_n4914_, new_n4915_, new_n4916_,
    new_n4917_, new_n4918_, new_n4919_, new_n4920_, new_n4921_, new_n4922_,
    new_n4923_, new_n4924_, new_n4925_, new_n4926_, new_n4927_, new_n4928_,
    new_n4929_, new_n4930_, new_n4931_, new_n4932_, new_n4933_, new_n4934_,
    new_n4935_, new_n4936_, new_n4937_, new_n4938_, new_n4939_, new_n4940_,
    new_n4941_, new_n4942_, new_n4943_, new_n4944_, new_n4945_, new_n4946_,
    new_n4947_, new_n4948_, new_n4949_, new_n4950_, new_n4951_, new_n4952_,
    new_n4953_, new_n4954_, new_n4955_, new_n4956_, new_n4957_, new_n4958_,
    new_n4959_, new_n4960_, new_n4961_, new_n4962_, new_n4963_, new_n4964_,
    new_n4965_, new_n4966_, new_n4967_, new_n4968_, new_n4969_, new_n4970_,
    new_n4971_, new_n4972_, new_n4973_, new_n4974_, new_n4975_, new_n4976_,
    new_n4977_, new_n4978_, new_n4979_, new_n4980_, new_n4981_, new_n4982_,
    new_n4983_, new_n4984_, new_n4985_, new_n4986_, new_n4987_, new_n4988_,
    new_n4989_, new_n4990_, new_n4991_, new_n4992_, new_n4993_, new_n4994_,
    new_n4995_, new_n4996_, new_n4997_, new_n4998_, new_n4999_, new_n5000_,
    new_n5001_, new_n5002_, new_n5003_, new_n5004_, new_n5005_, new_n5006_,
    new_n5007_, new_n5008_, new_n5009_, new_n5010_, new_n5011_, new_n5012_,
    new_n5013_, new_n5014_, new_n5015_, new_n5016_, new_n5017_, new_n5018_,
    new_n5019_, new_n5020_, new_n5021_, new_n5022_, new_n5023_, new_n5024_,
    new_n5025_, new_n5026_, new_n5027_, new_n5028_, new_n5029_, new_n5030_,
    new_n5031_, new_n5032_, new_n5033_, new_n5034_, new_n5035_, new_n5036_,
    new_n5037_, new_n5038_, new_n5039_, new_n5040_, new_n5041_, new_n5042_,
    new_n5043_, new_n5044_, new_n5045_, new_n5046_, new_n5047_, new_n5048_,
    new_n5049_, new_n5050_, new_n5051_, new_n5052_, new_n5053_, new_n5054_,
    new_n5055_, new_n5056_, new_n5057_, new_n5058_, new_n5059_, new_n5060_,
    new_n5061_, new_n5062_, new_n5063_, new_n5064_, new_n5065_, new_n5066_,
    new_n5067_, new_n5068_, new_n5069_, new_n5070_, new_n5071_, new_n5072_,
    new_n5073_, new_n5074_, new_n5075_, new_n5076_, new_n5077_, new_n5078_,
    new_n5079_, new_n5080_, new_n5081_, new_n5082_, new_n5083_, new_n5084_,
    new_n5085_, new_n5086_, new_n5087_, new_n5088_, new_n5089_, new_n5090_,
    new_n5091_, new_n5092_, new_n5093_, new_n5094_, new_n5095_, new_n5096_,
    new_n5097_, new_n5098_, new_n5099_, new_n5100_, new_n5101_, new_n5102_,
    new_n5103_, new_n5104_, new_n5105_, new_n5106_, new_n5107_, new_n5108_,
    new_n5109_, new_n5110_, new_n5111_, new_n5112_, new_n5113_, new_n5114_,
    new_n5115_, new_n5116_, new_n5117_, new_n5118_, new_n5119_, new_n5120_,
    new_n5121_, new_n5122_, new_n5123_, new_n5124_, new_n5125_, new_n5126_,
    new_n5127_, new_n5128_, new_n5129_, new_n5130_, new_n5131_, new_n5132_,
    new_n5133_, new_n5134_, new_n5135_, new_n5136_, new_n5137_, new_n5138_,
    new_n5139_, new_n5140_, new_n5141_, new_n5142_, new_n5143_, new_n5144_,
    new_n5145_, new_n5146_, new_n5147_, new_n5148_, new_n5149_, new_n5150_,
    new_n5151_, new_n5152_, new_n5153_, new_n5154_, new_n5155_, new_n5156_,
    new_n5157_, new_n5158_, new_n5159_, new_n5160_, new_n5161_, new_n5162_,
    new_n5163_, new_n5164_, new_n5165_, new_n5166_, new_n5167_, new_n5168_,
    new_n5169_, new_n5170_, new_n5171_, new_n5172_, new_n5174_, new_n5175_,
    new_n5176_, new_n5177_, new_n5178_, new_n5179_, new_n5180_, new_n5181_,
    new_n5182_, new_n5183_, new_n5184_, new_n5185_, new_n5186_, new_n5187_,
    new_n5188_, new_n5189_, new_n5190_, new_n5191_, new_n5192_, new_n5193_,
    new_n5194_, new_n5195_, new_n5196_, new_n5197_, new_n5198_, new_n5199_,
    new_n5200_, new_n5201_, new_n5202_, new_n5203_, new_n5204_, new_n5205_,
    new_n5206_, new_n5207_, new_n5208_, new_n5209_, new_n5210_, new_n5211_,
    new_n5212_, new_n5213_, new_n5214_, new_n5215_, new_n5216_, new_n5217_,
    new_n5218_, new_n5219_, new_n5220_, new_n5221_, new_n5222_, new_n5223_,
    new_n5224_, new_n5225_, new_n5226_, new_n5227_, new_n5228_, new_n5229_,
    new_n5230_, new_n5231_, new_n5232_, new_n5233_, new_n5234_, new_n5235_,
    new_n5236_, new_n5237_, new_n5238_, new_n5239_, new_n5240_, new_n5241_,
    new_n5242_, new_n5243_, new_n5244_, new_n5245_, new_n5246_, new_n5247_,
    new_n5248_, new_n5249_, new_n5250_, new_n5251_, new_n5252_, new_n5253_,
    new_n5254_, new_n5255_, new_n5256_, new_n5257_, new_n5258_, new_n5259_,
    new_n5260_, new_n5261_, new_n5262_, new_n5263_, new_n5264_, new_n5265_,
    new_n5266_, new_n5267_, new_n5268_, new_n5269_, new_n5270_, new_n5271_,
    new_n5272_, new_n5273_, new_n5274_, new_n5275_, new_n5276_, new_n5277_,
    new_n5278_, new_n5279_, new_n5280_, new_n5281_, new_n5282_, new_n5283_,
    new_n5284_, new_n5285_, new_n5286_, new_n5287_, new_n5288_, new_n5289_,
    new_n5290_, new_n5291_, new_n5292_, new_n5293_, new_n5294_, new_n5295_,
    new_n5296_, new_n5297_, new_n5298_, new_n5299_, new_n5300_, new_n5301_,
    new_n5302_, new_n5303_, new_n5304_, new_n5305_, new_n5306_, new_n5307_,
    new_n5308_, new_n5309_, new_n5310_, new_n5311_, new_n5312_, new_n5313_,
    new_n5314_, new_n5315_, new_n5316_, new_n5317_, new_n5318_, new_n5319_,
    new_n5320_, new_n5321_, new_n5322_, new_n5323_, new_n5324_, new_n5325_,
    new_n5326_, new_n5327_, new_n5328_, new_n5329_, new_n5330_, new_n5331_,
    new_n5332_, new_n5333_, new_n5334_, new_n5335_, new_n5336_, new_n5337_,
    new_n5338_, new_n5339_, new_n5340_, new_n5341_, new_n5342_, new_n5343_,
    new_n5344_, new_n5345_, new_n5346_, new_n5347_, new_n5348_, new_n5349_,
    new_n5350_, new_n5351_, new_n5352_, new_n5353_, new_n5354_, new_n5355_,
    new_n5356_, new_n5357_, new_n5358_, new_n5359_, new_n5360_, new_n5361_,
    new_n5362_, new_n5363_, new_n5364_, new_n5365_, new_n5366_, new_n5367_,
    new_n5368_, new_n5369_, new_n5370_, new_n5371_, new_n5372_, new_n5373_,
    new_n5374_, new_n5375_, new_n5376_, new_n5377_, new_n5378_, new_n5379_,
    new_n5380_, new_n5381_, new_n5382_, new_n5383_, new_n5384_, new_n5385_,
    new_n5386_, new_n5387_, new_n5388_, new_n5389_, new_n5390_, new_n5391_,
    new_n5392_, new_n5393_, new_n5394_, new_n5395_, new_n5396_, new_n5397_,
    new_n5398_, new_n5399_, new_n5400_, new_n5401_, new_n5402_, new_n5403_,
    new_n5404_, new_n5405_, new_n5406_, new_n5407_, new_n5408_, new_n5409_,
    new_n5410_, new_n5411_, new_n5412_, new_n5413_, new_n5414_, new_n5415_,
    new_n5416_, new_n5417_, new_n5418_, new_n5419_, new_n5420_, new_n5421_,
    new_n5422_, new_n5423_, new_n5424_, new_n5425_, new_n5426_, new_n5427_,
    new_n5428_, new_n5429_, new_n5430_, new_n5431_, new_n5432_, new_n5433_,
    new_n5434_, new_n5435_, new_n5436_, new_n5437_, new_n5438_, new_n5439_,
    new_n5440_, new_n5441_, new_n5442_, new_n5443_, new_n5444_, new_n5445_,
    new_n5446_, new_n5447_, new_n5448_, new_n5449_, new_n5450_, new_n5451_,
    new_n5452_, new_n5453_, new_n5454_, new_n5455_, new_n5456_, new_n5457_,
    new_n5458_, new_n5459_, new_n5460_, new_n5461_, new_n5462_, new_n5463_,
    new_n5464_, new_n5465_, new_n5466_, new_n5467_, new_n5468_, new_n5469_,
    new_n5470_, new_n5471_, new_n5472_, new_n5473_, new_n5474_, new_n5475_,
    new_n5476_, new_n5477_, new_n5478_, new_n5479_, new_n5480_, new_n5481_,
    new_n5482_, new_n5483_, new_n5484_, new_n5485_, new_n5486_, new_n5487_,
    new_n5488_, new_n5489_, new_n5490_, new_n5491_, new_n5492_, new_n5493_,
    new_n5494_, new_n5495_, new_n5496_, new_n5497_, new_n5498_, new_n5499_,
    new_n5500_, new_n5501_, new_n5502_, new_n5503_, new_n5504_, new_n5505_,
    new_n5506_, new_n5507_, new_n5508_, new_n5509_, new_n5510_, new_n5511_,
    new_n5512_, new_n5513_, new_n5514_, new_n5515_, new_n5516_, new_n5517_,
    new_n5518_, new_n5519_, new_n5520_, new_n5521_, new_n5522_, new_n5523_,
    new_n5524_, new_n5525_, new_n5526_, new_n5527_, new_n5528_, new_n5529_,
    new_n5530_, new_n5531_, new_n5532_, new_n5533_, new_n5534_, new_n5535_,
    new_n5536_, new_n5537_, new_n5538_, new_n5539_, new_n5540_, new_n5541_,
    new_n5542_, new_n5543_, new_n5544_, new_n5545_, new_n5546_, new_n5548_,
    new_n5549_, new_n5550_, new_n5551_, new_n5552_, new_n5553_, new_n5554_,
    new_n5555_, new_n5556_, new_n5557_, new_n5558_, new_n5559_, new_n5560_,
    new_n5561_, new_n5562_, new_n5563_, new_n5564_, new_n5565_, new_n5566_,
    new_n5567_, new_n5568_, new_n5569_, new_n5570_, new_n5571_, new_n5572_,
    new_n5573_, new_n5574_, new_n5575_, new_n5576_, new_n5577_, new_n5578_,
    new_n5579_, new_n5580_, new_n5581_, new_n5582_, new_n5583_, new_n5584_,
    new_n5585_, new_n5586_, new_n5587_, new_n5588_, new_n5589_, new_n5590_,
    new_n5591_, new_n5592_, new_n5593_, new_n5594_, new_n5595_, new_n5596_,
    new_n5597_, new_n5598_, new_n5599_, new_n5600_, new_n5601_, new_n5602_,
    new_n5603_, new_n5604_, new_n5605_, new_n5606_, new_n5607_, new_n5608_,
    new_n5609_, new_n5610_, new_n5611_, new_n5612_, new_n5613_, new_n5614_,
    new_n5615_, new_n5616_, new_n5617_, new_n5618_, new_n5619_, new_n5620_,
    new_n5621_, new_n5622_, new_n5623_, new_n5624_, new_n5625_, new_n5626_,
    new_n5627_, new_n5628_, new_n5629_, new_n5630_, new_n5631_, new_n5632_,
    new_n5633_, new_n5634_, new_n5635_, new_n5636_, new_n5637_, new_n5638_,
    new_n5639_, new_n5640_, new_n5641_, new_n5642_, new_n5643_, new_n5644_,
    new_n5645_, new_n5646_, new_n5647_, new_n5648_, new_n5649_, new_n5650_,
    new_n5651_, new_n5652_, new_n5653_, new_n5654_, new_n5655_, new_n5656_,
    new_n5657_, new_n5658_, new_n5659_, new_n5660_, new_n5661_, new_n5662_,
    new_n5663_, new_n5664_, new_n5665_, new_n5666_, new_n5667_, new_n5668_,
    new_n5669_, new_n5670_, new_n5671_, new_n5672_, new_n5673_, new_n5674_,
    new_n5675_, new_n5676_, new_n5677_, new_n5678_, new_n5679_, new_n5680_,
    new_n5681_, new_n5682_, new_n5683_, new_n5684_, new_n5685_, new_n5686_,
    new_n5687_, new_n5688_, new_n5689_, new_n5690_, new_n5691_, new_n5692_,
    new_n5693_, new_n5694_, new_n5695_, new_n5696_, new_n5697_, new_n5698_,
    new_n5699_, new_n5700_, new_n5701_, new_n5702_, new_n5703_, new_n5704_,
    new_n5705_, new_n5706_, new_n5707_, new_n5708_, new_n5709_, new_n5710_,
    new_n5711_, new_n5712_, new_n5713_, new_n5714_, new_n5715_, new_n5716_,
    new_n5717_, new_n5718_, new_n5719_, new_n5720_, new_n5721_, new_n5722_,
    new_n5723_, new_n5724_, new_n5725_, new_n5726_, new_n5727_, new_n5728_,
    new_n5729_, new_n5730_, new_n5731_, new_n5732_, new_n5733_, new_n5734_,
    new_n5735_, new_n5736_, new_n5737_, new_n5738_, new_n5739_, new_n5740_,
    new_n5741_, new_n5742_, new_n5743_, new_n5744_, new_n5745_, new_n5746_,
    new_n5747_, new_n5748_, new_n5749_, new_n5750_, new_n5751_, new_n5752_,
    new_n5753_, new_n5754_, new_n5755_, new_n5756_, new_n5757_, new_n5758_,
    new_n5759_, new_n5760_, new_n5761_, new_n5762_, new_n5763_, new_n5764_,
    new_n5765_, new_n5766_, new_n5767_, new_n5768_, new_n5769_, new_n5770_,
    new_n5771_, new_n5772_, new_n5773_, new_n5774_, new_n5775_, new_n5776_,
    new_n5777_, new_n5778_, new_n5779_, new_n5780_, new_n5781_, new_n5782_,
    new_n5783_, new_n5784_, new_n5785_, new_n5786_, new_n5787_, new_n5788_,
    new_n5789_, new_n5790_, new_n5791_, new_n5792_, new_n5793_, new_n5794_,
    new_n5795_, new_n5796_, new_n5797_, new_n5798_, new_n5799_, new_n5800_,
    new_n5801_, new_n5802_, new_n5803_, new_n5804_, new_n5805_, new_n5806_,
    new_n5807_, new_n5808_, new_n5809_, new_n5810_, new_n5811_, new_n5812_,
    new_n5813_, new_n5814_, new_n5815_, new_n5816_, new_n5817_, new_n5818_,
    new_n5819_, new_n5820_, new_n5821_, new_n5822_, new_n5823_, new_n5824_,
    new_n5825_, new_n5826_, new_n5827_, new_n5828_, new_n5829_, new_n5830_,
    new_n5831_, new_n5832_, new_n5833_, new_n5834_, new_n5835_, new_n5836_,
    new_n5837_, new_n5838_, new_n5839_, new_n5840_, new_n5841_, new_n5842_,
    new_n5843_, new_n5844_, new_n5845_, new_n5846_, new_n5847_, new_n5848_,
    new_n5849_, new_n5850_, new_n5851_, new_n5852_, new_n5853_, new_n5854_,
    new_n5855_, new_n5856_, new_n5857_, new_n5858_, new_n5859_, new_n5860_,
    new_n5861_, new_n5862_, new_n5863_, new_n5864_, new_n5865_, new_n5866_,
    new_n5867_, new_n5868_, new_n5869_, new_n5870_, new_n5871_, new_n5872_,
    new_n5873_, new_n5874_, new_n5875_, new_n5876_, new_n5877_, new_n5878_,
    new_n5879_, new_n5880_, new_n5881_, new_n5882_, new_n5883_, new_n5884_,
    new_n5885_, new_n5886_, new_n5887_, new_n5888_, new_n5889_, new_n5890_,
    new_n5891_, new_n5892_, new_n5893_, new_n5894_, new_n5895_, new_n5896_,
    new_n5897_, new_n5898_, new_n5899_, new_n5900_, new_n5901_, new_n5902_,
    new_n5903_, new_n5904_, new_n5905_, new_n5906_, new_n5907_, new_n5908_,
    new_n5909_, new_n5910_, new_n5911_, new_n5912_, new_n5913_, new_n5914_,
    new_n5915_, new_n5916_, new_n5917_, new_n5918_, new_n5919_, new_n5920_,
    new_n5921_, new_n5922_, new_n5923_, new_n5924_, new_n5925_, new_n5926_,
    new_n5928_, new_n5929_, new_n5930_, new_n5931_, new_n5932_, new_n5933_,
    new_n5934_, new_n5935_, new_n5936_, new_n5937_, new_n5938_, new_n5939_,
    new_n5940_, new_n5941_, new_n5942_, new_n5943_, new_n5944_, new_n5945_,
    new_n5946_, new_n5947_, new_n5948_, new_n5949_, new_n5950_, new_n5951_,
    new_n5952_, new_n5953_, new_n5954_, new_n5955_, new_n5956_, new_n5957_,
    new_n5958_, new_n5959_, new_n5960_, new_n5961_, new_n5962_, new_n5963_,
    new_n5964_, new_n5965_, new_n5966_, new_n5967_, new_n5968_, new_n5969_,
    new_n5970_, new_n5971_, new_n5972_, new_n5973_, new_n5974_, new_n5975_,
    new_n5976_, new_n5977_, new_n5978_, new_n5979_, new_n5980_, new_n5981_,
    new_n5982_, new_n5983_, new_n5984_, new_n5985_, new_n5986_, new_n5987_,
    new_n5988_, new_n5989_, new_n5990_, new_n5991_, new_n5992_, new_n5993_,
    new_n5994_, new_n5995_, new_n5996_, new_n5997_, new_n5998_, new_n5999_,
    new_n6000_, new_n6001_, new_n6002_, new_n6003_, new_n6004_, new_n6005_,
    new_n6006_, new_n6007_, new_n6008_, new_n6009_, new_n6010_, new_n6011_,
    new_n6012_, new_n6013_, new_n6014_, new_n6015_, new_n6016_, new_n6017_,
    new_n6018_, new_n6019_, new_n6020_, new_n6021_, new_n6022_, new_n6023_,
    new_n6024_, new_n6025_, new_n6026_, new_n6027_, new_n6028_, new_n6029_,
    new_n6030_, new_n6031_, new_n6032_, new_n6033_, new_n6034_, new_n6035_,
    new_n6036_, new_n6037_, new_n6038_, new_n6039_, new_n6040_, new_n6041_,
    new_n6042_, new_n6043_, new_n6044_, new_n6045_, new_n6046_, new_n6047_,
    new_n6048_, new_n6049_, new_n6050_, new_n6051_, new_n6052_, new_n6053_,
    new_n6054_, new_n6055_, new_n6056_, new_n6057_, new_n6058_, new_n6059_,
    new_n6060_, new_n6061_, new_n6062_, new_n6063_, new_n6064_, new_n6065_,
    new_n6066_, new_n6067_, new_n6068_, new_n6069_, new_n6070_, new_n6071_,
    new_n6072_, new_n6073_, new_n6074_, new_n6075_, new_n6076_, new_n6077_,
    new_n6078_, new_n6079_, new_n6080_, new_n6081_, new_n6082_, new_n6083_,
    new_n6084_, new_n6085_, new_n6086_, new_n6087_, new_n6088_, new_n6089_,
    new_n6090_, new_n6091_, new_n6092_, new_n6093_, new_n6094_, new_n6095_,
    new_n6096_, new_n6097_, new_n6098_, new_n6099_, new_n6100_, new_n6101_,
    new_n6102_, new_n6103_, new_n6104_, new_n6105_, new_n6106_, new_n6107_,
    new_n6108_, new_n6109_, new_n6110_, new_n6111_, new_n6112_, new_n6113_,
    new_n6114_, new_n6115_, new_n6116_, new_n6117_, new_n6118_, new_n6119_,
    new_n6120_, new_n6121_, new_n6122_, new_n6123_, new_n6124_, new_n6125_,
    new_n6126_, new_n6127_, new_n6128_, new_n6129_, new_n6130_, new_n6131_,
    new_n6132_, new_n6133_, new_n6134_, new_n6135_, new_n6136_, new_n6137_,
    new_n6138_, new_n6139_, new_n6140_, new_n6141_, new_n6142_, new_n6143_,
    new_n6144_, new_n6145_, new_n6146_, new_n6147_, new_n6148_, new_n6149_,
    new_n6150_, new_n6151_, new_n6152_, new_n6153_, new_n6154_, new_n6155_,
    new_n6156_, new_n6157_, new_n6158_, new_n6159_, new_n6160_, new_n6161_,
    new_n6162_, new_n6163_, new_n6164_, new_n6165_, new_n6166_, new_n6167_,
    new_n6168_, new_n6169_, new_n6170_, new_n6171_, new_n6172_, new_n6173_,
    new_n6174_, new_n6175_, new_n6176_, new_n6177_, new_n6178_, new_n6179_,
    new_n6180_, new_n6181_, new_n6182_, new_n6183_, new_n6184_, new_n6185_,
    new_n6186_, new_n6187_, new_n6188_, new_n6189_, new_n6190_, new_n6191_,
    new_n6192_, new_n6193_, new_n6194_, new_n6195_, new_n6196_, new_n6197_,
    new_n6198_, new_n6199_, new_n6200_, new_n6201_, new_n6202_, new_n6203_,
    new_n6204_, new_n6205_, new_n6206_, new_n6207_, new_n6208_, new_n6209_,
    new_n6210_, new_n6211_, new_n6212_, new_n6213_, new_n6214_, new_n6215_,
    new_n6216_, new_n6217_, new_n6218_, new_n6219_, new_n6220_, new_n6221_,
    new_n6222_, new_n6223_, new_n6224_, new_n6225_, new_n6226_, new_n6227_,
    new_n6228_, new_n6229_, new_n6230_, new_n6231_, new_n6232_, new_n6233_,
    new_n6234_, new_n6235_, new_n6236_, new_n6237_, new_n6238_, new_n6239_,
    new_n6240_, new_n6241_, new_n6242_, new_n6243_, new_n6244_, new_n6245_,
    new_n6246_, new_n6247_, new_n6248_, new_n6249_, new_n6250_, new_n6251_,
    new_n6252_, new_n6253_, new_n6254_, new_n6255_, new_n6256_, new_n6257_,
    new_n6258_, new_n6259_, new_n6260_, new_n6261_, new_n6262_, new_n6263_,
    new_n6264_, new_n6265_, new_n6266_, new_n6267_, new_n6268_, new_n6269_,
    new_n6270_, new_n6271_, new_n6272_, new_n6273_, new_n6274_, new_n6275_,
    new_n6276_, new_n6277_, new_n6278_, new_n6279_, new_n6280_, new_n6281_,
    new_n6282_, new_n6283_, new_n6284_, new_n6285_, new_n6286_, new_n6287_,
    new_n6288_, new_n6289_, new_n6290_, new_n6291_, new_n6292_, new_n6293_,
    new_n6294_, new_n6295_, new_n6296_, new_n6297_, new_n6298_, new_n6299_,
    new_n6300_, new_n6301_, new_n6302_, new_n6303_, new_n6304_, new_n6305_,
    new_n6306_, new_n6307_, new_n6308_, new_n6309_, new_n6310_, new_n6311_,
    new_n6312_, new_n6313_, new_n6314_, new_n6315_, new_n6316_, new_n6317_,
    new_n6318_, new_n6319_, new_n6320_, new_n6321_, new_n6322_, new_n6323_,
    new_n6324_, new_n6326_, new_n6327_, new_n6328_, new_n6329_, new_n6330_,
    new_n6331_, new_n6332_, new_n6333_, new_n6334_, new_n6335_, new_n6336_,
    new_n6337_, new_n6338_, new_n6339_, new_n6340_, new_n6341_, new_n6342_,
    new_n6343_, new_n6344_, new_n6345_, new_n6346_, new_n6347_, new_n6348_,
    new_n6349_, new_n6350_, new_n6351_, new_n6352_, new_n6353_, new_n6354_,
    new_n6355_, new_n6356_, new_n6357_, new_n6358_, new_n6359_, new_n6360_,
    new_n6361_, new_n6362_, new_n6363_, new_n6364_, new_n6365_, new_n6366_,
    new_n6367_, new_n6368_, new_n6369_, new_n6370_, new_n6371_, new_n6372_,
    new_n6373_, new_n6374_, new_n6375_, new_n6376_, new_n6377_, new_n6378_,
    new_n6379_, new_n6380_, new_n6381_, new_n6382_, new_n6383_, new_n6384_,
    new_n6385_, new_n6386_, new_n6387_, new_n6388_, new_n6389_, new_n6390_,
    new_n6391_, new_n6392_, new_n6393_, new_n6394_, new_n6395_, new_n6396_,
    new_n6397_, new_n6398_, new_n6399_, new_n6400_, new_n6401_, new_n6402_,
    new_n6403_, new_n6404_, new_n6405_, new_n6406_, new_n6407_, new_n6408_,
    new_n6409_, new_n6410_, new_n6411_, new_n6412_, new_n6413_, new_n6414_,
    new_n6415_, new_n6416_, new_n6417_, new_n6418_, new_n6419_, new_n6420_,
    new_n6421_, new_n6422_, new_n6423_, new_n6424_, new_n6425_, new_n6426_,
    new_n6427_, new_n6428_, new_n6429_, new_n6430_, new_n6431_, new_n6432_,
    new_n6433_, new_n6434_, new_n6435_, new_n6436_, new_n6437_, new_n6438_,
    new_n6439_, new_n6440_, new_n6441_, new_n6442_, new_n6443_, new_n6444_,
    new_n6445_, new_n6446_, new_n6447_, new_n6448_, new_n6449_, new_n6450_,
    new_n6451_, new_n6452_, new_n6453_, new_n6454_, new_n6455_, new_n6456_,
    new_n6457_, new_n6458_, new_n6459_, new_n6460_, new_n6461_, new_n6462_,
    new_n6463_, new_n6464_, new_n6465_, new_n6466_, new_n6467_, new_n6468_,
    new_n6469_, new_n6470_, new_n6471_, new_n6472_, new_n6473_, new_n6474_,
    new_n6475_, new_n6476_, new_n6477_, new_n6478_, new_n6479_, new_n6480_,
    new_n6481_, new_n6482_, new_n6483_, new_n6484_, new_n6485_, new_n6486_,
    new_n6487_, new_n6488_, new_n6489_, new_n6490_, new_n6491_, new_n6492_,
    new_n6493_, new_n6494_, new_n6495_, new_n6496_, new_n6497_, new_n6498_,
    new_n6499_, new_n6500_, new_n6501_, new_n6502_, new_n6503_, new_n6504_,
    new_n6505_, new_n6506_, new_n6507_, new_n6508_, new_n6509_, new_n6510_,
    new_n6511_, new_n6512_, new_n6513_, new_n6514_, new_n6515_, new_n6516_,
    new_n6517_, new_n6518_, new_n6519_, new_n6520_, new_n6521_, new_n6522_,
    new_n6523_, new_n6524_, new_n6525_, new_n6526_, new_n6527_, new_n6528_,
    new_n6529_, new_n6530_, new_n6531_, new_n6532_, new_n6533_, new_n6534_,
    new_n6535_, new_n6536_, new_n6537_, new_n6538_, new_n6539_, new_n6540_,
    new_n6541_, new_n6542_, new_n6543_, new_n6544_, new_n6545_, new_n6546_,
    new_n6547_, new_n6548_, new_n6549_, new_n6550_, new_n6551_, new_n6552_,
    new_n6553_, new_n6554_, new_n6555_, new_n6556_, new_n6557_, new_n6558_,
    new_n6559_, new_n6560_, new_n6561_, new_n6562_, new_n6563_, new_n6564_,
    new_n6565_, new_n6566_, new_n6567_, new_n6568_, new_n6569_, new_n6570_,
    new_n6571_, new_n6572_, new_n6573_, new_n6574_, new_n6575_, new_n6576_,
    new_n6577_, new_n6578_, new_n6579_, new_n6580_, new_n6581_, new_n6582_,
    new_n6583_, new_n6584_, new_n6585_, new_n6586_, new_n6587_, new_n6588_,
    new_n6589_, new_n6590_, new_n6591_, new_n6592_, new_n6593_, new_n6594_,
    new_n6595_, new_n6596_, new_n6597_, new_n6598_, new_n6599_, new_n6600_,
    new_n6601_, new_n6602_, new_n6603_, new_n6604_, new_n6605_, new_n6606_,
    new_n6607_, new_n6608_, new_n6609_, new_n6610_, new_n6611_, new_n6612_,
    new_n6613_, new_n6614_, new_n6615_, new_n6616_, new_n6617_, new_n6618_,
    new_n6619_, new_n6620_, new_n6621_, new_n6622_, new_n6623_, new_n6624_,
    new_n6625_, new_n6626_, new_n6627_, new_n6628_, new_n6629_, new_n6630_,
    new_n6631_, new_n6632_, new_n6633_, new_n6634_, new_n6635_, new_n6636_,
    new_n6637_, new_n6638_, new_n6639_, new_n6640_, new_n6641_, new_n6642_,
    new_n6643_, new_n6644_, new_n6645_, new_n6646_, new_n6647_, new_n6648_,
    new_n6649_, new_n6650_, new_n6651_, new_n6652_, new_n6653_, new_n6654_,
    new_n6655_, new_n6656_, new_n6657_, new_n6658_, new_n6659_, new_n6660_,
    new_n6661_, new_n6662_, new_n6663_, new_n6664_, new_n6665_, new_n6666_,
    new_n6667_, new_n6668_, new_n6669_, new_n6670_, new_n6671_, new_n6672_,
    new_n6673_, new_n6674_, new_n6675_, new_n6676_, new_n6677_, new_n6678_,
    new_n6679_, new_n6680_, new_n6681_, new_n6682_, new_n6683_, new_n6684_,
    new_n6685_, new_n6686_, new_n6687_, new_n6688_, new_n6689_, new_n6690_,
    new_n6691_, new_n6692_, new_n6693_, new_n6694_, new_n6695_, new_n6696_,
    new_n6697_, new_n6698_, new_n6699_, new_n6700_, new_n6701_, new_n6702_,
    new_n6703_, new_n6704_, new_n6705_, new_n6706_, new_n6707_, new_n6708_,
    new_n6709_, new_n6710_, new_n6711_, new_n6712_, new_n6713_, new_n6714_,
    new_n6715_, new_n6716_, new_n6717_, new_n6718_, new_n6719_, new_n6720_,
    new_n6721_, new_n6722_, new_n6723_, new_n6724_, new_n6725_, new_n6726_,
    new_n6727_, new_n6728_, new_n6729_, new_n6730_, new_n6731_, new_n6732_,
    new_n6733_, new_n6734_, new_n6735_, new_n6736_, new_n6737_, new_n6738_,
    new_n6739_, new_n6741_, new_n6742_, new_n6743_, new_n6744_, new_n6745_,
    new_n6746_, new_n6747_, new_n6748_, new_n6749_, new_n6750_, new_n6751_,
    new_n6752_, new_n6753_, new_n6754_, new_n6755_, new_n6756_, new_n6757_,
    new_n6758_, new_n6759_, new_n6760_, new_n6761_, new_n6762_, new_n6763_,
    new_n6764_, new_n6765_, new_n6766_, new_n6767_, new_n6768_, new_n6769_,
    new_n6770_, new_n6771_, new_n6772_, new_n6773_, new_n6774_, new_n6775_,
    new_n6776_, new_n6777_, new_n6778_, new_n6779_, new_n6780_, new_n6781_,
    new_n6782_, new_n6783_, new_n6784_, new_n6785_, new_n6786_, new_n6787_,
    new_n6788_, new_n6789_, new_n6790_, new_n6791_, new_n6792_, new_n6793_,
    new_n6794_, new_n6795_, new_n6796_, new_n6797_, new_n6798_, new_n6799_,
    new_n6800_, new_n6801_, new_n6802_, new_n6803_, new_n6804_, new_n6805_,
    new_n6806_, new_n6807_, new_n6808_, new_n6809_, new_n6810_, new_n6811_,
    new_n6812_, new_n6813_, new_n6814_, new_n6815_, new_n6816_, new_n6817_,
    new_n6818_, new_n6819_, new_n6820_, new_n6821_, new_n6822_, new_n6823_,
    new_n6824_, new_n6825_, new_n6826_, new_n6827_, new_n6828_, new_n6829_,
    new_n6830_, new_n6831_, new_n6832_, new_n6833_, new_n6834_, new_n6835_,
    new_n6836_, new_n6837_, new_n6838_, new_n6839_, new_n6840_, new_n6841_,
    new_n6842_, new_n6843_, new_n6844_, new_n6845_, new_n6846_, new_n6847_,
    new_n6848_, new_n6849_, new_n6850_, new_n6851_, new_n6852_, new_n6853_,
    new_n6854_, new_n6855_, new_n6856_, new_n6857_, new_n6858_, new_n6859_,
    new_n6860_, new_n6861_, new_n6862_, new_n6863_, new_n6864_, new_n6865_,
    new_n6866_, new_n6867_, new_n6868_, new_n6869_, new_n6870_, new_n6871_,
    new_n6872_, new_n6873_, new_n6874_, new_n6875_, new_n6876_, new_n6877_,
    new_n6878_, new_n6879_, new_n6880_, new_n6881_, new_n6882_, new_n6883_,
    new_n6884_, new_n6885_, new_n6886_, new_n6887_, new_n6888_, new_n6889_,
    new_n6890_, new_n6891_, new_n6892_, new_n6893_, new_n6894_, new_n6895_,
    new_n6896_, new_n6897_, new_n6898_, new_n6899_, new_n6900_, new_n6901_,
    new_n6902_, new_n6903_, new_n6904_, new_n6905_, new_n6906_, new_n6907_,
    new_n6908_, new_n6909_, new_n6910_, new_n6911_, new_n6912_, new_n6913_,
    new_n6914_, new_n6915_, new_n6916_, new_n6917_, new_n6918_, new_n6919_,
    new_n6920_, new_n6921_, new_n6922_, new_n6923_, new_n6924_, new_n6925_,
    new_n6926_, new_n6927_, new_n6928_, new_n6929_, new_n6930_, new_n6931_,
    new_n6932_, new_n6933_, new_n6934_, new_n6935_, new_n6936_, new_n6937_,
    new_n6938_, new_n6939_, new_n6940_, new_n6941_, new_n6942_, new_n6943_,
    new_n6944_, new_n6945_, new_n6946_, new_n6947_, new_n6948_, new_n6949_,
    new_n6950_, new_n6951_, new_n6952_, new_n6953_, new_n6954_, new_n6955_,
    new_n6956_, new_n6957_, new_n6958_, new_n6959_, new_n6960_, new_n6961_,
    new_n6962_, new_n6963_, new_n6964_, new_n6965_, new_n6966_, new_n6967_,
    new_n6968_, new_n6969_, new_n6970_, new_n6971_, new_n6972_, new_n6973_,
    new_n6974_, new_n6975_, new_n6976_, new_n6977_, new_n6978_, new_n6979_,
    new_n6980_, new_n6981_, new_n6982_, new_n6983_, new_n6984_, new_n6985_,
    new_n6986_, new_n6987_, new_n6988_, new_n6989_, new_n6990_, new_n6991_,
    new_n6992_, new_n6993_, new_n6994_, new_n6995_, new_n6996_, new_n6997_,
    new_n6998_, new_n6999_, new_n7000_, new_n7001_, new_n7002_, new_n7003_,
    new_n7004_, new_n7005_, new_n7006_, new_n7007_, new_n7008_, new_n7009_,
    new_n7010_, new_n7011_, new_n7012_, new_n7013_, new_n7014_, new_n7015_,
    new_n7016_, new_n7017_, new_n7018_, new_n7019_, new_n7020_, new_n7021_,
    new_n7022_, new_n7023_, new_n7024_, new_n7025_, new_n7026_, new_n7027_,
    new_n7028_, new_n7029_, new_n7030_, new_n7031_, new_n7032_, new_n7033_,
    new_n7034_, new_n7035_, new_n7036_, new_n7037_, new_n7038_, new_n7039_,
    new_n7040_, new_n7041_, new_n7042_, new_n7043_, new_n7044_, new_n7045_,
    new_n7046_, new_n7047_, new_n7048_, new_n7049_, new_n7050_, new_n7051_,
    new_n7052_, new_n7053_, new_n7054_, new_n7055_, new_n7056_, new_n7057_,
    new_n7058_, new_n7059_, new_n7060_, new_n7061_, new_n7062_, new_n7063_,
    new_n7064_, new_n7065_, new_n7066_, new_n7067_, new_n7068_, new_n7069_,
    new_n7070_, new_n7071_, new_n7072_, new_n7073_, new_n7074_, new_n7075_,
    new_n7076_, new_n7077_, new_n7078_, new_n7079_, new_n7080_, new_n7081_,
    new_n7082_, new_n7083_, new_n7084_, new_n7085_, new_n7086_, new_n7087_,
    new_n7088_, new_n7089_, new_n7090_, new_n7091_, new_n7092_, new_n7093_,
    new_n7094_, new_n7095_, new_n7096_, new_n7097_, new_n7098_, new_n7099_,
    new_n7100_, new_n7101_, new_n7102_, new_n7103_, new_n7104_, new_n7105_,
    new_n7106_, new_n7107_, new_n7108_, new_n7109_, new_n7110_, new_n7111_,
    new_n7112_, new_n7113_, new_n7114_, new_n7115_, new_n7116_, new_n7117_,
    new_n7118_, new_n7119_, new_n7120_, new_n7121_, new_n7122_, new_n7123_,
    new_n7124_, new_n7125_, new_n7126_, new_n7127_, new_n7128_, new_n7129_,
    new_n7130_, new_n7131_, new_n7132_, new_n7133_, new_n7134_, new_n7135_,
    new_n7136_, new_n7137_, new_n7138_, new_n7139_, new_n7140_, new_n7141_,
    new_n7142_, new_n7143_, new_n7144_, new_n7145_, new_n7146_, new_n7147_,
    new_n7148_, new_n7149_, new_n7150_, new_n7151_, new_n7152_, new_n7153_,
    new_n7154_, new_n7155_, new_n7156_, new_n7157_, new_n7158_, new_n7159_,
    new_n7160_, new_n7161_, new_n7162_, new_n7164_, new_n7165_, new_n7166_,
    new_n7167_, new_n7168_, new_n7169_, new_n7170_, new_n7171_, new_n7172_,
    new_n7173_, new_n7174_, new_n7175_, new_n7176_, new_n7177_, new_n7178_,
    new_n7179_, new_n7180_, new_n7181_, new_n7182_, new_n7183_, new_n7184_,
    new_n7185_, new_n7186_, new_n7187_, new_n7188_, new_n7189_, new_n7190_,
    new_n7191_, new_n7192_, new_n7193_, new_n7194_, new_n7195_, new_n7196_,
    new_n7197_, new_n7198_, new_n7199_, new_n7200_, new_n7201_, new_n7202_,
    new_n7203_, new_n7204_, new_n7205_, new_n7206_, new_n7207_, new_n7208_,
    new_n7209_, new_n7210_, new_n7211_, new_n7212_, new_n7213_, new_n7214_,
    new_n7215_, new_n7216_, new_n7217_, new_n7218_, new_n7219_, new_n7220_,
    new_n7221_, new_n7222_, new_n7223_, new_n7224_, new_n7225_, new_n7226_,
    new_n7227_, new_n7228_, new_n7229_, new_n7230_, new_n7231_, new_n7232_,
    new_n7233_, new_n7234_, new_n7235_, new_n7236_, new_n7237_, new_n7238_,
    new_n7239_, new_n7240_, new_n7241_, new_n7242_, new_n7243_, new_n7244_,
    new_n7245_, new_n7246_, new_n7247_, new_n7248_, new_n7249_, new_n7250_,
    new_n7251_, new_n7252_, new_n7253_, new_n7254_, new_n7255_, new_n7256_,
    new_n7257_, new_n7258_, new_n7259_, new_n7260_, new_n7261_, new_n7262_,
    new_n7263_, new_n7264_, new_n7265_, new_n7266_, new_n7267_, new_n7268_,
    new_n7269_, new_n7270_, new_n7271_, new_n7272_, new_n7273_, new_n7274_,
    new_n7275_, new_n7276_, new_n7277_, new_n7278_, new_n7279_, new_n7280_,
    new_n7281_, new_n7282_, new_n7283_, new_n7284_, new_n7285_, new_n7286_,
    new_n7287_, new_n7288_, new_n7289_, new_n7290_, new_n7291_, new_n7292_,
    new_n7293_, new_n7294_, new_n7295_, new_n7296_, new_n7297_, new_n7298_,
    new_n7299_, new_n7300_, new_n7301_, new_n7302_, new_n7303_, new_n7304_,
    new_n7305_, new_n7306_, new_n7307_, new_n7308_, new_n7309_, new_n7310_,
    new_n7311_, new_n7312_, new_n7313_, new_n7314_, new_n7315_, new_n7316_,
    new_n7317_, new_n7318_, new_n7319_, new_n7320_, new_n7321_, new_n7322_,
    new_n7323_, new_n7324_, new_n7325_, new_n7326_, new_n7327_, new_n7328_,
    new_n7329_, new_n7330_, new_n7331_, new_n7332_, new_n7333_, new_n7334_,
    new_n7335_, new_n7336_, new_n7337_, new_n7338_, new_n7339_, new_n7340_,
    new_n7341_, new_n7342_, new_n7343_, new_n7344_, new_n7345_, new_n7346_,
    new_n7347_, new_n7348_, new_n7349_, new_n7350_, new_n7351_, new_n7352_,
    new_n7353_, new_n7354_, new_n7355_, new_n7356_, new_n7357_, new_n7358_,
    new_n7359_, new_n7360_, new_n7361_, new_n7362_, new_n7363_, new_n7364_,
    new_n7365_, new_n7366_, new_n7367_, new_n7368_, new_n7369_, new_n7370_,
    new_n7371_, new_n7372_, new_n7373_, new_n7374_, new_n7375_, new_n7376_,
    new_n7377_, new_n7378_, new_n7379_, new_n7380_, new_n7381_, new_n7382_,
    new_n7383_, new_n7384_, new_n7385_, new_n7386_, new_n7387_, new_n7388_,
    new_n7389_, new_n7390_, new_n7391_, new_n7392_, new_n7393_, new_n7394_,
    new_n7395_, new_n7396_, new_n7397_, new_n7398_, new_n7399_, new_n7400_,
    new_n7401_, new_n7402_, new_n7403_, new_n7404_, new_n7405_, new_n7406_,
    new_n7407_, new_n7408_, new_n7409_, new_n7410_, new_n7411_, new_n7412_,
    new_n7413_, new_n7414_, new_n7415_, new_n7416_, new_n7417_, new_n7418_,
    new_n7419_, new_n7420_, new_n7421_, new_n7422_, new_n7423_, new_n7424_,
    new_n7425_, new_n7426_, new_n7427_, new_n7428_, new_n7429_, new_n7430_,
    new_n7431_, new_n7432_, new_n7433_, new_n7434_, new_n7435_, new_n7436_,
    new_n7437_, new_n7438_, new_n7439_, new_n7440_, new_n7441_, new_n7442_,
    new_n7443_, new_n7444_, new_n7445_, new_n7446_, new_n7447_, new_n7448_,
    new_n7449_, new_n7450_, new_n7451_, new_n7452_, new_n7453_, new_n7454_,
    new_n7455_, new_n7456_, new_n7457_, new_n7458_, new_n7459_, new_n7460_,
    new_n7461_, new_n7462_, new_n7463_, new_n7464_, new_n7465_, new_n7466_,
    new_n7467_, new_n7468_, new_n7469_, new_n7470_, new_n7471_, new_n7472_,
    new_n7473_, new_n7474_, new_n7475_, new_n7476_, new_n7477_, new_n7478_,
    new_n7479_, new_n7480_, new_n7481_, new_n7482_, new_n7483_, new_n7484_,
    new_n7485_, new_n7486_, new_n7487_, new_n7488_, new_n7489_, new_n7490_,
    new_n7491_, new_n7492_, new_n7493_, new_n7494_, new_n7495_, new_n7496_,
    new_n7497_, new_n7498_, new_n7499_, new_n7500_, new_n7501_, new_n7502_,
    new_n7503_, new_n7504_, new_n7505_, new_n7506_, new_n7507_, new_n7508_,
    new_n7509_, new_n7510_, new_n7511_, new_n7512_, new_n7513_, new_n7514_,
    new_n7515_, new_n7516_, new_n7517_, new_n7518_, new_n7519_, new_n7520_,
    new_n7521_, new_n7522_, new_n7523_, new_n7524_, new_n7525_, new_n7526_,
    new_n7527_, new_n7528_, new_n7529_, new_n7530_, new_n7531_, new_n7532_,
    new_n7533_, new_n7534_, new_n7535_, new_n7536_, new_n7537_, new_n7538_,
    new_n7539_, new_n7540_, new_n7541_, new_n7542_, new_n7543_, new_n7544_,
    new_n7545_, new_n7546_, new_n7547_, new_n7548_, new_n7549_, new_n7550_,
    new_n7551_, new_n7552_, new_n7553_, new_n7554_, new_n7555_, new_n7556_,
    new_n7557_, new_n7558_, new_n7559_, new_n7560_, new_n7561_, new_n7562_,
    new_n7563_, new_n7564_, new_n7565_, new_n7566_, new_n7567_, new_n7568_,
    new_n7569_, new_n7570_, new_n7571_, new_n7572_, new_n7573_, new_n7574_,
    new_n7575_, new_n7576_, new_n7577_, new_n7578_, new_n7579_, new_n7580_,
    new_n7581_, new_n7582_, new_n7583_, new_n7584_, new_n7585_, new_n7586_,
    new_n7587_, new_n7588_, new_n7589_, new_n7590_, new_n7591_, new_n7592_,
    new_n7593_, new_n7594_, new_n7595_, new_n7596_, new_n7597_, new_n7598_,
    new_n7599_, new_n7600_, new_n7601_, new_n7603_, new_n7604_, new_n7605_,
    new_n7606_, new_n7607_, new_n7608_, new_n7609_, new_n7610_, new_n7611_,
    new_n7612_, new_n7613_, new_n7614_, new_n7615_, new_n7616_, new_n7617_,
    new_n7618_, new_n7619_, new_n7620_, new_n7621_, new_n7622_, new_n7623_,
    new_n7624_, new_n7625_, new_n7626_, new_n7627_, new_n7628_, new_n7629_,
    new_n7630_, new_n7631_, new_n7632_, new_n7633_, new_n7634_, new_n7635_,
    new_n7636_, new_n7637_, new_n7638_, new_n7639_, new_n7640_, new_n7641_,
    new_n7642_, new_n7643_, new_n7644_, new_n7645_, new_n7646_, new_n7647_,
    new_n7648_, new_n7649_, new_n7650_, new_n7651_, new_n7652_, new_n7653_,
    new_n7654_, new_n7655_, new_n7656_, new_n7657_, new_n7658_, new_n7659_,
    new_n7660_, new_n7661_, new_n7662_, new_n7663_, new_n7664_, new_n7665_,
    new_n7666_, new_n7667_, new_n7668_, new_n7669_, new_n7670_, new_n7671_,
    new_n7672_, new_n7673_, new_n7674_, new_n7675_, new_n7676_, new_n7677_,
    new_n7678_, new_n7679_, new_n7680_, new_n7681_, new_n7682_, new_n7683_,
    new_n7684_, new_n7685_, new_n7686_, new_n7687_, new_n7688_, new_n7689_,
    new_n7690_, new_n7691_, new_n7692_, new_n7693_, new_n7694_, new_n7695_,
    new_n7696_, new_n7697_, new_n7698_, new_n7699_, new_n7700_, new_n7701_,
    new_n7702_, new_n7703_, new_n7704_, new_n7705_, new_n7706_, new_n7707_,
    new_n7708_, new_n7709_, new_n7710_, new_n7711_, new_n7712_, new_n7713_,
    new_n7714_, new_n7715_, new_n7716_, new_n7717_, new_n7718_, new_n7719_,
    new_n7720_, new_n7721_, new_n7722_, new_n7723_, new_n7724_, new_n7725_,
    new_n7726_, new_n7727_, new_n7728_, new_n7729_, new_n7730_, new_n7731_,
    new_n7732_, new_n7733_, new_n7734_, new_n7735_, new_n7736_, new_n7737_,
    new_n7738_, new_n7739_, new_n7740_, new_n7741_, new_n7742_, new_n7743_,
    new_n7744_, new_n7745_, new_n7746_, new_n7747_, new_n7748_, new_n7749_,
    new_n7750_, new_n7751_, new_n7752_, new_n7753_, new_n7754_, new_n7755_,
    new_n7756_, new_n7757_, new_n7758_, new_n7759_, new_n7760_, new_n7761_,
    new_n7762_, new_n7763_, new_n7764_, new_n7765_, new_n7766_, new_n7767_,
    new_n7768_, new_n7769_, new_n7770_, new_n7771_, new_n7772_, new_n7773_,
    new_n7774_, new_n7775_, new_n7776_, new_n7777_, new_n7778_, new_n7779_,
    new_n7780_, new_n7781_, new_n7782_, new_n7783_, new_n7784_, new_n7785_,
    new_n7786_, new_n7787_, new_n7788_, new_n7789_, new_n7790_, new_n7791_,
    new_n7792_, new_n7793_, new_n7794_, new_n7795_, new_n7796_, new_n7797_,
    new_n7798_, new_n7799_, new_n7800_, new_n7801_, new_n7802_, new_n7803_,
    new_n7804_, new_n7805_, new_n7806_, new_n7807_, new_n7808_, new_n7809_,
    new_n7810_, new_n7811_, new_n7812_, new_n7813_, new_n7814_, new_n7815_,
    new_n7816_, new_n7817_, new_n7818_, new_n7819_, new_n7820_, new_n7821_,
    new_n7822_, new_n7823_, new_n7824_, new_n7825_, new_n7826_, new_n7827_,
    new_n7828_, new_n7829_, new_n7830_, new_n7831_, new_n7832_, new_n7833_,
    new_n7834_, new_n7835_, new_n7836_, new_n7837_, new_n7838_, new_n7839_,
    new_n7840_, new_n7841_, new_n7842_, new_n7843_, new_n7844_, new_n7845_,
    new_n7846_, new_n7847_, new_n7848_, new_n7849_, new_n7850_, new_n7851_,
    new_n7852_, new_n7853_, new_n7854_, new_n7855_, new_n7856_, new_n7857_,
    new_n7858_, new_n7859_, new_n7860_, new_n7861_, new_n7862_, new_n7863_,
    new_n7864_, new_n7865_, new_n7866_, new_n7867_, new_n7868_, new_n7869_,
    new_n7870_, new_n7871_, new_n7872_, new_n7873_, new_n7874_, new_n7875_,
    new_n7876_, new_n7877_, new_n7878_, new_n7879_, new_n7880_, new_n7881_,
    new_n7882_, new_n7883_, new_n7884_, new_n7885_, new_n7886_, new_n7887_,
    new_n7888_, new_n7889_, new_n7890_, new_n7891_, new_n7892_, new_n7893_,
    new_n7894_, new_n7895_, new_n7896_, new_n7897_, new_n7898_, new_n7899_,
    new_n7900_, new_n7901_, new_n7902_, new_n7903_, new_n7904_, new_n7905_,
    new_n7906_, new_n7907_, new_n7908_, new_n7909_, new_n7910_, new_n7911_,
    new_n7912_, new_n7913_, new_n7914_, new_n7915_, new_n7916_, new_n7917_,
    new_n7918_, new_n7919_, new_n7920_, new_n7921_, new_n7922_, new_n7923_,
    new_n7924_, new_n7925_, new_n7926_, new_n7927_, new_n7928_, new_n7929_,
    new_n7930_, new_n7931_, new_n7932_, new_n7933_, new_n7934_, new_n7935_,
    new_n7936_, new_n7937_, new_n7938_, new_n7939_, new_n7940_, new_n7941_,
    new_n7942_, new_n7943_, new_n7944_, new_n7945_, new_n7946_, new_n7947_,
    new_n7948_, new_n7949_, new_n7950_, new_n7951_, new_n7952_, new_n7953_,
    new_n7954_, new_n7955_, new_n7956_, new_n7957_, new_n7958_, new_n7959_,
    new_n7960_, new_n7961_, new_n7962_, new_n7963_, new_n7964_, new_n7965_,
    new_n7966_, new_n7967_, new_n7968_, new_n7969_, new_n7970_, new_n7971_,
    new_n7972_, new_n7973_, new_n7974_, new_n7975_, new_n7976_, new_n7977_,
    new_n7978_, new_n7979_, new_n7980_, new_n7981_, new_n7982_, new_n7983_,
    new_n7984_, new_n7985_, new_n7986_, new_n7987_, new_n7988_, new_n7989_,
    new_n7990_, new_n7991_, new_n7992_, new_n7993_, new_n7994_, new_n7995_,
    new_n7996_, new_n7997_, new_n7998_, new_n7999_, new_n8000_, new_n8001_,
    new_n8002_, new_n8003_, new_n8004_, new_n8005_, new_n8006_, new_n8007_,
    new_n8008_, new_n8009_, new_n8010_, new_n8011_, new_n8012_, new_n8013_,
    new_n8014_, new_n8015_, new_n8016_, new_n8017_, new_n8018_, new_n8019_,
    new_n8020_, new_n8021_, new_n8022_, new_n8023_, new_n8024_, new_n8025_,
    new_n8026_, new_n8027_, new_n8028_, new_n8029_, new_n8030_, new_n8031_,
    new_n8032_, new_n8033_, new_n8034_, new_n8035_, new_n8036_, new_n8037_,
    new_n8038_, new_n8039_, new_n8040_, new_n8041_, new_n8042_, new_n8043_,
    new_n8044_, new_n8045_, new_n8046_, new_n8047_, new_n8048_, new_n8049_,
    new_n8050_, new_n8051_, new_n8052_, new_n8053_, new_n8054_, new_n8056_,
    new_n8057_, new_n8058_, new_n8059_, new_n8060_, new_n8061_, new_n8062_,
    new_n8063_, new_n8064_, new_n8065_, new_n8066_, new_n8067_, new_n8068_,
    new_n8069_, new_n8070_, new_n8071_, new_n8072_, new_n8073_, new_n8074_,
    new_n8075_, new_n8076_, new_n8077_, new_n8078_, new_n8079_, new_n8080_,
    new_n8081_, new_n8082_, new_n8083_, new_n8084_, new_n8085_, new_n8086_,
    new_n8087_, new_n8088_, new_n8089_, new_n8090_, new_n8091_, new_n8092_,
    new_n8093_, new_n8094_, new_n8095_, new_n8096_, new_n8097_, new_n8098_,
    new_n8099_, new_n8100_, new_n8101_, new_n8102_, new_n8103_, new_n8104_,
    new_n8105_, new_n8106_, new_n8107_, new_n8108_, new_n8109_, new_n8110_,
    new_n8111_, new_n8112_, new_n8113_, new_n8114_, new_n8115_, new_n8116_,
    new_n8117_, new_n8118_, new_n8119_, new_n8120_, new_n8121_, new_n8122_,
    new_n8123_, new_n8124_, new_n8125_, new_n8126_, new_n8127_, new_n8128_,
    new_n8129_, new_n8130_, new_n8131_, new_n8132_, new_n8133_, new_n8134_,
    new_n8135_, new_n8136_, new_n8137_, new_n8138_, new_n8139_, new_n8140_,
    new_n8141_, new_n8142_, new_n8143_, new_n8144_, new_n8145_, new_n8146_,
    new_n8147_, new_n8148_, new_n8149_, new_n8150_, new_n8151_, new_n8152_,
    new_n8153_, new_n8154_, new_n8155_, new_n8156_, new_n8157_, new_n8158_,
    new_n8159_, new_n8160_, new_n8161_, new_n8162_, new_n8163_, new_n8164_,
    new_n8165_, new_n8166_, new_n8167_, new_n8168_, new_n8169_, new_n8170_,
    new_n8171_, new_n8172_, new_n8173_, new_n8174_, new_n8175_, new_n8176_,
    new_n8177_, new_n8178_, new_n8179_, new_n8180_, new_n8181_, new_n8182_,
    new_n8183_, new_n8184_, new_n8185_, new_n8186_, new_n8187_, new_n8188_,
    new_n8189_, new_n8190_, new_n8191_, new_n8192_, new_n8193_, new_n8194_,
    new_n8195_, new_n8196_, new_n8197_, new_n8198_, new_n8199_, new_n8200_,
    new_n8201_, new_n8202_, new_n8203_, new_n8204_, new_n8205_, new_n8206_,
    new_n8207_, new_n8208_, new_n8209_, new_n8210_, new_n8211_, new_n8212_,
    new_n8213_, new_n8214_, new_n8215_, new_n8216_, new_n8217_, new_n8218_,
    new_n8219_, new_n8220_, new_n8221_, new_n8222_, new_n8223_, new_n8224_,
    new_n8225_, new_n8226_, new_n8227_, new_n8228_, new_n8229_, new_n8230_,
    new_n8231_, new_n8232_, new_n8233_, new_n8234_, new_n8235_, new_n8236_,
    new_n8237_, new_n8238_, new_n8239_, new_n8240_, new_n8241_, new_n8242_,
    new_n8243_, new_n8244_, new_n8245_, new_n8246_, new_n8247_, new_n8248_,
    new_n8249_, new_n8250_, new_n8251_, new_n8252_, new_n8253_, new_n8254_,
    new_n8255_, new_n8256_, new_n8257_, new_n8258_, new_n8259_, new_n8260_,
    new_n8261_, new_n8262_, new_n8263_, new_n8264_, new_n8265_, new_n8266_,
    new_n8267_, new_n8268_, new_n8269_, new_n8270_, new_n8271_, new_n8272_,
    new_n8273_, new_n8274_, new_n8275_, new_n8276_, new_n8277_, new_n8278_,
    new_n8279_, new_n8280_, new_n8281_, new_n8282_, new_n8283_, new_n8284_,
    new_n8285_, new_n8286_, new_n8287_, new_n8288_, new_n8289_, new_n8290_,
    new_n8291_, new_n8292_, new_n8293_, new_n8294_, new_n8295_, new_n8296_,
    new_n8297_, new_n8298_, new_n8299_, new_n8300_, new_n8301_, new_n8302_,
    new_n8303_, new_n8304_, new_n8305_, new_n8306_, new_n8307_, new_n8308_,
    new_n8309_, new_n8310_, new_n8311_, new_n8312_, new_n8313_, new_n8314_,
    new_n8315_, new_n8316_, new_n8317_, new_n8318_, new_n8319_, new_n8320_,
    new_n8321_, new_n8322_, new_n8323_, new_n8324_, new_n8325_, new_n8326_,
    new_n8327_, new_n8328_, new_n8329_, new_n8330_, new_n8331_, new_n8332_,
    new_n8333_, new_n8334_, new_n8335_, new_n8336_, new_n8337_, new_n8338_,
    new_n8339_, new_n8340_, new_n8341_, new_n8342_, new_n8343_, new_n8344_,
    new_n8345_, new_n8346_, new_n8347_, new_n8348_, new_n8349_, new_n8350_,
    new_n8351_, new_n8352_, new_n8353_, new_n8354_, new_n8355_, new_n8356_,
    new_n8357_, new_n8358_, new_n8359_, new_n8360_, new_n8361_, new_n8362_,
    new_n8363_, new_n8364_, new_n8365_, new_n8366_, new_n8367_, new_n8368_,
    new_n8369_, new_n8370_, new_n8371_, new_n8372_, new_n8373_, new_n8374_,
    new_n8375_, new_n8376_, new_n8377_, new_n8378_, new_n8379_, new_n8380_,
    new_n8381_, new_n8382_, new_n8383_, new_n8384_, new_n8385_, new_n8386_,
    new_n8387_, new_n8388_, new_n8389_, new_n8390_, new_n8391_, new_n8392_,
    new_n8393_, new_n8394_, new_n8395_, new_n8396_, new_n8397_, new_n8398_,
    new_n8399_, new_n8400_, new_n8401_, new_n8402_, new_n8403_, new_n8404_,
    new_n8405_, new_n8406_, new_n8407_, new_n8408_, new_n8409_, new_n8410_,
    new_n8411_, new_n8412_, new_n8413_, new_n8414_, new_n8415_, new_n8416_,
    new_n8417_, new_n8418_, new_n8419_, new_n8420_, new_n8421_, new_n8422_,
    new_n8423_, new_n8424_, new_n8425_, new_n8426_, new_n8427_, new_n8428_,
    new_n8429_, new_n8430_, new_n8431_, new_n8432_, new_n8433_, new_n8434_,
    new_n8435_, new_n8436_, new_n8437_, new_n8438_, new_n8439_, new_n8440_,
    new_n8441_, new_n8442_, new_n8443_, new_n8444_, new_n8445_, new_n8446_,
    new_n8447_, new_n8448_, new_n8449_, new_n8450_, new_n8451_, new_n8452_,
    new_n8453_, new_n8454_, new_n8455_, new_n8456_, new_n8457_, new_n8458_,
    new_n8459_, new_n8460_, new_n8461_, new_n8462_, new_n8463_, new_n8464_,
    new_n8465_, new_n8466_, new_n8467_, new_n8468_, new_n8469_, new_n8470_,
    new_n8471_, new_n8472_, new_n8473_, new_n8474_, new_n8475_, new_n8476_,
    new_n8477_, new_n8478_, new_n8479_, new_n8480_, new_n8481_, new_n8482_,
    new_n8483_, new_n8484_, new_n8485_, new_n8486_, new_n8487_, new_n8488_,
    new_n8489_, new_n8490_, new_n8491_, new_n8492_, new_n8493_, new_n8494_,
    new_n8495_, new_n8496_, new_n8497_, new_n8498_, new_n8499_, new_n8500_,
    new_n8501_, new_n8502_, new_n8503_, new_n8504_, new_n8505_, new_n8506_,
    new_n8507_, new_n8508_, new_n8509_, new_n8510_, new_n8511_, new_n8512_,
    new_n8513_, new_n8514_, new_n8515_, new_n8516_, new_n8517_, new_n8518_,
    new_n8519_, new_n8521_, new_n8522_, new_n8523_, new_n8524_, new_n8525_,
    new_n8526_, new_n8527_, new_n8528_, new_n8529_, new_n8530_, new_n8531_,
    new_n8532_, new_n8533_, new_n8534_, new_n8535_, new_n8536_, new_n8537_,
    new_n8538_, new_n8539_, new_n8540_, new_n8541_, new_n8542_, new_n8543_,
    new_n8544_, new_n8545_, new_n8546_, new_n8547_, new_n8548_, new_n8549_,
    new_n8550_, new_n8551_, new_n8552_, new_n8553_, new_n8554_, new_n8555_,
    new_n8556_, new_n8557_, new_n8558_, new_n8559_, new_n8560_, new_n8561_,
    new_n8562_, new_n8563_, new_n8564_, new_n8565_, new_n8566_, new_n8567_,
    new_n8568_, new_n8569_, new_n8570_, new_n8571_, new_n8572_, new_n8573_,
    new_n8574_, new_n8575_, new_n8576_, new_n8577_, new_n8578_, new_n8579_,
    new_n8580_, new_n8581_, new_n8582_, new_n8583_, new_n8584_, new_n8585_,
    new_n8586_, new_n8587_, new_n8588_, new_n8589_, new_n8590_, new_n8591_,
    new_n8592_, new_n8593_, new_n8594_, new_n8595_, new_n8596_, new_n8597_,
    new_n8598_, new_n8599_, new_n8600_, new_n8601_, new_n8602_, new_n8603_,
    new_n8604_, new_n8605_, new_n8606_, new_n8607_, new_n8608_, new_n8609_,
    new_n8610_, new_n8611_, new_n8612_, new_n8613_, new_n8614_, new_n8615_,
    new_n8616_, new_n8617_, new_n8618_, new_n8619_, new_n8620_, new_n8621_,
    new_n8622_, new_n8623_, new_n8624_, new_n8625_, new_n8626_, new_n8627_,
    new_n8628_, new_n8629_, new_n8630_, new_n8631_, new_n8632_, new_n8633_,
    new_n8634_, new_n8635_, new_n8636_, new_n8637_, new_n8638_, new_n8639_,
    new_n8640_, new_n8641_, new_n8642_, new_n8643_, new_n8644_, new_n8645_,
    new_n8646_, new_n8647_, new_n8648_, new_n8649_, new_n8650_, new_n8651_,
    new_n8652_, new_n8653_, new_n8654_, new_n8655_, new_n8656_, new_n8657_,
    new_n8658_, new_n8659_, new_n8660_, new_n8661_, new_n8662_, new_n8663_,
    new_n8664_, new_n8665_, new_n8666_, new_n8667_, new_n8668_, new_n8669_,
    new_n8670_, new_n8671_, new_n8672_, new_n8673_, new_n8674_, new_n8675_,
    new_n8676_, new_n8677_, new_n8678_, new_n8679_, new_n8680_, new_n8681_,
    new_n8682_, new_n8683_, new_n8684_, new_n8685_, new_n8686_, new_n8687_,
    new_n8688_, new_n8689_, new_n8690_, new_n8691_, new_n8692_, new_n8693_,
    new_n8694_, new_n8695_, new_n8696_, new_n8697_, new_n8698_, new_n8699_,
    new_n8700_, new_n8701_, new_n8702_, new_n8703_, new_n8704_, new_n8705_,
    new_n8706_, new_n8707_, new_n8708_, new_n8709_, new_n8710_, new_n8711_,
    new_n8712_, new_n8713_, new_n8714_, new_n8715_, new_n8716_, new_n8717_,
    new_n8718_, new_n8719_, new_n8720_, new_n8721_, new_n8722_, new_n8723_,
    new_n8724_, new_n8725_, new_n8726_, new_n8727_, new_n8728_, new_n8729_,
    new_n8730_, new_n8731_, new_n8732_, new_n8733_, new_n8734_, new_n8735_,
    new_n8736_, new_n8737_, new_n8738_, new_n8739_, new_n8740_, new_n8741_,
    new_n8742_, new_n8743_, new_n8744_, new_n8745_, new_n8746_, new_n8747_,
    new_n8748_, new_n8749_, new_n8750_, new_n8751_, new_n8752_, new_n8753_,
    new_n8754_, new_n8755_, new_n8756_, new_n8757_, new_n8758_, new_n8759_,
    new_n8760_, new_n8761_, new_n8762_, new_n8763_, new_n8764_, new_n8765_,
    new_n8766_, new_n8767_, new_n8768_, new_n8769_, new_n8770_, new_n8771_,
    new_n8772_, new_n8773_, new_n8774_, new_n8775_, new_n8776_, new_n8777_,
    new_n8778_, new_n8779_, new_n8780_, new_n8781_, new_n8782_, new_n8783_,
    new_n8784_, new_n8785_, new_n8786_, new_n8787_, new_n8788_, new_n8789_,
    new_n8790_, new_n8791_, new_n8792_, new_n8793_, new_n8794_, new_n8795_,
    new_n8796_, new_n8797_, new_n8798_, new_n8799_, new_n8800_, new_n8801_,
    new_n8802_, new_n8803_, new_n8804_, new_n8805_, new_n8806_, new_n8807_,
    new_n8808_, new_n8809_, new_n8810_, new_n8811_, new_n8812_, new_n8813_,
    new_n8814_, new_n8815_, new_n8816_, new_n8817_, new_n8818_, new_n8819_,
    new_n8820_, new_n8821_, new_n8822_, new_n8823_, new_n8824_, new_n8825_,
    new_n8826_, new_n8827_, new_n8828_, new_n8829_, new_n8830_, new_n8831_,
    new_n8832_, new_n8833_, new_n8834_, new_n8835_, new_n8836_, new_n8837_,
    new_n8838_, new_n8839_, new_n8840_, new_n8841_, new_n8842_, new_n8843_,
    new_n8844_, new_n8845_, new_n8846_, new_n8847_, new_n8848_, new_n8849_,
    new_n8850_, new_n8851_, new_n8852_, new_n8853_, new_n8854_, new_n8855_,
    new_n8856_, new_n8857_, new_n8858_, new_n8859_, new_n8860_, new_n8861_,
    new_n8862_, new_n8863_, new_n8864_, new_n8865_, new_n8866_, new_n8867_,
    new_n8868_, new_n8869_, new_n8870_, new_n8871_, new_n8872_, new_n8873_,
    new_n8874_, new_n8875_, new_n8876_, new_n8877_, new_n8878_, new_n8879_,
    new_n8880_, new_n8881_, new_n8882_, new_n8883_, new_n8884_, new_n8885_,
    new_n8886_, new_n8887_, new_n8888_, new_n8889_, new_n8890_, new_n8891_,
    new_n8892_, new_n8893_, new_n8894_, new_n8895_, new_n8896_, new_n8897_,
    new_n8898_, new_n8899_, new_n8900_, new_n8901_, new_n8902_, new_n8903_,
    new_n8904_, new_n8905_, new_n8906_, new_n8907_, new_n8908_, new_n8909_,
    new_n8910_, new_n8911_, new_n8912_, new_n8913_, new_n8914_, new_n8915_,
    new_n8916_, new_n8917_, new_n8918_, new_n8919_, new_n8920_, new_n8921_,
    new_n8922_, new_n8923_, new_n8924_, new_n8925_, new_n8926_, new_n8927_,
    new_n8928_, new_n8929_, new_n8930_, new_n8931_, new_n8932_, new_n8933_,
    new_n8934_, new_n8935_, new_n8936_, new_n8937_, new_n8938_, new_n8939_,
    new_n8940_, new_n8941_, new_n8942_, new_n8943_, new_n8944_, new_n8945_,
    new_n8946_, new_n8947_, new_n8948_, new_n8949_, new_n8950_, new_n8951_,
    new_n8952_, new_n8953_, new_n8954_, new_n8955_, new_n8956_, new_n8957_,
    new_n8958_, new_n8959_, new_n8960_, new_n8961_, new_n8962_, new_n8963_,
    new_n8964_, new_n8965_, new_n8966_, new_n8967_, new_n8968_, new_n8969_,
    new_n8970_, new_n8971_, new_n8972_, new_n8973_, new_n8974_, new_n8975_,
    new_n8976_, new_n8977_, new_n8978_, new_n8979_, new_n8980_, new_n8981_,
    new_n8982_, new_n8983_, new_n8984_, new_n8985_, new_n8986_, new_n8987_,
    new_n8988_, new_n8989_, new_n8990_, new_n8991_, new_n8992_, new_n8993_,
    new_n8994_, new_n8995_, new_n8996_, new_n8997_, new_n8998_, new_n8999_,
    new_n9000_, new_n9001_, new_n9002_, new_n9003_, new_n9004_, new_n9006_,
    new_n9007_, new_n9008_, new_n9009_, new_n9010_, new_n9011_, new_n9012_,
    new_n9013_, new_n9014_, new_n9015_, new_n9016_, new_n9017_, new_n9018_,
    new_n9019_, new_n9020_, new_n9021_, new_n9022_, new_n9023_, new_n9024_,
    new_n9025_, new_n9026_, new_n9027_, new_n9028_, new_n9029_, new_n9030_,
    new_n9031_, new_n9032_, new_n9033_, new_n9034_, new_n9035_, new_n9036_,
    new_n9037_, new_n9038_, new_n9039_, new_n9040_, new_n9041_, new_n9042_,
    new_n9043_, new_n9044_, new_n9045_, new_n9046_, new_n9047_, new_n9048_,
    new_n9049_, new_n9050_, new_n9051_, new_n9052_, new_n9053_, new_n9054_,
    new_n9055_, new_n9056_, new_n9057_, new_n9058_, new_n9059_, new_n9060_,
    new_n9061_, new_n9062_, new_n9063_, new_n9064_, new_n9065_, new_n9066_,
    new_n9067_, new_n9068_, new_n9069_, new_n9070_, new_n9071_, new_n9072_,
    new_n9073_, new_n9074_, new_n9075_, new_n9076_, new_n9077_, new_n9078_,
    new_n9079_, new_n9080_, new_n9081_, new_n9082_, new_n9083_, new_n9084_,
    new_n9085_, new_n9086_, new_n9087_, new_n9088_, new_n9089_, new_n9090_,
    new_n9091_, new_n9092_, new_n9093_, new_n9094_, new_n9095_, new_n9096_,
    new_n9097_, new_n9098_, new_n9099_, new_n9100_, new_n9101_, new_n9102_,
    new_n9103_, new_n9104_, new_n9105_, new_n9106_, new_n9107_, new_n9108_,
    new_n9109_, new_n9110_, new_n9111_, new_n9112_, new_n9113_, new_n9114_,
    new_n9115_, new_n9116_, new_n9117_, new_n9118_, new_n9119_, new_n9120_,
    new_n9121_, new_n9122_, new_n9123_, new_n9124_, new_n9125_, new_n9126_,
    new_n9127_, new_n9128_, new_n9129_, new_n9130_, new_n9131_, new_n9132_,
    new_n9133_, new_n9134_, new_n9135_, new_n9136_, new_n9137_, new_n9138_,
    new_n9139_, new_n9140_, new_n9141_, new_n9142_, new_n9143_, new_n9144_,
    new_n9145_, new_n9146_, new_n9147_, new_n9148_, new_n9149_, new_n9150_,
    new_n9151_, new_n9152_, new_n9153_, new_n9154_, new_n9155_, new_n9156_,
    new_n9157_, new_n9158_, new_n9159_, new_n9160_, new_n9161_, new_n9162_,
    new_n9163_, new_n9164_, new_n9165_, new_n9166_, new_n9167_, new_n9168_,
    new_n9169_, new_n9170_, new_n9171_, new_n9172_, new_n9173_, new_n9174_,
    new_n9175_, new_n9176_, new_n9177_, new_n9178_, new_n9179_, new_n9180_,
    new_n9181_, new_n9182_, new_n9183_, new_n9184_, new_n9185_, new_n9186_,
    new_n9187_, new_n9188_, new_n9189_, new_n9190_, new_n9191_, new_n9192_,
    new_n9193_, new_n9194_, new_n9195_, new_n9196_, new_n9197_, new_n9198_,
    new_n9199_, new_n9200_, new_n9201_, new_n9202_, new_n9203_, new_n9204_,
    new_n9205_, new_n9206_, new_n9207_, new_n9208_, new_n9209_, new_n9210_,
    new_n9211_, new_n9212_, new_n9213_, new_n9214_, new_n9215_, new_n9216_,
    new_n9217_, new_n9218_, new_n9219_, new_n9220_, new_n9221_, new_n9222_,
    new_n9223_, new_n9224_, new_n9225_, new_n9226_, new_n9227_, new_n9228_,
    new_n9229_, new_n9230_, new_n9231_, new_n9232_, new_n9233_, new_n9234_,
    new_n9235_, new_n9236_, new_n9237_, new_n9238_, new_n9239_, new_n9240_,
    new_n9241_, new_n9242_, new_n9243_, new_n9244_, new_n9245_, new_n9246_,
    new_n9247_, new_n9248_, new_n9249_, new_n9250_, new_n9251_, new_n9252_,
    new_n9253_, new_n9254_, new_n9255_, new_n9256_, new_n9257_, new_n9258_,
    new_n9259_, new_n9260_, new_n9261_, new_n9262_, new_n9263_, new_n9264_,
    new_n9265_, new_n9266_, new_n9267_, new_n9268_, new_n9269_, new_n9270_,
    new_n9271_, new_n9272_, new_n9273_, new_n9274_, new_n9275_, new_n9276_,
    new_n9277_, new_n9278_, new_n9279_, new_n9280_, new_n9281_, new_n9282_,
    new_n9283_, new_n9284_, new_n9285_, new_n9286_, new_n9287_, new_n9288_,
    new_n9289_, new_n9290_, new_n9291_, new_n9292_, new_n9293_, new_n9294_,
    new_n9295_, new_n9296_, new_n9297_, new_n9298_, new_n9299_, new_n9300_,
    new_n9301_, new_n9302_, new_n9303_, new_n9304_, new_n9305_, new_n9306_,
    new_n9307_, new_n9308_, new_n9309_, new_n9310_, new_n9311_, new_n9312_,
    new_n9313_, new_n9314_, new_n9315_, new_n9316_, new_n9317_, new_n9318_,
    new_n9319_, new_n9320_, new_n9321_, new_n9322_, new_n9323_, new_n9324_,
    new_n9325_, new_n9326_, new_n9327_, new_n9328_, new_n9329_, new_n9330_,
    new_n9331_, new_n9332_, new_n9333_, new_n9334_, new_n9335_, new_n9336_,
    new_n9337_, new_n9338_, new_n9339_, new_n9340_, new_n9341_, new_n9342_,
    new_n9343_, new_n9344_, new_n9345_, new_n9346_, new_n9347_, new_n9348_,
    new_n9349_, new_n9350_, new_n9351_, new_n9352_, new_n9353_, new_n9354_,
    new_n9355_, new_n9356_, new_n9357_, new_n9358_, new_n9359_, new_n9360_,
    new_n9361_, new_n9362_, new_n9363_, new_n9364_, new_n9365_, new_n9366_,
    new_n9367_, new_n9368_, new_n9369_, new_n9370_, new_n9371_, new_n9372_,
    new_n9373_, new_n9374_, new_n9375_, new_n9376_, new_n9377_, new_n9378_,
    new_n9379_, new_n9380_, new_n9381_, new_n9382_, new_n9383_, new_n9384_,
    new_n9385_, new_n9386_, new_n9387_, new_n9388_, new_n9389_, new_n9390_,
    new_n9391_, new_n9392_, new_n9393_, new_n9394_, new_n9395_, new_n9396_,
    new_n9397_, new_n9398_, new_n9399_, new_n9400_, new_n9401_, new_n9402_,
    new_n9403_, new_n9404_, new_n9405_, new_n9406_, new_n9407_, new_n9408_,
    new_n9409_, new_n9410_, new_n9411_, new_n9412_, new_n9413_, new_n9414_,
    new_n9415_, new_n9416_, new_n9417_, new_n9418_, new_n9419_, new_n9420_,
    new_n9421_, new_n9422_, new_n9423_, new_n9424_, new_n9425_, new_n9426_,
    new_n9427_, new_n9428_, new_n9429_, new_n9430_, new_n9431_, new_n9432_,
    new_n9433_, new_n9434_, new_n9435_, new_n9436_, new_n9437_, new_n9438_,
    new_n9439_, new_n9440_, new_n9441_, new_n9442_, new_n9443_, new_n9444_,
    new_n9445_, new_n9446_, new_n9447_, new_n9448_, new_n9449_, new_n9450_,
    new_n9451_, new_n9452_, new_n9453_, new_n9454_, new_n9455_, new_n9456_,
    new_n9457_, new_n9458_, new_n9459_, new_n9460_, new_n9461_, new_n9462_,
    new_n9463_, new_n9464_, new_n9465_, new_n9466_, new_n9467_, new_n9468_,
    new_n9469_, new_n9470_, new_n9471_, new_n9472_, new_n9473_, new_n9474_,
    new_n9475_, new_n9476_, new_n9477_, new_n9478_, new_n9479_, new_n9480_,
    new_n9481_, new_n9482_, new_n9483_, new_n9484_, new_n9485_, new_n9486_,
    new_n9487_, new_n9488_, new_n9489_, new_n9490_, new_n9491_, new_n9492_,
    new_n9493_, new_n9494_, new_n9495_, new_n9496_, new_n9497_, new_n9498_,
    new_n9499_, new_n9500_, new_n9502_, new_n9503_, new_n9504_, new_n9505_,
    new_n9506_, new_n9507_, new_n9508_, new_n9509_, new_n9510_, new_n9511_,
    new_n9512_, new_n9513_, new_n9514_, new_n9515_, new_n9516_, new_n9517_,
    new_n9518_, new_n9519_, new_n9520_, new_n9521_, new_n9522_, new_n9523_,
    new_n9524_, new_n9525_, new_n9526_, new_n9527_, new_n9528_, new_n9529_,
    new_n9530_, new_n9531_, new_n9532_, new_n9533_, new_n9534_, new_n9535_,
    new_n9536_, new_n9537_, new_n9538_, new_n9539_, new_n9540_, new_n9541_,
    new_n9542_, new_n9543_, new_n9544_, new_n9545_, new_n9546_, new_n9547_,
    new_n9548_, new_n9549_, new_n9550_, new_n9551_, new_n9552_, new_n9553_,
    new_n9554_, new_n9555_, new_n9556_, new_n9557_, new_n9558_, new_n9559_,
    new_n9560_, new_n9561_, new_n9562_, new_n9563_, new_n9564_, new_n9565_,
    new_n9566_, new_n9567_, new_n9568_, new_n9569_, new_n9570_, new_n9571_,
    new_n9572_, new_n9573_, new_n9574_, new_n9575_, new_n9576_, new_n9577_,
    new_n9578_, new_n9579_, new_n9580_, new_n9581_, new_n9582_, new_n9583_,
    new_n9584_, new_n9585_, new_n9586_, new_n9587_, new_n9588_, new_n9589_,
    new_n9590_, new_n9591_, new_n9592_, new_n9593_, new_n9594_, new_n9595_,
    new_n9596_, new_n9597_, new_n9598_, new_n9599_, new_n9600_, new_n9601_,
    new_n9602_, new_n9603_, new_n9604_, new_n9605_, new_n9606_, new_n9607_,
    new_n9608_, new_n9609_, new_n9610_, new_n9611_, new_n9612_, new_n9613_,
    new_n9614_, new_n9615_, new_n9616_, new_n9617_, new_n9618_, new_n9619_,
    new_n9620_, new_n9621_, new_n9622_, new_n9623_, new_n9624_, new_n9625_,
    new_n9626_, new_n9627_, new_n9628_, new_n9629_, new_n9630_, new_n9631_,
    new_n9632_, new_n9633_, new_n9634_, new_n9635_, new_n9636_, new_n9637_,
    new_n9638_, new_n9639_, new_n9640_, new_n9641_, new_n9642_, new_n9643_,
    new_n9644_, new_n9645_, new_n9646_, new_n9647_, new_n9648_, new_n9649_,
    new_n9650_, new_n9651_, new_n9652_, new_n9653_, new_n9654_, new_n9655_,
    new_n9656_, new_n9657_, new_n9658_, new_n9659_, new_n9660_, new_n9661_,
    new_n9662_, new_n9663_, new_n9664_, new_n9665_, new_n9666_, new_n9667_,
    new_n9668_, new_n9669_, new_n9670_, new_n9671_, new_n9672_, new_n9673_,
    new_n9674_, new_n9675_, new_n9676_, new_n9677_, new_n9678_, new_n9679_,
    new_n9680_, new_n9681_, new_n9682_, new_n9683_, new_n9684_, new_n9685_,
    new_n9686_, new_n9687_, new_n9688_, new_n9689_, new_n9690_, new_n9691_,
    new_n9692_, new_n9693_, new_n9694_, new_n9695_, new_n9696_, new_n9697_,
    new_n9698_, new_n9699_, new_n9700_, new_n9701_, new_n9702_, new_n9703_,
    new_n9704_, new_n9705_, new_n9706_, new_n9707_, new_n9708_, new_n9709_,
    new_n9710_, new_n9711_, new_n9712_, new_n9713_, new_n9714_, new_n9715_,
    new_n9716_, new_n9717_, new_n9718_, new_n9719_, new_n9720_, new_n9721_,
    new_n9722_, new_n9723_, new_n9724_, new_n9725_, new_n9726_, new_n9727_,
    new_n9728_, new_n9729_, new_n9730_, new_n9731_, new_n9732_, new_n9733_,
    new_n9734_, new_n9735_, new_n9736_, new_n9737_, new_n9738_, new_n9739_,
    new_n9740_, new_n9741_, new_n9742_, new_n9743_, new_n9744_, new_n9745_,
    new_n9746_, new_n9747_, new_n9748_, new_n9749_, new_n9750_, new_n9751_,
    new_n9752_, new_n9753_, new_n9754_, new_n9755_, new_n9756_, new_n9757_,
    new_n9758_, new_n9759_, new_n9760_, new_n9761_, new_n9762_, new_n9763_,
    new_n9764_, new_n9765_, new_n9766_, new_n9767_, new_n9768_, new_n9769_,
    new_n9770_, new_n9771_, new_n9772_, new_n9773_, new_n9774_, new_n9775_,
    new_n9776_, new_n9777_, new_n9778_, new_n9779_, new_n9780_, new_n9781_,
    new_n9782_, new_n9783_, new_n9784_, new_n9785_, new_n9786_, new_n9787_,
    new_n9788_, new_n9789_, new_n9790_, new_n9791_, new_n9792_, new_n9793_,
    new_n9794_, new_n9795_, new_n9796_, new_n9797_, new_n9798_, new_n9799_,
    new_n9800_, new_n9801_, new_n9802_, new_n9803_, new_n9804_, new_n9805_,
    new_n9806_, new_n9807_, new_n9808_, new_n9809_, new_n9810_, new_n9811_,
    new_n9812_, new_n9813_, new_n9814_, new_n9815_, new_n9816_, new_n9817_,
    new_n9818_, new_n9819_, new_n9820_, new_n9821_, new_n9822_, new_n9823_,
    new_n9824_, new_n9825_, new_n9826_, new_n9827_, new_n9828_, new_n9829_,
    new_n9830_, new_n9831_, new_n9832_, new_n9833_, new_n9834_, new_n9835_,
    new_n9836_, new_n9837_, new_n9838_, new_n9839_, new_n9840_, new_n9841_,
    new_n9842_, new_n9843_, new_n9844_, new_n9845_, new_n9846_, new_n9847_,
    new_n9848_, new_n9849_, new_n9850_, new_n9851_, new_n9852_, new_n9853_,
    new_n9854_, new_n9855_, new_n9856_, new_n9857_, new_n9858_, new_n9859_,
    new_n9860_, new_n9861_, new_n9862_, new_n9863_, new_n9864_, new_n9865_,
    new_n9866_, new_n9867_, new_n9868_, new_n9869_, new_n9870_, new_n9871_,
    new_n9872_, new_n9873_, new_n9874_, new_n9875_, new_n9876_, new_n9877_,
    new_n9878_, new_n9879_, new_n9880_, new_n9881_, new_n9882_, new_n9883_,
    new_n9884_, new_n9885_, new_n9886_, new_n9887_, new_n9888_, new_n9889_,
    new_n9890_, new_n9891_, new_n9892_, new_n9893_, new_n9894_, new_n9895_,
    new_n9896_, new_n9897_, new_n9898_, new_n9899_, new_n9900_, new_n9901_,
    new_n9902_, new_n9903_, new_n9904_, new_n9905_, new_n9906_, new_n9907_,
    new_n9908_, new_n9909_, new_n9910_, new_n9911_, new_n9912_, new_n9913_,
    new_n9914_, new_n9915_, new_n9916_, new_n9917_, new_n9918_, new_n9919_,
    new_n9920_, new_n9921_, new_n9922_, new_n9923_, new_n9924_, new_n9925_,
    new_n9926_, new_n9927_, new_n9928_, new_n9929_, new_n9930_, new_n9931_,
    new_n9932_, new_n9933_, new_n9934_, new_n9935_, new_n9936_, new_n9937_,
    new_n9938_, new_n9939_, new_n9940_, new_n9941_, new_n9942_, new_n9943_,
    new_n9944_, new_n9945_, new_n9946_, new_n9947_, new_n9948_, new_n9949_,
    new_n9950_, new_n9951_, new_n9952_, new_n9953_, new_n9954_, new_n9955_,
    new_n9956_, new_n9957_, new_n9958_, new_n9959_, new_n9960_, new_n9961_,
    new_n9962_, new_n9963_, new_n9964_, new_n9965_, new_n9966_, new_n9967_,
    new_n9968_, new_n9969_, new_n9970_, new_n9971_, new_n9972_, new_n9973_,
    new_n9974_, new_n9975_, new_n9976_, new_n9977_, new_n9978_, new_n9979_,
    new_n9980_, new_n9981_, new_n9982_, new_n9983_, new_n9984_, new_n9985_,
    new_n9986_, new_n9987_, new_n9988_, new_n9989_, new_n9990_, new_n9991_,
    new_n9992_, new_n9993_, new_n9994_, new_n9995_, new_n9996_, new_n9997_,
    new_n9998_, new_n9999_, new_n10000_, new_n10001_, new_n10002_,
    new_n10003_, new_n10004_, new_n10006_, new_n10007_, new_n10008_,
    new_n10009_, new_n10010_, new_n10011_, new_n10012_, new_n10013_,
    new_n10014_, new_n10015_, new_n10016_, new_n10017_, new_n10018_,
    new_n10019_, new_n10020_, new_n10021_, new_n10022_, new_n10023_,
    new_n10024_, new_n10025_, new_n10026_, new_n10027_, new_n10028_,
    new_n10029_, new_n10030_, new_n10031_, new_n10032_, new_n10033_,
    new_n10034_, new_n10035_, new_n10036_, new_n10037_, new_n10038_,
    new_n10039_, new_n10040_, new_n10041_, new_n10042_, new_n10043_,
    new_n10044_, new_n10045_, new_n10046_, new_n10047_, new_n10048_,
    new_n10049_, new_n10050_, new_n10051_, new_n10052_, new_n10053_,
    new_n10054_, new_n10055_, new_n10056_, new_n10057_, new_n10058_,
    new_n10059_, new_n10060_, new_n10061_, new_n10062_, new_n10063_,
    new_n10064_, new_n10065_, new_n10066_, new_n10067_, new_n10068_,
    new_n10069_, new_n10070_, new_n10071_, new_n10072_, new_n10073_,
    new_n10074_, new_n10075_, new_n10076_, new_n10077_, new_n10078_,
    new_n10079_, new_n10080_, new_n10081_, new_n10082_, new_n10083_,
    new_n10084_, new_n10085_, new_n10086_, new_n10087_, new_n10088_,
    new_n10089_, new_n10090_, new_n10091_, new_n10092_, new_n10093_,
    new_n10094_, new_n10095_, new_n10096_, new_n10097_, new_n10098_,
    new_n10099_, new_n10100_, new_n10101_, new_n10102_, new_n10103_,
    new_n10104_, new_n10105_, new_n10106_, new_n10107_, new_n10108_,
    new_n10109_, new_n10110_, new_n10111_, new_n10112_, new_n10113_,
    new_n10114_, new_n10115_, new_n10116_, new_n10117_, new_n10118_,
    new_n10119_, new_n10120_, new_n10121_, new_n10122_, new_n10123_,
    new_n10124_, new_n10125_, new_n10126_, new_n10127_, new_n10128_,
    new_n10129_, new_n10130_, new_n10131_, new_n10132_, new_n10133_,
    new_n10134_, new_n10135_, new_n10136_, new_n10137_, new_n10138_,
    new_n10139_, new_n10140_, new_n10141_, new_n10142_, new_n10143_,
    new_n10144_, new_n10145_, new_n10146_, new_n10147_, new_n10148_,
    new_n10149_, new_n10150_, new_n10151_, new_n10152_, new_n10153_,
    new_n10154_, new_n10155_, new_n10156_, new_n10157_, new_n10158_,
    new_n10159_, new_n10160_, new_n10161_, new_n10162_, new_n10163_,
    new_n10164_, new_n10165_, new_n10166_, new_n10167_, new_n10168_,
    new_n10169_, new_n10170_, new_n10171_, new_n10172_, new_n10173_,
    new_n10174_, new_n10175_, new_n10176_, new_n10177_, new_n10178_,
    new_n10179_, new_n10180_, new_n10181_, new_n10182_, new_n10183_,
    new_n10184_, new_n10185_, new_n10186_, new_n10187_, new_n10188_,
    new_n10189_, new_n10190_, new_n10191_, new_n10192_, new_n10193_,
    new_n10194_, new_n10195_, new_n10196_, new_n10197_, new_n10198_,
    new_n10199_, new_n10200_, new_n10201_, new_n10202_, new_n10203_,
    new_n10204_, new_n10205_, new_n10206_, new_n10207_, new_n10208_,
    new_n10209_, new_n10210_, new_n10211_, new_n10212_, new_n10213_,
    new_n10214_, new_n10215_, new_n10216_, new_n10217_, new_n10218_,
    new_n10219_, new_n10220_, new_n10221_, new_n10222_, new_n10223_,
    new_n10224_, new_n10225_, new_n10226_, new_n10227_, new_n10228_,
    new_n10229_, new_n10230_, new_n10231_, new_n10232_, new_n10233_,
    new_n10234_, new_n10235_, new_n10236_, new_n10237_, new_n10238_,
    new_n10239_, new_n10240_, new_n10241_, new_n10242_, new_n10243_,
    new_n10244_, new_n10245_, new_n10246_, new_n10247_, new_n10248_,
    new_n10249_, new_n10250_, new_n10251_, new_n10252_, new_n10253_,
    new_n10254_, new_n10255_, new_n10256_, new_n10257_, new_n10258_,
    new_n10259_, new_n10260_, new_n10261_, new_n10262_, new_n10263_,
    new_n10264_, new_n10265_, new_n10266_, new_n10267_, new_n10268_,
    new_n10269_, new_n10270_, new_n10271_, new_n10272_, new_n10273_,
    new_n10274_, new_n10275_, new_n10276_, new_n10277_, new_n10278_,
    new_n10279_, new_n10280_, new_n10281_, new_n10282_, new_n10283_,
    new_n10284_, new_n10285_, new_n10286_, new_n10287_, new_n10288_,
    new_n10289_, new_n10290_, new_n10291_, new_n10292_, new_n10293_,
    new_n10294_, new_n10295_, new_n10296_, new_n10297_, new_n10298_,
    new_n10299_, new_n10300_, new_n10301_, new_n10302_, new_n10303_,
    new_n10304_, new_n10305_, new_n10306_, new_n10307_, new_n10308_,
    new_n10309_, new_n10310_, new_n10311_, new_n10312_, new_n10313_,
    new_n10314_, new_n10315_, new_n10316_, new_n10317_, new_n10318_,
    new_n10319_, new_n10320_, new_n10321_, new_n10322_, new_n10323_,
    new_n10324_, new_n10325_, new_n10326_, new_n10327_, new_n10328_,
    new_n10329_, new_n10330_, new_n10331_, new_n10332_, new_n10333_,
    new_n10334_, new_n10335_, new_n10336_, new_n10337_, new_n10338_,
    new_n10339_, new_n10340_, new_n10341_, new_n10342_, new_n10343_,
    new_n10344_, new_n10345_, new_n10346_, new_n10347_, new_n10348_,
    new_n10349_, new_n10350_, new_n10351_, new_n10352_, new_n10353_,
    new_n10354_, new_n10355_, new_n10356_, new_n10357_, new_n10358_,
    new_n10359_, new_n10360_, new_n10361_, new_n10362_, new_n10363_,
    new_n10364_, new_n10365_, new_n10366_, new_n10367_, new_n10368_,
    new_n10369_, new_n10370_, new_n10371_, new_n10372_, new_n10373_,
    new_n10374_, new_n10375_, new_n10376_, new_n10377_, new_n10378_,
    new_n10379_, new_n10380_, new_n10381_, new_n10382_, new_n10383_,
    new_n10384_, new_n10385_, new_n10386_, new_n10387_, new_n10388_,
    new_n10389_, new_n10390_, new_n10391_, new_n10392_, new_n10393_,
    new_n10394_, new_n10395_, new_n10396_, new_n10397_, new_n10398_,
    new_n10399_, new_n10400_, new_n10401_, new_n10402_, new_n10403_,
    new_n10404_, new_n10405_, new_n10406_, new_n10407_, new_n10408_,
    new_n10409_, new_n10410_, new_n10411_, new_n10412_, new_n10413_,
    new_n10414_, new_n10415_, new_n10416_, new_n10417_, new_n10418_,
    new_n10419_, new_n10420_, new_n10421_, new_n10422_, new_n10423_,
    new_n10424_, new_n10425_, new_n10426_, new_n10427_, new_n10428_,
    new_n10429_, new_n10430_, new_n10431_, new_n10432_, new_n10433_,
    new_n10434_, new_n10435_, new_n10436_, new_n10437_, new_n10438_,
    new_n10439_, new_n10440_, new_n10441_, new_n10442_, new_n10443_,
    new_n10444_, new_n10445_, new_n10446_, new_n10447_, new_n10448_,
    new_n10449_, new_n10450_, new_n10451_, new_n10452_, new_n10453_,
    new_n10454_, new_n10455_, new_n10456_, new_n10457_, new_n10458_,
    new_n10459_, new_n10460_, new_n10461_, new_n10462_, new_n10463_,
    new_n10464_, new_n10465_, new_n10466_, new_n10467_, new_n10468_,
    new_n10469_, new_n10470_, new_n10471_, new_n10472_, new_n10473_,
    new_n10474_, new_n10475_, new_n10476_, new_n10477_, new_n10478_,
    new_n10479_, new_n10480_, new_n10481_, new_n10482_, new_n10483_,
    new_n10484_, new_n10485_, new_n10486_, new_n10487_, new_n10488_,
    new_n10489_, new_n10490_, new_n10491_, new_n10492_, new_n10493_,
    new_n10494_, new_n10495_, new_n10496_, new_n10497_, new_n10498_,
    new_n10499_, new_n10500_, new_n10501_, new_n10502_, new_n10503_,
    new_n10504_, new_n10505_, new_n10506_, new_n10507_, new_n10508_,
    new_n10509_, new_n10510_, new_n10511_, new_n10512_, new_n10513_,
    new_n10514_, new_n10515_, new_n10516_, new_n10517_, new_n10518_,
    new_n10519_, new_n10520_, new_n10521_, new_n10522_, new_n10523_,
    new_n10524_, new_n10525_, new_n10526_, new_n10527_, new_n10528_,
    new_n10529_, new_n10530_, new_n10532_, new_n10533_, new_n10534_,
    new_n10535_, new_n10536_, new_n10537_, new_n10538_, new_n10539_,
    new_n10540_, new_n10541_, new_n10542_, new_n10543_, new_n10544_,
    new_n10545_, new_n10546_, new_n10547_, new_n10548_, new_n10549_,
    new_n10550_, new_n10551_, new_n10552_, new_n10553_, new_n10554_,
    new_n10555_, new_n10556_, new_n10557_, new_n10558_, new_n10559_,
    new_n10560_, new_n10561_, new_n10562_, new_n10563_, new_n10564_,
    new_n10565_, new_n10566_, new_n10567_, new_n10568_, new_n10569_,
    new_n10570_, new_n10571_, new_n10572_, new_n10573_, new_n10574_,
    new_n10575_, new_n10576_, new_n10577_, new_n10578_, new_n10579_,
    new_n10580_, new_n10581_, new_n10582_, new_n10583_, new_n10584_,
    new_n10585_, new_n10586_, new_n10587_, new_n10588_, new_n10589_,
    new_n10590_, new_n10591_, new_n10592_, new_n10593_, new_n10594_,
    new_n10595_, new_n10596_, new_n10597_, new_n10598_, new_n10599_,
    new_n10600_, new_n10601_, new_n10602_, new_n10603_, new_n10604_,
    new_n10605_, new_n10606_, new_n10607_, new_n10608_, new_n10609_,
    new_n10610_, new_n10611_, new_n10612_, new_n10613_, new_n10614_,
    new_n10615_, new_n10616_, new_n10617_, new_n10618_, new_n10619_,
    new_n10620_, new_n10621_, new_n10622_, new_n10623_, new_n10624_,
    new_n10625_, new_n10626_, new_n10627_, new_n10628_, new_n10629_,
    new_n10630_, new_n10631_, new_n10632_, new_n10633_, new_n10634_,
    new_n10635_, new_n10636_, new_n10637_, new_n10638_, new_n10639_,
    new_n10640_, new_n10641_, new_n10642_, new_n10643_, new_n10644_,
    new_n10645_, new_n10646_, new_n10647_, new_n10648_, new_n10649_,
    new_n10650_, new_n10651_, new_n10652_, new_n10653_, new_n10654_,
    new_n10655_, new_n10656_, new_n10657_, new_n10658_, new_n10659_,
    new_n10660_, new_n10661_, new_n10662_, new_n10663_, new_n10664_,
    new_n10665_, new_n10666_, new_n10667_, new_n10668_, new_n10669_,
    new_n10670_, new_n10671_, new_n10672_, new_n10673_, new_n10674_,
    new_n10675_, new_n10676_, new_n10677_, new_n10678_, new_n10679_,
    new_n10680_, new_n10681_, new_n10682_, new_n10683_, new_n10684_,
    new_n10685_, new_n10686_, new_n10687_, new_n10688_, new_n10689_,
    new_n10690_, new_n10691_, new_n10692_, new_n10693_, new_n10694_,
    new_n10695_, new_n10696_, new_n10697_, new_n10698_, new_n10699_,
    new_n10700_, new_n10701_, new_n10702_, new_n10703_, new_n10704_,
    new_n10705_, new_n10706_, new_n10707_, new_n10708_, new_n10709_,
    new_n10710_, new_n10711_, new_n10712_, new_n10713_, new_n10714_,
    new_n10715_, new_n10716_, new_n10717_, new_n10718_, new_n10719_,
    new_n10720_, new_n10721_, new_n10722_, new_n10723_, new_n10724_,
    new_n10725_, new_n10726_, new_n10727_, new_n10728_, new_n10729_,
    new_n10730_, new_n10731_, new_n10732_, new_n10733_, new_n10734_,
    new_n10735_, new_n10736_, new_n10737_, new_n10738_, new_n10739_,
    new_n10740_, new_n10741_, new_n10742_, new_n10743_, new_n10744_,
    new_n10745_, new_n10746_, new_n10747_, new_n10748_, new_n10749_,
    new_n10750_, new_n10751_, new_n10752_, new_n10753_, new_n10754_,
    new_n10755_, new_n10756_, new_n10757_, new_n10758_, new_n10759_,
    new_n10760_, new_n10761_, new_n10762_, new_n10763_, new_n10764_,
    new_n10765_, new_n10766_, new_n10767_, new_n10768_, new_n10769_,
    new_n10770_, new_n10771_, new_n10772_, new_n10773_, new_n10774_,
    new_n10775_, new_n10776_, new_n10777_, new_n10778_, new_n10779_,
    new_n10780_, new_n10781_, new_n10782_, new_n10783_, new_n10784_,
    new_n10785_, new_n10786_, new_n10787_, new_n10788_, new_n10789_,
    new_n10790_, new_n10791_, new_n10792_, new_n10793_, new_n10794_,
    new_n10795_, new_n10796_, new_n10797_, new_n10798_, new_n10799_,
    new_n10800_, new_n10801_, new_n10802_, new_n10803_, new_n10804_,
    new_n10805_, new_n10806_, new_n10807_, new_n10808_, new_n10809_,
    new_n10810_, new_n10811_, new_n10812_, new_n10813_, new_n10814_,
    new_n10815_, new_n10816_, new_n10817_, new_n10818_, new_n10819_,
    new_n10820_, new_n10821_, new_n10822_, new_n10823_, new_n10824_,
    new_n10825_, new_n10826_, new_n10827_, new_n10828_, new_n10829_,
    new_n10830_, new_n10831_, new_n10832_, new_n10833_, new_n10834_,
    new_n10835_, new_n10836_, new_n10837_, new_n10838_, new_n10839_,
    new_n10840_, new_n10841_, new_n10842_, new_n10843_, new_n10844_,
    new_n10845_, new_n10846_, new_n10847_, new_n10848_, new_n10849_,
    new_n10850_, new_n10851_, new_n10852_, new_n10853_, new_n10854_,
    new_n10855_, new_n10856_, new_n10857_, new_n10858_, new_n10859_,
    new_n10860_, new_n10861_, new_n10862_, new_n10863_, new_n10864_,
    new_n10865_, new_n10866_, new_n10867_, new_n10868_, new_n10869_,
    new_n10870_, new_n10871_, new_n10872_, new_n10873_, new_n10874_,
    new_n10875_, new_n10876_, new_n10877_, new_n10878_, new_n10879_,
    new_n10880_, new_n10881_, new_n10882_, new_n10883_, new_n10884_,
    new_n10885_, new_n10886_, new_n10887_, new_n10888_, new_n10889_,
    new_n10890_, new_n10891_, new_n10892_, new_n10893_, new_n10894_,
    new_n10895_, new_n10896_, new_n10897_, new_n10898_, new_n10899_,
    new_n10900_, new_n10901_, new_n10902_, new_n10903_, new_n10904_,
    new_n10905_, new_n10906_, new_n10907_, new_n10908_, new_n10909_,
    new_n10910_, new_n10911_, new_n10912_, new_n10913_, new_n10914_,
    new_n10915_, new_n10916_, new_n10917_, new_n10918_, new_n10919_,
    new_n10920_, new_n10921_, new_n10922_, new_n10923_, new_n10924_,
    new_n10925_, new_n10926_, new_n10927_, new_n10928_, new_n10929_,
    new_n10930_, new_n10931_, new_n10932_, new_n10933_, new_n10934_,
    new_n10935_, new_n10936_, new_n10937_, new_n10938_, new_n10939_,
    new_n10940_, new_n10941_, new_n10942_, new_n10943_, new_n10944_,
    new_n10945_, new_n10946_, new_n10947_, new_n10948_, new_n10949_,
    new_n10950_, new_n10951_, new_n10952_, new_n10953_, new_n10954_,
    new_n10955_, new_n10956_, new_n10957_, new_n10958_, new_n10959_,
    new_n10960_, new_n10961_, new_n10962_, new_n10963_, new_n10964_,
    new_n10965_, new_n10966_, new_n10967_, new_n10968_, new_n10969_,
    new_n10970_, new_n10971_, new_n10972_, new_n10973_, new_n10974_,
    new_n10975_, new_n10976_, new_n10977_, new_n10978_, new_n10979_,
    new_n10980_, new_n10981_, new_n10982_, new_n10983_, new_n10984_,
    new_n10985_, new_n10986_, new_n10987_, new_n10988_, new_n10989_,
    new_n10990_, new_n10991_, new_n10992_, new_n10993_, new_n10994_,
    new_n10995_, new_n10996_, new_n10997_, new_n10998_, new_n10999_,
    new_n11000_, new_n11001_, new_n11002_, new_n11003_, new_n11004_,
    new_n11005_, new_n11006_, new_n11007_, new_n11008_, new_n11009_,
    new_n11010_, new_n11011_, new_n11012_, new_n11013_, new_n11014_,
    new_n11015_, new_n11016_, new_n11017_, new_n11018_, new_n11019_,
    new_n11020_, new_n11021_, new_n11022_, new_n11023_, new_n11024_,
    new_n11025_, new_n11026_, new_n11027_, new_n11028_, new_n11029_,
    new_n11030_, new_n11031_, new_n11032_, new_n11033_, new_n11034_,
    new_n11035_, new_n11036_, new_n11037_, new_n11038_, new_n11039_,
    new_n11040_, new_n11041_, new_n11042_, new_n11043_, new_n11044_,
    new_n11045_, new_n11046_, new_n11047_, new_n11048_, new_n11049_,
    new_n11050_, new_n11051_, new_n11052_, new_n11053_, new_n11054_,
    new_n11055_, new_n11056_, new_n11057_, new_n11058_, new_n11059_,
    new_n11060_, new_n11061_, new_n11062_, new_n11063_, new_n11064_,
    new_n11065_, new_n11066_, new_n11067_, new_n11068_, new_n11069_,
    new_n11070_, new_n11071_, new_n11072_, new_n11074_, new_n11075_,
    new_n11076_, new_n11077_, new_n11078_, new_n11079_, new_n11080_,
    new_n11081_, new_n11082_, new_n11083_, new_n11084_, new_n11085_,
    new_n11086_, new_n11087_, new_n11088_, new_n11089_, new_n11090_,
    new_n11091_, new_n11092_, new_n11093_, new_n11094_, new_n11095_,
    new_n11096_, new_n11097_, new_n11098_, new_n11099_, new_n11100_,
    new_n11101_, new_n11102_, new_n11103_, new_n11104_, new_n11105_,
    new_n11106_, new_n11107_, new_n11108_, new_n11109_, new_n11110_,
    new_n11111_, new_n11112_, new_n11113_, new_n11114_, new_n11115_,
    new_n11116_, new_n11117_, new_n11118_, new_n11119_, new_n11120_,
    new_n11121_, new_n11122_, new_n11123_, new_n11124_, new_n11125_,
    new_n11126_, new_n11127_, new_n11128_, new_n11129_, new_n11130_,
    new_n11131_, new_n11132_, new_n11133_, new_n11134_, new_n11135_,
    new_n11136_, new_n11137_, new_n11138_, new_n11139_, new_n11140_,
    new_n11141_, new_n11142_, new_n11143_, new_n11144_, new_n11145_,
    new_n11146_, new_n11147_, new_n11148_, new_n11149_, new_n11150_,
    new_n11151_, new_n11152_, new_n11153_, new_n11154_, new_n11155_,
    new_n11156_, new_n11157_, new_n11158_, new_n11159_, new_n11160_,
    new_n11161_, new_n11162_, new_n11163_, new_n11164_, new_n11165_,
    new_n11166_, new_n11167_, new_n11168_, new_n11169_, new_n11170_,
    new_n11171_, new_n11172_, new_n11173_, new_n11174_, new_n11175_,
    new_n11176_, new_n11177_, new_n11178_, new_n11179_, new_n11180_,
    new_n11181_, new_n11182_, new_n11183_, new_n11184_, new_n11185_,
    new_n11186_, new_n11187_, new_n11188_, new_n11189_, new_n11190_,
    new_n11191_, new_n11192_, new_n11193_, new_n11194_, new_n11195_,
    new_n11196_, new_n11197_, new_n11198_, new_n11199_, new_n11200_,
    new_n11201_, new_n11202_, new_n11203_, new_n11204_, new_n11205_,
    new_n11206_, new_n11207_, new_n11208_, new_n11209_, new_n11210_,
    new_n11211_, new_n11212_, new_n11213_, new_n11214_, new_n11215_,
    new_n11216_, new_n11217_, new_n11218_, new_n11219_, new_n11220_,
    new_n11221_, new_n11222_, new_n11223_, new_n11224_, new_n11225_,
    new_n11226_, new_n11227_, new_n11228_, new_n11229_, new_n11230_,
    new_n11231_, new_n11232_, new_n11233_, new_n11234_, new_n11235_,
    new_n11236_, new_n11237_, new_n11238_, new_n11239_, new_n11240_,
    new_n11241_, new_n11242_, new_n11243_, new_n11244_, new_n11245_,
    new_n11246_, new_n11247_, new_n11248_, new_n11249_, new_n11250_,
    new_n11251_, new_n11252_, new_n11253_, new_n11254_, new_n11255_,
    new_n11256_, new_n11257_, new_n11258_, new_n11259_, new_n11260_,
    new_n11261_, new_n11262_, new_n11263_, new_n11264_, new_n11265_,
    new_n11266_, new_n11267_, new_n11268_, new_n11269_, new_n11270_,
    new_n11271_, new_n11272_, new_n11273_, new_n11274_, new_n11275_,
    new_n11276_, new_n11277_, new_n11278_, new_n11279_, new_n11280_,
    new_n11281_, new_n11282_, new_n11283_, new_n11284_, new_n11285_,
    new_n11286_, new_n11287_, new_n11288_, new_n11289_, new_n11290_,
    new_n11291_, new_n11292_, new_n11293_, new_n11294_, new_n11295_,
    new_n11296_, new_n11297_, new_n11298_, new_n11299_, new_n11300_,
    new_n11301_, new_n11302_, new_n11303_, new_n11304_, new_n11305_,
    new_n11306_, new_n11307_, new_n11308_, new_n11309_, new_n11310_,
    new_n11311_, new_n11312_, new_n11313_, new_n11314_, new_n11315_,
    new_n11316_, new_n11317_, new_n11318_, new_n11319_, new_n11320_,
    new_n11321_, new_n11322_, new_n11323_, new_n11324_, new_n11325_,
    new_n11326_, new_n11327_, new_n11328_, new_n11329_, new_n11330_,
    new_n11331_, new_n11332_, new_n11333_, new_n11334_, new_n11335_,
    new_n11336_, new_n11337_, new_n11338_, new_n11339_, new_n11340_,
    new_n11341_, new_n11342_, new_n11343_, new_n11344_, new_n11345_,
    new_n11346_, new_n11347_, new_n11348_, new_n11349_, new_n11350_,
    new_n11351_, new_n11352_, new_n11353_, new_n11354_, new_n11355_,
    new_n11356_, new_n11357_, new_n11358_, new_n11359_, new_n11360_,
    new_n11361_, new_n11362_, new_n11363_, new_n11364_, new_n11365_,
    new_n11366_, new_n11367_, new_n11368_, new_n11369_, new_n11370_,
    new_n11371_, new_n11372_, new_n11373_, new_n11374_, new_n11375_,
    new_n11376_, new_n11377_, new_n11378_, new_n11379_, new_n11380_,
    new_n11381_, new_n11382_, new_n11383_, new_n11384_, new_n11385_,
    new_n11386_, new_n11387_, new_n11388_, new_n11389_, new_n11390_,
    new_n11391_, new_n11392_, new_n11393_, new_n11394_, new_n11395_,
    new_n11396_, new_n11397_, new_n11398_, new_n11399_, new_n11400_,
    new_n11401_, new_n11402_, new_n11403_, new_n11404_, new_n11405_,
    new_n11406_, new_n11407_, new_n11408_, new_n11409_, new_n11410_,
    new_n11411_, new_n11412_, new_n11413_, new_n11414_, new_n11415_,
    new_n11416_, new_n11417_, new_n11418_, new_n11419_, new_n11420_,
    new_n11421_, new_n11422_, new_n11423_, new_n11424_, new_n11425_,
    new_n11426_, new_n11427_, new_n11428_, new_n11429_, new_n11430_,
    new_n11431_, new_n11432_, new_n11433_, new_n11434_, new_n11435_,
    new_n11436_, new_n11437_, new_n11438_, new_n11439_, new_n11440_,
    new_n11441_, new_n11442_, new_n11443_, new_n11444_, new_n11445_,
    new_n11446_, new_n11447_, new_n11448_, new_n11449_, new_n11450_,
    new_n11451_, new_n11452_, new_n11453_, new_n11454_, new_n11455_,
    new_n11456_, new_n11457_, new_n11458_, new_n11459_, new_n11460_,
    new_n11461_, new_n11462_, new_n11463_, new_n11464_, new_n11465_,
    new_n11466_, new_n11467_, new_n11468_, new_n11469_, new_n11470_,
    new_n11471_, new_n11472_, new_n11473_, new_n11474_, new_n11475_,
    new_n11476_, new_n11477_, new_n11478_, new_n11479_, new_n11480_,
    new_n11481_, new_n11482_, new_n11483_, new_n11484_, new_n11485_,
    new_n11486_, new_n11487_, new_n11488_, new_n11489_, new_n11490_,
    new_n11491_, new_n11492_, new_n11493_, new_n11494_, new_n11495_,
    new_n11496_, new_n11497_, new_n11498_, new_n11499_, new_n11500_,
    new_n11501_, new_n11502_, new_n11503_, new_n11504_, new_n11505_,
    new_n11506_, new_n11507_, new_n11508_, new_n11509_, new_n11510_,
    new_n11511_, new_n11512_, new_n11513_, new_n11514_, new_n11515_,
    new_n11516_, new_n11517_, new_n11518_, new_n11519_, new_n11520_,
    new_n11521_, new_n11522_, new_n11523_, new_n11524_, new_n11525_,
    new_n11526_, new_n11527_, new_n11528_, new_n11529_, new_n11530_,
    new_n11531_, new_n11532_, new_n11533_, new_n11534_, new_n11535_,
    new_n11536_, new_n11537_, new_n11538_, new_n11539_, new_n11540_,
    new_n11541_, new_n11542_, new_n11543_, new_n11544_, new_n11545_,
    new_n11546_, new_n11547_, new_n11548_, new_n11549_, new_n11550_,
    new_n11551_, new_n11552_, new_n11553_, new_n11554_, new_n11555_,
    new_n11556_, new_n11557_, new_n11558_, new_n11559_, new_n11560_,
    new_n11561_, new_n11562_, new_n11563_, new_n11564_, new_n11565_,
    new_n11566_, new_n11567_, new_n11568_, new_n11569_, new_n11570_,
    new_n11571_, new_n11572_, new_n11573_, new_n11574_, new_n11575_,
    new_n11576_, new_n11577_, new_n11578_, new_n11579_, new_n11580_,
    new_n11581_, new_n11582_, new_n11583_, new_n11584_, new_n11585_,
    new_n11586_, new_n11587_, new_n11588_, new_n11589_, new_n11590_,
    new_n11591_, new_n11592_, new_n11593_, new_n11594_, new_n11595_,
    new_n11596_, new_n11597_, new_n11598_, new_n11599_, new_n11600_,
    new_n11601_, new_n11602_, new_n11603_, new_n11604_, new_n11605_,
    new_n11606_, new_n11607_, new_n11608_, new_n11609_, new_n11610_,
    new_n11611_, new_n11612_, new_n11613_, new_n11614_, new_n11615_,
    new_n11616_, new_n11617_, new_n11618_, new_n11619_, new_n11621_,
    new_n11622_, new_n11623_, new_n11624_, new_n11625_, new_n11626_,
    new_n11627_, new_n11628_, new_n11629_, new_n11630_, new_n11631_,
    new_n11632_, new_n11633_, new_n11634_, new_n11635_, new_n11636_,
    new_n11637_, new_n11638_, new_n11639_, new_n11640_, new_n11641_,
    new_n11642_, new_n11643_, new_n11644_, new_n11645_, new_n11646_,
    new_n11647_, new_n11648_, new_n11649_, new_n11650_, new_n11651_,
    new_n11652_, new_n11653_, new_n11654_, new_n11655_, new_n11656_,
    new_n11657_, new_n11658_, new_n11659_, new_n11660_, new_n11661_,
    new_n11662_, new_n11663_, new_n11664_, new_n11665_, new_n11666_,
    new_n11667_, new_n11668_, new_n11669_, new_n11670_, new_n11671_,
    new_n11672_, new_n11673_, new_n11674_, new_n11675_, new_n11676_,
    new_n11677_, new_n11678_, new_n11679_, new_n11680_, new_n11681_,
    new_n11682_, new_n11683_, new_n11684_, new_n11685_, new_n11686_,
    new_n11687_, new_n11688_, new_n11689_, new_n11690_, new_n11691_,
    new_n11692_, new_n11693_, new_n11694_, new_n11695_, new_n11696_,
    new_n11697_, new_n11698_, new_n11699_, new_n11700_, new_n11701_,
    new_n11702_, new_n11703_, new_n11704_, new_n11705_, new_n11706_,
    new_n11707_, new_n11708_, new_n11709_, new_n11710_, new_n11711_,
    new_n11712_, new_n11713_, new_n11714_, new_n11715_, new_n11716_,
    new_n11717_, new_n11718_, new_n11719_, new_n11720_, new_n11721_,
    new_n11722_, new_n11723_, new_n11724_, new_n11725_, new_n11726_,
    new_n11727_, new_n11728_, new_n11729_, new_n11730_, new_n11731_,
    new_n11732_, new_n11733_, new_n11734_, new_n11735_, new_n11736_,
    new_n11737_, new_n11738_, new_n11739_, new_n11740_, new_n11741_,
    new_n11742_, new_n11743_, new_n11744_, new_n11745_, new_n11746_,
    new_n11747_, new_n11748_, new_n11749_, new_n11750_, new_n11751_,
    new_n11752_, new_n11753_, new_n11754_, new_n11755_, new_n11756_,
    new_n11757_, new_n11758_, new_n11759_, new_n11760_, new_n11761_,
    new_n11762_, new_n11763_, new_n11764_, new_n11765_, new_n11766_,
    new_n11767_, new_n11768_, new_n11769_, new_n11770_, new_n11771_,
    new_n11772_, new_n11773_, new_n11774_, new_n11775_, new_n11776_,
    new_n11777_, new_n11778_, new_n11779_, new_n11780_, new_n11781_,
    new_n11782_, new_n11783_, new_n11784_, new_n11785_, new_n11786_,
    new_n11787_, new_n11788_, new_n11789_, new_n11790_, new_n11791_,
    new_n11792_, new_n11793_, new_n11794_, new_n11795_, new_n11796_,
    new_n11797_, new_n11798_, new_n11799_, new_n11800_, new_n11801_,
    new_n11802_, new_n11803_, new_n11804_, new_n11805_, new_n11806_,
    new_n11807_, new_n11808_, new_n11809_, new_n11810_, new_n11811_,
    new_n11812_, new_n11813_, new_n11814_, new_n11815_, new_n11816_,
    new_n11817_, new_n11818_, new_n11819_, new_n11820_, new_n11821_,
    new_n11822_, new_n11823_, new_n11824_, new_n11825_, new_n11826_,
    new_n11827_, new_n11828_, new_n11829_, new_n11830_, new_n11831_,
    new_n11832_, new_n11833_, new_n11834_, new_n11835_, new_n11836_,
    new_n11837_, new_n11838_, new_n11839_, new_n11840_, new_n11841_,
    new_n11842_, new_n11843_, new_n11844_, new_n11845_, new_n11846_,
    new_n11847_, new_n11848_, new_n11849_, new_n11850_, new_n11851_,
    new_n11852_, new_n11853_, new_n11854_, new_n11855_, new_n11856_,
    new_n11857_, new_n11858_, new_n11859_, new_n11860_, new_n11861_,
    new_n11862_, new_n11863_, new_n11864_, new_n11865_, new_n11866_,
    new_n11867_, new_n11868_, new_n11869_, new_n11870_, new_n11871_,
    new_n11872_, new_n11873_, new_n11874_, new_n11875_, new_n11876_,
    new_n11877_, new_n11878_, new_n11879_, new_n11880_, new_n11881_,
    new_n11882_, new_n11883_, new_n11884_, new_n11885_, new_n11886_,
    new_n11887_, new_n11888_, new_n11889_, new_n11890_, new_n11891_,
    new_n11892_, new_n11893_, new_n11894_, new_n11895_, new_n11896_,
    new_n11897_, new_n11898_, new_n11899_, new_n11900_, new_n11901_,
    new_n11902_, new_n11903_, new_n11904_, new_n11905_, new_n11906_,
    new_n11907_, new_n11908_, new_n11909_, new_n11910_, new_n11911_,
    new_n11912_, new_n11913_, new_n11914_, new_n11915_, new_n11916_,
    new_n11917_, new_n11918_, new_n11919_, new_n11920_, new_n11921_,
    new_n11922_, new_n11923_, new_n11924_, new_n11925_, new_n11926_,
    new_n11927_, new_n11928_, new_n11929_, new_n11930_, new_n11931_,
    new_n11932_, new_n11933_, new_n11934_, new_n11935_, new_n11936_,
    new_n11937_, new_n11938_, new_n11939_, new_n11940_, new_n11941_,
    new_n11942_, new_n11943_, new_n11944_, new_n11945_, new_n11946_,
    new_n11947_, new_n11948_, new_n11949_, new_n11950_, new_n11951_,
    new_n11952_, new_n11953_, new_n11954_, new_n11955_, new_n11956_,
    new_n11957_, new_n11958_, new_n11959_, new_n11960_, new_n11961_,
    new_n11962_, new_n11963_, new_n11964_, new_n11965_, new_n11966_,
    new_n11967_, new_n11968_, new_n11969_, new_n11970_, new_n11971_,
    new_n11972_, new_n11973_, new_n11974_, new_n11975_, new_n11976_,
    new_n11977_, new_n11978_, new_n11979_, new_n11980_, new_n11981_,
    new_n11982_, new_n11983_, new_n11984_, new_n11985_, new_n11986_,
    new_n11987_, new_n11988_, new_n11989_, new_n11990_, new_n11991_,
    new_n11992_, new_n11993_, new_n11994_, new_n11995_, new_n11996_,
    new_n11997_, new_n11998_, new_n11999_, new_n12000_, new_n12001_,
    new_n12002_, new_n12003_, new_n12004_, new_n12005_, new_n12006_,
    new_n12007_, new_n12008_, new_n12009_, new_n12010_, new_n12011_,
    new_n12012_, new_n12013_, new_n12014_, new_n12015_, new_n12016_,
    new_n12017_, new_n12018_, new_n12019_, new_n12020_, new_n12021_,
    new_n12022_, new_n12023_, new_n12024_, new_n12025_, new_n12026_,
    new_n12027_, new_n12028_, new_n12029_, new_n12030_, new_n12031_,
    new_n12032_, new_n12033_, new_n12034_, new_n12035_, new_n12036_,
    new_n12037_, new_n12038_, new_n12039_, new_n12040_, new_n12041_,
    new_n12042_, new_n12043_, new_n12044_, new_n12045_, new_n12046_,
    new_n12047_, new_n12048_, new_n12049_, new_n12050_, new_n12051_,
    new_n12052_, new_n12053_, new_n12054_, new_n12055_, new_n12056_,
    new_n12057_, new_n12058_, new_n12059_, new_n12060_, new_n12061_,
    new_n12062_, new_n12063_, new_n12064_, new_n12065_, new_n12066_,
    new_n12067_, new_n12068_, new_n12069_, new_n12070_, new_n12071_,
    new_n12072_, new_n12073_, new_n12074_, new_n12075_, new_n12076_,
    new_n12077_, new_n12078_, new_n12079_, new_n12080_, new_n12081_,
    new_n12082_, new_n12083_, new_n12084_, new_n12085_, new_n12086_,
    new_n12087_, new_n12088_, new_n12089_, new_n12090_, new_n12091_,
    new_n12092_, new_n12093_, new_n12094_, new_n12095_, new_n12096_,
    new_n12097_, new_n12098_, new_n12099_, new_n12100_, new_n12101_,
    new_n12102_, new_n12103_, new_n12104_, new_n12105_, new_n12106_,
    new_n12107_, new_n12108_, new_n12109_, new_n12110_, new_n12111_,
    new_n12112_, new_n12113_, new_n12114_, new_n12115_, new_n12116_,
    new_n12117_, new_n12118_, new_n12119_, new_n12120_, new_n12121_,
    new_n12122_, new_n12123_, new_n12124_, new_n12125_, new_n12126_,
    new_n12127_, new_n12128_, new_n12129_, new_n12130_, new_n12131_,
    new_n12132_, new_n12133_, new_n12134_, new_n12135_, new_n12136_,
    new_n12137_, new_n12138_, new_n12139_, new_n12140_, new_n12141_,
    new_n12142_, new_n12143_, new_n12144_, new_n12145_, new_n12146_,
    new_n12147_, new_n12148_, new_n12149_, new_n12150_, new_n12151_,
    new_n12152_, new_n12153_, new_n12154_, new_n12155_, new_n12156_,
    new_n12157_, new_n12158_, new_n12159_, new_n12160_, new_n12161_,
    new_n12162_, new_n12163_, new_n12164_, new_n12165_, new_n12166_,
    new_n12167_, new_n12168_, new_n12169_, new_n12170_, new_n12171_,
    new_n12172_, new_n12173_, new_n12174_, new_n12175_, new_n12176_,
    new_n12177_, new_n12178_, new_n12179_, new_n12180_, new_n12181_,
    new_n12182_, new_n12183_, new_n12184_, new_n12186_, new_n12187_,
    new_n12188_, new_n12189_, new_n12190_, new_n12191_, new_n12192_,
    new_n12193_, new_n12194_, new_n12195_, new_n12196_, new_n12197_,
    new_n12198_, new_n12199_, new_n12200_, new_n12201_, new_n12202_,
    new_n12203_, new_n12204_, new_n12205_, new_n12206_, new_n12207_,
    new_n12208_, new_n12209_, new_n12210_, new_n12211_, new_n12212_,
    new_n12213_, new_n12214_, new_n12215_, new_n12216_, new_n12217_,
    new_n12218_, new_n12219_, new_n12220_, new_n12221_, new_n12222_,
    new_n12223_, new_n12224_, new_n12225_, new_n12226_, new_n12227_,
    new_n12228_, new_n12229_, new_n12230_, new_n12231_, new_n12232_,
    new_n12233_, new_n12234_, new_n12235_, new_n12236_, new_n12237_,
    new_n12238_, new_n12239_, new_n12240_, new_n12241_, new_n12242_,
    new_n12243_, new_n12244_, new_n12245_, new_n12246_, new_n12247_,
    new_n12248_, new_n12249_, new_n12250_, new_n12251_, new_n12252_,
    new_n12253_, new_n12254_, new_n12255_, new_n12256_, new_n12257_,
    new_n12258_, new_n12259_, new_n12260_, new_n12261_, new_n12262_,
    new_n12263_, new_n12264_, new_n12265_, new_n12266_, new_n12267_,
    new_n12268_, new_n12269_, new_n12270_, new_n12271_, new_n12272_,
    new_n12273_, new_n12274_, new_n12275_, new_n12276_, new_n12277_,
    new_n12278_, new_n12279_, new_n12280_, new_n12281_, new_n12282_,
    new_n12283_, new_n12284_, new_n12285_, new_n12286_, new_n12287_,
    new_n12288_, new_n12289_, new_n12290_, new_n12291_, new_n12292_,
    new_n12293_, new_n12294_, new_n12295_, new_n12296_, new_n12297_,
    new_n12298_, new_n12299_, new_n12300_, new_n12301_, new_n12302_,
    new_n12303_, new_n12304_, new_n12305_, new_n12306_, new_n12307_,
    new_n12308_, new_n12309_, new_n12310_, new_n12311_, new_n12312_,
    new_n12313_, new_n12314_, new_n12315_, new_n12316_, new_n12317_,
    new_n12318_, new_n12319_, new_n12320_, new_n12321_, new_n12322_,
    new_n12323_, new_n12324_, new_n12325_, new_n12326_, new_n12327_,
    new_n12328_, new_n12329_, new_n12330_, new_n12331_, new_n12332_,
    new_n12333_, new_n12334_, new_n12335_, new_n12336_, new_n12337_,
    new_n12338_, new_n12339_, new_n12340_, new_n12341_, new_n12342_,
    new_n12343_, new_n12344_, new_n12345_, new_n12346_, new_n12347_,
    new_n12348_, new_n12349_, new_n12350_, new_n12351_, new_n12352_,
    new_n12353_, new_n12354_, new_n12355_, new_n12356_, new_n12357_,
    new_n12358_, new_n12359_, new_n12360_, new_n12361_, new_n12362_,
    new_n12363_, new_n12364_, new_n12365_, new_n12366_, new_n12367_,
    new_n12368_, new_n12369_, new_n12370_, new_n12371_, new_n12372_,
    new_n12373_, new_n12374_, new_n12375_, new_n12376_, new_n12377_,
    new_n12378_, new_n12379_, new_n12380_, new_n12381_, new_n12382_,
    new_n12383_, new_n12384_, new_n12385_, new_n12386_, new_n12387_,
    new_n12388_, new_n12389_, new_n12390_, new_n12391_, new_n12392_,
    new_n12393_, new_n12394_, new_n12395_, new_n12396_, new_n12397_,
    new_n12398_, new_n12399_, new_n12400_, new_n12401_, new_n12402_,
    new_n12403_, new_n12404_, new_n12405_, new_n12406_, new_n12407_,
    new_n12408_, new_n12409_, new_n12410_, new_n12411_, new_n12412_,
    new_n12413_, new_n12414_, new_n12415_, new_n12416_, new_n12417_,
    new_n12418_, new_n12419_, new_n12420_, new_n12421_, new_n12422_,
    new_n12423_, new_n12424_, new_n12425_, new_n12426_, new_n12427_,
    new_n12428_, new_n12429_, new_n12430_, new_n12431_, new_n12432_,
    new_n12433_, new_n12434_, new_n12435_, new_n12436_, new_n12437_,
    new_n12438_, new_n12439_, new_n12440_, new_n12441_, new_n12442_,
    new_n12443_, new_n12444_, new_n12445_, new_n12446_, new_n12447_,
    new_n12448_, new_n12449_, new_n12450_, new_n12451_, new_n12452_,
    new_n12453_, new_n12454_, new_n12455_, new_n12456_, new_n12457_,
    new_n12458_, new_n12459_, new_n12460_, new_n12461_, new_n12462_,
    new_n12463_, new_n12464_, new_n12465_, new_n12466_, new_n12467_,
    new_n12468_, new_n12469_, new_n12470_, new_n12471_, new_n12472_,
    new_n12473_, new_n12474_, new_n12475_, new_n12476_, new_n12477_,
    new_n12478_, new_n12479_, new_n12480_, new_n12481_, new_n12482_,
    new_n12483_, new_n12484_, new_n12485_, new_n12486_, new_n12487_,
    new_n12488_, new_n12489_, new_n12490_, new_n12491_, new_n12492_,
    new_n12493_, new_n12494_, new_n12495_, new_n12496_, new_n12497_,
    new_n12498_, new_n12499_, new_n12500_, new_n12501_, new_n12502_,
    new_n12503_, new_n12504_, new_n12505_, new_n12506_, new_n12507_,
    new_n12508_, new_n12509_, new_n12510_, new_n12511_, new_n12512_,
    new_n12513_, new_n12514_, new_n12515_, new_n12516_, new_n12517_,
    new_n12518_, new_n12519_, new_n12520_, new_n12521_, new_n12522_,
    new_n12523_, new_n12524_, new_n12525_, new_n12526_, new_n12527_,
    new_n12528_, new_n12529_, new_n12530_, new_n12531_, new_n12532_,
    new_n12533_, new_n12534_, new_n12535_, new_n12536_, new_n12537_,
    new_n12538_, new_n12539_, new_n12540_, new_n12541_, new_n12542_,
    new_n12543_, new_n12544_, new_n12545_, new_n12546_, new_n12547_,
    new_n12548_, new_n12549_, new_n12550_, new_n12551_, new_n12552_,
    new_n12553_, new_n12554_, new_n12555_, new_n12556_, new_n12557_,
    new_n12558_, new_n12559_, new_n12560_, new_n12561_, new_n12562_,
    new_n12563_, new_n12564_, new_n12565_, new_n12566_, new_n12567_,
    new_n12568_, new_n12569_, new_n12570_, new_n12571_, new_n12572_,
    new_n12573_, new_n12574_, new_n12575_, new_n12576_, new_n12577_,
    new_n12578_, new_n12579_, new_n12580_, new_n12581_, new_n12582_,
    new_n12583_, new_n12584_, new_n12585_, new_n12586_, new_n12587_,
    new_n12588_, new_n12589_, new_n12590_, new_n12591_, new_n12592_,
    new_n12593_, new_n12594_, new_n12595_, new_n12596_, new_n12597_,
    new_n12598_, new_n12599_, new_n12600_, new_n12601_, new_n12602_,
    new_n12603_, new_n12604_, new_n12605_, new_n12606_, new_n12607_,
    new_n12608_, new_n12609_, new_n12610_, new_n12611_, new_n12612_,
    new_n12613_, new_n12614_, new_n12615_, new_n12616_, new_n12617_,
    new_n12618_, new_n12619_, new_n12620_, new_n12621_, new_n12622_,
    new_n12623_, new_n12624_, new_n12625_, new_n12626_, new_n12627_,
    new_n12628_, new_n12629_, new_n12630_, new_n12631_, new_n12632_,
    new_n12633_, new_n12634_, new_n12635_, new_n12636_, new_n12637_,
    new_n12638_, new_n12639_, new_n12640_, new_n12641_, new_n12642_,
    new_n12643_, new_n12644_, new_n12645_, new_n12646_, new_n12647_,
    new_n12648_, new_n12649_, new_n12650_, new_n12651_, new_n12652_,
    new_n12653_, new_n12654_, new_n12655_, new_n12656_, new_n12657_,
    new_n12658_, new_n12659_, new_n12660_, new_n12661_, new_n12662_,
    new_n12663_, new_n12664_, new_n12665_, new_n12666_, new_n12667_,
    new_n12668_, new_n12669_, new_n12670_, new_n12671_, new_n12672_,
    new_n12673_, new_n12674_, new_n12675_, new_n12676_, new_n12677_,
    new_n12678_, new_n12679_, new_n12680_, new_n12681_, new_n12682_,
    new_n12683_, new_n12684_, new_n12685_, new_n12686_, new_n12687_,
    new_n12688_, new_n12689_, new_n12690_, new_n12691_, new_n12692_,
    new_n12693_, new_n12694_, new_n12695_, new_n12696_, new_n12697_,
    new_n12698_, new_n12699_, new_n12700_, new_n12701_, new_n12702_,
    new_n12703_, new_n12704_, new_n12705_, new_n12706_, new_n12707_,
    new_n12708_, new_n12709_, new_n12710_, new_n12711_, new_n12712_,
    new_n12713_, new_n12714_, new_n12715_, new_n12716_, new_n12717_,
    new_n12718_, new_n12719_, new_n12720_, new_n12721_, new_n12722_,
    new_n12723_, new_n12724_, new_n12725_, new_n12726_, new_n12727_,
    new_n12728_, new_n12729_, new_n12730_, new_n12731_, new_n12732_,
    new_n12733_, new_n12734_, new_n12735_, new_n12736_, new_n12737_,
    new_n12738_, new_n12739_, new_n12740_, new_n12741_, new_n12742_,
    new_n12743_, new_n12744_, new_n12745_, new_n12746_, new_n12747_,
    new_n12748_, new_n12749_, new_n12750_, new_n12751_, new_n12752_,
    new_n12753_, new_n12754_, new_n12755_, new_n12756_, new_n12757_,
    new_n12758_, new_n12759_, new_n12760_, new_n12761_, new_n12762_,
    new_n12763_, new_n12764_, new_n12765_, new_n12767_, new_n12768_,
    new_n12769_, new_n12770_, new_n12771_, new_n12772_, new_n12773_,
    new_n12774_, new_n12775_, new_n12776_, new_n12777_, new_n12778_,
    new_n12779_, new_n12780_, new_n12781_, new_n12782_, new_n12783_,
    new_n12784_, new_n12785_, new_n12786_, new_n12787_, new_n12788_,
    new_n12789_, new_n12790_, new_n12791_, new_n12792_, new_n12793_,
    new_n12794_, new_n12795_, new_n12796_, new_n12797_, new_n12798_,
    new_n12799_, new_n12800_, new_n12801_, new_n12802_, new_n12803_,
    new_n12804_, new_n12805_, new_n12806_, new_n12807_, new_n12808_,
    new_n12809_, new_n12810_, new_n12811_, new_n12812_, new_n12813_,
    new_n12814_, new_n12815_, new_n12816_, new_n12817_, new_n12818_,
    new_n12819_, new_n12820_, new_n12821_, new_n12822_, new_n12823_,
    new_n12824_, new_n12825_, new_n12826_, new_n12827_, new_n12828_,
    new_n12829_, new_n12830_, new_n12831_, new_n12832_, new_n12833_,
    new_n12834_, new_n12835_, new_n12836_, new_n12837_, new_n12838_,
    new_n12839_, new_n12840_, new_n12841_, new_n12842_, new_n12843_,
    new_n12844_, new_n12845_, new_n12846_, new_n12847_, new_n12848_,
    new_n12849_, new_n12850_, new_n12851_, new_n12852_, new_n12853_,
    new_n12854_, new_n12855_, new_n12856_, new_n12857_, new_n12858_,
    new_n12859_, new_n12860_, new_n12861_, new_n12862_, new_n12863_,
    new_n12864_, new_n12865_, new_n12866_, new_n12867_, new_n12868_,
    new_n12869_, new_n12870_, new_n12871_, new_n12872_, new_n12873_,
    new_n12874_, new_n12875_, new_n12876_, new_n12877_, new_n12878_,
    new_n12879_, new_n12880_, new_n12881_, new_n12882_, new_n12883_,
    new_n12884_, new_n12885_, new_n12886_, new_n12887_, new_n12888_,
    new_n12889_, new_n12890_, new_n12891_, new_n12892_, new_n12893_,
    new_n12894_, new_n12895_, new_n12896_, new_n12897_, new_n12898_,
    new_n12899_, new_n12900_, new_n12901_, new_n12902_, new_n12903_,
    new_n12904_, new_n12905_, new_n12906_, new_n12907_, new_n12908_,
    new_n12909_, new_n12910_, new_n12911_, new_n12912_, new_n12913_,
    new_n12914_, new_n12915_, new_n12916_, new_n12917_, new_n12918_,
    new_n12919_, new_n12920_, new_n12921_, new_n12922_, new_n12923_,
    new_n12924_, new_n12925_, new_n12926_, new_n12927_, new_n12928_,
    new_n12929_, new_n12930_, new_n12931_, new_n12932_, new_n12933_,
    new_n12934_, new_n12935_, new_n12936_, new_n12937_, new_n12938_,
    new_n12939_, new_n12940_, new_n12941_, new_n12942_, new_n12943_,
    new_n12944_, new_n12945_, new_n12946_, new_n12947_, new_n12948_,
    new_n12949_, new_n12950_, new_n12951_, new_n12952_, new_n12953_,
    new_n12954_, new_n12955_, new_n12956_, new_n12957_, new_n12958_,
    new_n12959_, new_n12960_, new_n12961_, new_n12962_, new_n12963_,
    new_n12964_, new_n12965_, new_n12966_, new_n12967_, new_n12968_,
    new_n12969_, new_n12970_, new_n12971_, new_n12972_, new_n12973_,
    new_n12974_, new_n12975_, new_n12976_, new_n12977_, new_n12978_,
    new_n12979_, new_n12980_, new_n12981_, new_n12982_, new_n12983_,
    new_n12984_, new_n12985_, new_n12986_, new_n12987_, new_n12988_,
    new_n12989_, new_n12990_, new_n12991_, new_n12992_, new_n12993_,
    new_n12994_, new_n12995_, new_n12996_, new_n12997_, new_n12998_,
    new_n12999_, new_n13000_, new_n13001_, new_n13002_, new_n13003_,
    new_n13004_, new_n13005_, new_n13006_, new_n13007_, new_n13008_,
    new_n13009_, new_n13010_, new_n13011_, new_n13012_, new_n13013_,
    new_n13014_, new_n13015_, new_n13016_, new_n13017_, new_n13018_,
    new_n13019_, new_n13020_, new_n13021_, new_n13022_, new_n13023_,
    new_n13024_, new_n13025_, new_n13026_, new_n13027_, new_n13028_,
    new_n13029_, new_n13030_, new_n13031_, new_n13032_, new_n13033_,
    new_n13034_, new_n13035_, new_n13036_, new_n13037_, new_n13038_,
    new_n13039_, new_n13040_, new_n13041_, new_n13042_, new_n13043_,
    new_n13044_, new_n13045_, new_n13046_, new_n13047_, new_n13048_,
    new_n13049_, new_n13050_, new_n13051_, new_n13052_, new_n13053_,
    new_n13054_, new_n13055_, new_n13056_, new_n13057_, new_n13058_,
    new_n13059_, new_n13060_, new_n13061_, new_n13062_, new_n13063_,
    new_n13064_, new_n13065_, new_n13066_, new_n13067_, new_n13068_,
    new_n13069_, new_n13070_, new_n13071_, new_n13072_, new_n13073_,
    new_n13074_, new_n13075_, new_n13076_, new_n13077_, new_n13078_,
    new_n13079_, new_n13080_, new_n13081_, new_n13082_, new_n13083_,
    new_n13084_, new_n13085_, new_n13086_, new_n13087_, new_n13088_,
    new_n13089_, new_n13090_, new_n13091_, new_n13092_, new_n13093_,
    new_n13094_, new_n13095_, new_n13096_, new_n13097_, new_n13098_,
    new_n13099_, new_n13100_, new_n13101_, new_n13102_, new_n13103_,
    new_n13104_, new_n13105_, new_n13106_, new_n13107_, new_n13108_,
    new_n13109_, new_n13110_, new_n13111_, new_n13112_, new_n13113_,
    new_n13114_, new_n13115_, new_n13116_, new_n13117_, new_n13118_,
    new_n13119_, new_n13120_, new_n13121_, new_n13122_, new_n13123_,
    new_n13124_, new_n13125_, new_n13126_, new_n13127_, new_n13128_,
    new_n13129_, new_n13130_, new_n13131_, new_n13132_, new_n13133_,
    new_n13134_, new_n13135_, new_n13136_, new_n13137_, new_n13138_,
    new_n13139_, new_n13140_, new_n13141_, new_n13142_, new_n13143_,
    new_n13144_, new_n13145_, new_n13146_, new_n13147_, new_n13148_,
    new_n13149_, new_n13150_, new_n13151_, new_n13152_, new_n13153_,
    new_n13154_, new_n13155_, new_n13156_, new_n13157_, new_n13158_,
    new_n13159_, new_n13160_, new_n13161_, new_n13162_, new_n13163_,
    new_n13164_, new_n13165_, new_n13166_, new_n13167_, new_n13168_,
    new_n13169_, new_n13170_, new_n13171_, new_n13172_, new_n13173_,
    new_n13174_, new_n13175_, new_n13176_, new_n13177_, new_n13178_,
    new_n13179_, new_n13180_, new_n13181_, new_n13182_, new_n13183_,
    new_n13184_, new_n13185_, new_n13186_, new_n13187_, new_n13188_,
    new_n13189_, new_n13190_, new_n13191_, new_n13192_, new_n13193_,
    new_n13194_, new_n13195_, new_n13196_, new_n13197_, new_n13198_,
    new_n13199_, new_n13200_, new_n13201_, new_n13202_, new_n13203_,
    new_n13204_, new_n13205_, new_n13206_, new_n13207_, new_n13208_,
    new_n13209_, new_n13210_, new_n13211_, new_n13212_, new_n13213_,
    new_n13214_, new_n13215_, new_n13216_, new_n13217_, new_n13218_,
    new_n13219_, new_n13220_, new_n13221_, new_n13222_, new_n13223_,
    new_n13224_, new_n13225_, new_n13226_, new_n13227_, new_n13228_,
    new_n13229_, new_n13230_, new_n13231_, new_n13232_, new_n13233_,
    new_n13234_, new_n13235_, new_n13236_, new_n13237_, new_n13238_,
    new_n13239_, new_n13240_, new_n13241_, new_n13242_, new_n13243_,
    new_n13244_, new_n13245_, new_n13246_, new_n13247_, new_n13248_,
    new_n13249_, new_n13250_, new_n13251_, new_n13252_, new_n13253_,
    new_n13254_, new_n13255_, new_n13256_, new_n13257_, new_n13258_,
    new_n13259_, new_n13260_, new_n13261_, new_n13262_, new_n13263_,
    new_n13264_, new_n13265_, new_n13266_, new_n13267_, new_n13268_,
    new_n13269_, new_n13270_, new_n13271_, new_n13272_, new_n13273_,
    new_n13274_, new_n13275_, new_n13276_, new_n13277_, new_n13278_,
    new_n13279_, new_n13280_, new_n13281_, new_n13282_, new_n13283_,
    new_n13284_, new_n13285_, new_n13286_, new_n13287_, new_n13288_,
    new_n13289_, new_n13290_, new_n13291_, new_n13292_, new_n13293_,
    new_n13294_, new_n13295_, new_n13296_, new_n13297_, new_n13298_,
    new_n13299_, new_n13300_, new_n13301_, new_n13302_, new_n13303_,
    new_n13304_, new_n13305_, new_n13306_, new_n13307_, new_n13308_,
    new_n13309_, new_n13310_, new_n13311_, new_n13312_, new_n13313_,
    new_n13314_, new_n13315_, new_n13316_, new_n13317_, new_n13318_,
    new_n13319_, new_n13320_, new_n13321_, new_n13322_, new_n13323_,
    new_n13324_, new_n13325_, new_n13326_, new_n13327_, new_n13328_,
    new_n13329_, new_n13330_, new_n13331_, new_n13332_, new_n13333_,
    new_n13334_, new_n13335_, new_n13336_, new_n13337_, new_n13338_,
    new_n13339_, new_n13340_, new_n13341_, new_n13342_, new_n13343_,
    new_n13344_, new_n13345_, new_n13346_, new_n13347_, new_n13348_,
    new_n13349_, new_n13350_, new_n13351_, new_n13352_, new_n13353_,
    new_n13354_, new_n13355_, new_n13357_, new_n13358_, new_n13359_,
    new_n13360_, new_n13361_, new_n13362_, new_n13363_, new_n13364_,
    new_n13365_, new_n13366_, new_n13367_, new_n13368_, new_n13369_,
    new_n13370_, new_n13371_, new_n13372_, new_n13373_, new_n13374_,
    new_n13375_, new_n13376_, new_n13377_, new_n13378_, new_n13379_,
    new_n13380_, new_n13381_, new_n13382_, new_n13383_, new_n13384_,
    new_n13385_, new_n13386_, new_n13387_, new_n13388_, new_n13389_,
    new_n13390_, new_n13391_, new_n13392_, new_n13393_, new_n13394_,
    new_n13395_, new_n13396_, new_n13397_, new_n13398_, new_n13399_,
    new_n13400_, new_n13401_, new_n13402_, new_n13403_, new_n13404_,
    new_n13405_, new_n13406_, new_n13407_, new_n13408_, new_n13409_,
    new_n13410_, new_n13411_, new_n13412_, new_n13413_, new_n13414_,
    new_n13415_, new_n13416_, new_n13417_, new_n13418_, new_n13419_,
    new_n13420_, new_n13421_, new_n13422_, new_n13423_, new_n13424_,
    new_n13425_, new_n13426_, new_n13427_, new_n13428_, new_n13429_,
    new_n13430_, new_n13431_, new_n13432_, new_n13433_, new_n13434_,
    new_n13435_, new_n13436_, new_n13437_, new_n13438_, new_n13439_,
    new_n13440_, new_n13441_, new_n13442_, new_n13443_, new_n13444_,
    new_n13445_, new_n13446_, new_n13447_, new_n13448_, new_n13449_,
    new_n13450_, new_n13451_, new_n13452_, new_n13453_, new_n13454_,
    new_n13455_, new_n13456_, new_n13457_, new_n13458_, new_n13459_,
    new_n13460_, new_n13461_, new_n13462_, new_n13463_, new_n13464_,
    new_n13465_, new_n13466_, new_n13467_, new_n13468_, new_n13469_,
    new_n13470_, new_n13471_, new_n13472_, new_n13473_, new_n13474_,
    new_n13475_, new_n13476_, new_n13477_, new_n13478_, new_n13479_,
    new_n13480_, new_n13481_, new_n13482_, new_n13483_, new_n13484_,
    new_n13485_, new_n13486_, new_n13487_, new_n13488_, new_n13489_,
    new_n13490_, new_n13491_, new_n13492_, new_n13493_, new_n13494_,
    new_n13495_, new_n13496_, new_n13497_, new_n13498_, new_n13499_,
    new_n13500_, new_n13501_, new_n13502_, new_n13503_, new_n13504_,
    new_n13505_, new_n13506_, new_n13507_, new_n13508_, new_n13509_,
    new_n13510_, new_n13511_, new_n13512_, new_n13513_, new_n13514_,
    new_n13515_, new_n13516_, new_n13517_, new_n13518_, new_n13519_,
    new_n13520_, new_n13521_, new_n13522_, new_n13523_, new_n13524_,
    new_n13525_, new_n13526_, new_n13527_, new_n13528_, new_n13529_,
    new_n13530_, new_n13531_, new_n13532_, new_n13533_, new_n13534_,
    new_n13535_, new_n13536_, new_n13537_, new_n13538_, new_n13539_,
    new_n13540_, new_n13541_, new_n13542_, new_n13543_, new_n13544_,
    new_n13545_, new_n13546_, new_n13547_, new_n13548_, new_n13549_,
    new_n13550_, new_n13551_, new_n13552_, new_n13553_, new_n13554_,
    new_n13555_, new_n13556_, new_n13557_, new_n13558_, new_n13559_,
    new_n13560_, new_n13561_, new_n13562_, new_n13563_, new_n13564_,
    new_n13565_, new_n13566_, new_n13567_, new_n13568_, new_n13569_,
    new_n13570_, new_n13571_, new_n13572_, new_n13573_, new_n13574_,
    new_n13575_, new_n13576_, new_n13577_, new_n13578_, new_n13579_,
    new_n13580_, new_n13581_, new_n13582_, new_n13583_, new_n13584_,
    new_n13585_, new_n13586_, new_n13587_, new_n13588_, new_n13589_,
    new_n13590_, new_n13591_, new_n13592_, new_n13593_, new_n13594_,
    new_n13595_, new_n13596_, new_n13597_, new_n13598_, new_n13599_,
    new_n13600_, new_n13601_, new_n13602_, new_n13603_, new_n13604_,
    new_n13605_, new_n13606_, new_n13607_, new_n13608_, new_n13609_,
    new_n13610_, new_n13611_, new_n13612_, new_n13613_, new_n13614_,
    new_n13615_, new_n13616_, new_n13617_, new_n13618_, new_n13619_,
    new_n13620_, new_n13621_, new_n13622_, new_n13623_, new_n13624_,
    new_n13625_, new_n13626_, new_n13627_, new_n13628_, new_n13629_,
    new_n13630_, new_n13631_, new_n13632_, new_n13633_, new_n13634_,
    new_n13635_, new_n13636_, new_n13637_, new_n13638_, new_n13639_,
    new_n13640_, new_n13641_, new_n13642_, new_n13643_, new_n13644_,
    new_n13645_, new_n13646_, new_n13647_, new_n13648_, new_n13649_,
    new_n13650_, new_n13651_, new_n13652_, new_n13653_, new_n13654_,
    new_n13655_, new_n13656_, new_n13657_, new_n13658_, new_n13659_,
    new_n13660_, new_n13661_, new_n13662_, new_n13663_, new_n13664_,
    new_n13665_, new_n13666_, new_n13667_, new_n13668_, new_n13669_,
    new_n13670_, new_n13671_, new_n13672_, new_n13673_, new_n13674_,
    new_n13675_, new_n13676_, new_n13677_, new_n13678_, new_n13679_,
    new_n13680_, new_n13681_, new_n13682_, new_n13683_, new_n13684_,
    new_n13685_, new_n13686_, new_n13687_, new_n13688_, new_n13689_,
    new_n13690_, new_n13691_, new_n13692_, new_n13693_, new_n13694_,
    new_n13695_, new_n13696_, new_n13697_, new_n13698_, new_n13699_,
    new_n13700_, new_n13701_, new_n13702_, new_n13703_, new_n13704_,
    new_n13705_, new_n13706_, new_n13707_, new_n13708_, new_n13709_,
    new_n13710_, new_n13711_, new_n13712_, new_n13713_, new_n13714_,
    new_n13715_, new_n13716_, new_n13717_, new_n13718_, new_n13719_,
    new_n13720_, new_n13721_, new_n13722_, new_n13723_, new_n13724_,
    new_n13725_, new_n13726_, new_n13727_, new_n13728_, new_n13729_,
    new_n13730_, new_n13731_, new_n13732_, new_n13733_, new_n13734_,
    new_n13735_, new_n13736_, new_n13737_, new_n13738_, new_n13739_,
    new_n13740_, new_n13741_, new_n13742_, new_n13743_, new_n13744_,
    new_n13745_, new_n13746_, new_n13747_, new_n13748_, new_n13749_,
    new_n13750_, new_n13751_, new_n13752_, new_n13753_, new_n13754_,
    new_n13755_, new_n13756_, new_n13757_, new_n13758_, new_n13759_,
    new_n13760_, new_n13761_, new_n13762_, new_n13763_, new_n13764_,
    new_n13765_, new_n13766_, new_n13767_, new_n13768_, new_n13769_,
    new_n13770_, new_n13771_, new_n13772_, new_n13773_, new_n13774_,
    new_n13775_, new_n13776_, new_n13777_, new_n13778_, new_n13779_,
    new_n13780_, new_n13781_, new_n13782_, new_n13783_, new_n13784_,
    new_n13785_, new_n13786_, new_n13787_, new_n13788_, new_n13789_,
    new_n13790_, new_n13791_, new_n13792_, new_n13793_, new_n13794_,
    new_n13795_, new_n13796_, new_n13797_, new_n13798_, new_n13799_,
    new_n13800_, new_n13801_, new_n13802_, new_n13803_, new_n13804_,
    new_n13805_, new_n13806_, new_n13807_, new_n13808_, new_n13809_,
    new_n13810_, new_n13811_, new_n13812_, new_n13813_, new_n13814_,
    new_n13815_, new_n13816_, new_n13817_, new_n13818_, new_n13819_,
    new_n13820_, new_n13821_, new_n13822_, new_n13823_, new_n13824_,
    new_n13825_, new_n13826_, new_n13827_, new_n13828_, new_n13829_,
    new_n13830_, new_n13831_, new_n13832_, new_n13833_, new_n13834_,
    new_n13835_, new_n13836_, new_n13837_, new_n13838_, new_n13839_,
    new_n13840_, new_n13841_, new_n13842_, new_n13843_, new_n13844_,
    new_n13845_, new_n13846_, new_n13847_, new_n13848_, new_n13849_,
    new_n13850_, new_n13851_, new_n13852_, new_n13853_, new_n13854_,
    new_n13855_, new_n13856_, new_n13857_, new_n13858_, new_n13859_,
    new_n13860_, new_n13861_, new_n13862_, new_n13863_, new_n13864_,
    new_n13865_, new_n13866_, new_n13867_, new_n13868_, new_n13869_,
    new_n13870_, new_n13871_, new_n13872_, new_n13873_, new_n13874_,
    new_n13875_, new_n13876_, new_n13877_, new_n13878_, new_n13879_,
    new_n13880_, new_n13881_, new_n13882_, new_n13883_, new_n13884_,
    new_n13885_, new_n13886_, new_n13887_, new_n13888_, new_n13889_,
    new_n13890_, new_n13891_, new_n13892_, new_n13893_, new_n13894_,
    new_n13895_, new_n13896_, new_n13897_, new_n13898_, new_n13899_,
    new_n13900_, new_n13901_, new_n13902_, new_n13903_, new_n13904_,
    new_n13905_, new_n13906_, new_n13907_, new_n13908_, new_n13909_,
    new_n13910_, new_n13911_, new_n13912_, new_n13913_, new_n13914_,
    new_n13915_, new_n13916_, new_n13917_, new_n13918_, new_n13919_,
    new_n13920_, new_n13921_, new_n13922_, new_n13923_, new_n13924_,
    new_n13925_, new_n13926_, new_n13927_, new_n13928_, new_n13929_,
    new_n13930_, new_n13931_, new_n13932_, new_n13933_, new_n13934_,
    new_n13935_, new_n13936_, new_n13937_, new_n13938_, new_n13939_,
    new_n13940_, new_n13941_, new_n13942_, new_n13943_, new_n13944_,
    new_n13945_, new_n13946_, new_n13947_, new_n13948_, new_n13949_,
    new_n13950_, new_n13951_, new_n13952_, new_n13953_, new_n13954_,
    new_n13955_, new_n13956_, new_n13957_, new_n13958_, new_n13959_,
    new_n13960_, new_n13961_, new_n13962_, new_n13964_, new_n13965_,
    new_n13966_, new_n13967_, new_n13968_, new_n13969_, new_n13970_,
    new_n13971_, new_n13972_, new_n13973_, new_n13974_, new_n13975_,
    new_n13976_, new_n13977_, new_n13978_, new_n13979_, new_n13980_,
    new_n13981_, new_n13982_, new_n13983_, new_n13984_, new_n13985_,
    new_n13986_, new_n13987_, new_n13988_, new_n13989_, new_n13990_,
    new_n13991_, new_n13992_, new_n13993_, new_n13994_, new_n13995_,
    new_n13996_, new_n13997_, new_n13998_, new_n13999_, new_n14000_,
    new_n14001_, new_n14002_, new_n14003_, new_n14004_, new_n14005_,
    new_n14006_, new_n14007_, new_n14008_, new_n14009_, new_n14010_,
    new_n14011_, new_n14012_, new_n14013_, new_n14014_, new_n14015_,
    new_n14016_, new_n14017_, new_n14018_, new_n14019_, new_n14020_,
    new_n14021_, new_n14022_, new_n14023_, new_n14024_, new_n14025_,
    new_n14026_, new_n14027_, new_n14028_, new_n14029_, new_n14030_,
    new_n14031_, new_n14032_, new_n14033_, new_n14034_, new_n14035_,
    new_n14036_, new_n14037_, new_n14038_, new_n14039_, new_n14040_,
    new_n14041_, new_n14042_, new_n14043_, new_n14044_, new_n14045_,
    new_n14046_, new_n14047_, new_n14048_, new_n14049_, new_n14050_,
    new_n14051_, new_n14052_, new_n14053_, new_n14054_, new_n14055_,
    new_n14056_, new_n14057_, new_n14058_, new_n14059_, new_n14060_,
    new_n14061_, new_n14062_, new_n14063_, new_n14064_, new_n14065_,
    new_n14066_, new_n14067_, new_n14068_, new_n14069_, new_n14070_,
    new_n14071_, new_n14072_, new_n14073_, new_n14074_, new_n14075_,
    new_n14076_, new_n14077_, new_n14078_, new_n14079_, new_n14080_,
    new_n14081_, new_n14082_, new_n14083_, new_n14084_, new_n14085_,
    new_n14086_, new_n14087_, new_n14088_, new_n14089_, new_n14090_,
    new_n14091_, new_n14092_, new_n14093_, new_n14094_, new_n14095_,
    new_n14096_, new_n14097_, new_n14098_, new_n14099_, new_n14100_,
    new_n14101_, new_n14102_, new_n14103_, new_n14104_, new_n14105_,
    new_n14106_, new_n14107_, new_n14108_, new_n14109_, new_n14110_,
    new_n14111_, new_n14112_, new_n14113_, new_n14114_, new_n14115_,
    new_n14116_, new_n14117_, new_n14118_, new_n14119_, new_n14120_,
    new_n14121_, new_n14122_, new_n14123_, new_n14124_, new_n14125_,
    new_n14126_, new_n14127_, new_n14128_, new_n14129_, new_n14130_,
    new_n14131_, new_n14132_, new_n14133_, new_n14134_, new_n14135_,
    new_n14136_, new_n14137_, new_n14138_, new_n14139_, new_n14140_,
    new_n14141_, new_n14142_, new_n14143_, new_n14144_, new_n14145_,
    new_n14146_, new_n14147_, new_n14148_, new_n14149_, new_n14150_,
    new_n14151_, new_n14152_, new_n14153_, new_n14154_, new_n14155_,
    new_n14156_, new_n14157_, new_n14158_, new_n14159_, new_n14160_,
    new_n14161_, new_n14162_, new_n14163_, new_n14164_, new_n14165_,
    new_n14166_, new_n14167_, new_n14168_, new_n14169_, new_n14170_,
    new_n14171_, new_n14172_, new_n14173_, new_n14174_, new_n14175_,
    new_n14176_, new_n14177_, new_n14178_, new_n14179_, new_n14180_,
    new_n14181_, new_n14182_, new_n14183_, new_n14184_, new_n14185_,
    new_n14186_, new_n14187_, new_n14188_, new_n14189_, new_n14190_,
    new_n14191_, new_n14192_, new_n14193_, new_n14194_, new_n14195_,
    new_n14196_, new_n14197_, new_n14198_, new_n14199_, new_n14200_,
    new_n14201_, new_n14202_, new_n14203_, new_n14204_, new_n14205_,
    new_n14206_, new_n14207_, new_n14208_, new_n14209_, new_n14210_,
    new_n14211_, new_n14212_, new_n14213_, new_n14214_, new_n14215_,
    new_n14216_, new_n14217_, new_n14218_, new_n14219_, new_n14220_,
    new_n14221_, new_n14222_, new_n14223_, new_n14224_, new_n14225_,
    new_n14226_, new_n14227_, new_n14228_, new_n14229_, new_n14230_,
    new_n14231_, new_n14232_, new_n14233_, new_n14234_, new_n14235_,
    new_n14236_, new_n14237_, new_n14238_, new_n14239_, new_n14240_,
    new_n14241_, new_n14242_, new_n14243_, new_n14244_, new_n14245_,
    new_n14246_, new_n14247_, new_n14248_, new_n14249_, new_n14250_,
    new_n14251_, new_n14252_, new_n14253_, new_n14254_, new_n14255_,
    new_n14256_, new_n14257_, new_n14258_, new_n14259_, new_n14260_,
    new_n14261_, new_n14262_, new_n14263_, new_n14264_, new_n14265_,
    new_n14266_, new_n14267_, new_n14268_, new_n14269_, new_n14270_,
    new_n14271_, new_n14272_, new_n14273_, new_n14274_, new_n14275_,
    new_n14276_, new_n14277_, new_n14278_, new_n14279_, new_n14280_,
    new_n14281_, new_n14282_, new_n14283_, new_n14284_, new_n14285_,
    new_n14286_, new_n14287_, new_n14288_, new_n14289_, new_n14290_,
    new_n14291_, new_n14292_, new_n14293_, new_n14294_, new_n14295_,
    new_n14296_, new_n14297_, new_n14298_, new_n14299_, new_n14300_,
    new_n14301_, new_n14302_, new_n14303_, new_n14304_, new_n14305_,
    new_n14306_, new_n14307_, new_n14308_, new_n14309_, new_n14310_,
    new_n14311_, new_n14312_, new_n14313_, new_n14314_, new_n14315_,
    new_n14316_, new_n14317_, new_n14318_, new_n14319_, new_n14320_,
    new_n14321_, new_n14322_, new_n14323_, new_n14324_, new_n14325_,
    new_n14326_, new_n14327_, new_n14328_, new_n14329_, new_n14330_,
    new_n14331_, new_n14332_, new_n14333_, new_n14334_, new_n14335_,
    new_n14336_, new_n14337_, new_n14338_, new_n14339_, new_n14340_,
    new_n14341_, new_n14342_, new_n14343_, new_n14344_, new_n14345_,
    new_n14346_, new_n14347_, new_n14348_, new_n14349_, new_n14350_,
    new_n14351_, new_n14352_, new_n14353_, new_n14354_, new_n14355_,
    new_n14356_, new_n14357_, new_n14358_, new_n14359_, new_n14360_,
    new_n14361_, new_n14362_, new_n14363_, new_n14364_, new_n14365_,
    new_n14366_, new_n14367_, new_n14368_, new_n14369_, new_n14370_,
    new_n14371_, new_n14372_, new_n14373_, new_n14374_, new_n14375_,
    new_n14376_, new_n14377_, new_n14378_, new_n14379_, new_n14380_,
    new_n14381_, new_n14382_, new_n14383_, new_n14384_, new_n14385_,
    new_n14386_, new_n14387_, new_n14388_, new_n14389_, new_n14390_,
    new_n14391_, new_n14392_, new_n14393_, new_n14394_, new_n14395_,
    new_n14396_, new_n14397_, new_n14398_, new_n14399_, new_n14400_,
    new_n14401_, new_n14402_, new_n14403_, new_n14404_, new_n14405_,
    new_n14406_, new_n14407_, new_n14408_, new_n14409_, new_n14410_,
    new_n14411_, new_n14412_, new_n14413_, new_n14414_, new_n14415_,
    new_n14416_, new_n14417_, new_n14418_, new_n14419_, new_n14420_,
    new_n14421_, new_n14422_, new_n14423_, new_n14424_, new_n14425_,
    new_n14426_, new_n14427_, new_n14428_, new_n14429_, new_n14430_,
    new_n14431_, new_n14432_, new_n14433_, new_n14434_, new_n14435_,
    new_n14436_, new_n14437_, new_n14438_, new_n14439_, new_n14440_,
    new_n14441_, new_n14442_, new_n14443_, new_n14444_, new_n14445_,
    new_n14446_, new_n14447_, new_n14448_, new_n14449_, new_n14450_,
    new_n14451_, new_n14452_, new_n14453_, new_n14454_, new_n14455_,
    new_n14456_, new_n14457_, new_n14458_, new_n14459_, new_n14460_,
    new_n14461_, new_n14462_, new_n14463_, new_n14464_, new_n14465_,
    new_n14466_, new_n14467_, new_n14468_, new_n14469_, new_n14470_,
    new_n14471_, new_n14472_, new_n14473_, new_n14474_, new_n14475_,
    new_n14476_, new_n14477_, new_n14478_, new_n14479_, new_n14480_,
    new_n14481_, new_n14482_, new_n14483_, new_n14484_, new_n14485_,
    new_n14486_, new_n14487_, new_n14488_, new_n14489_, new_n14490_,
    new_n14491_, new_n14492_, new_n14493_, new_n14494_, new_n14495_,
    new_n14496_, new_n14497_, new_n14498_, new_n14499_, new_n14500_,
    new_n14501_, new_n14502_, new_n14503_, new_n14504_, new_n14505_,
    new_n14506_, new_n14507_, new_n14508_, new_n14509_, new_n14510_,
    new_n14511_, new_n14512_, new_n14513_, new_n14514_, new_n14515_,
    new_n14516_, new_n14517_, new_n14518_, new_n14519_, new_n14520_,
    new_n14521_, new_n14522_, new_n14523_, new_n14524_, new_n14525_,
    new_n14526_, new_n14527_, new_n14528_, new_n14529_, new_n14530_,
    new_n14531_, new_n14532_, new_n14533_, new_n14534_, new_n14535_,
    new_n14536_, new_n14537_, new_n14538_, new_n14539_, new_n14540_,
    new_n14541_, new_n14542_, new_n14543_, new_n14544_, new_n14545_,
    new_n14546_, new_n14547_, new_n14548_, new_n14549_, new_n14550_,
    new_n14551_, new_n14552_, new_n14553_, new_n14554_, new_n14555_,
    new_n14556_, new_n14557_, new_n14558_, new_n14559_, new_n14560_,
    new_n14561_, new_n14562_, new_n14563_, new_n14564_, new_n14565_,
    new_n14566_, new_n14567_, new_n14568_, new_n14569_, new_n14570_,
    new_n14571_, new_n14572_, new_n14573_, new_n14574_, new_n14575_,
    new_n14576_, new_n14577_, new_n14578_, new_n14579_, new_n14580_,
    new_n14582_, new_n14583_, new_n14584_, new_n14585_, new_n14586_,
    new_n14587_, new_n14588_, new_n14589_, new_n14590_, new_n14591_,
    new_n14592_, new_n14593_, new_n14594_, new_n14595_, new_n14596_,
    new_n14597_, new_n14598_, new_n14599_, new_n14600_, new_n14601_,
    new_n14602_, new_n14603_, new_n14604_, new_n14605_, new_n14606_,
    new_n14607_, new_n14608_, new_n14609_, new_n14610_, new_n14611_,
    new_n14612_, new_n14613_, new_n14614_, new_n14615_, new_n14616_,
    new_n14617_, new_n14618_, new_n14619_, new_n14620_, new_n14621_,
    new_n14622_, new_n14623_, new_n14624_, new_n14625_, new_n14626_,
    new_n14627_, new_n14628_, new_n14629_, new_n14630_, new_n14631_,
    new_n14632_, new_n14633_, new_n14634_, new_n14635_, new_n14636_,
    new_n14637_, new_n14638_, new_n14639_, new_n14640_, new_n14641_,
    new_n14642_, new_n14643_, new_n14644_, new_n14645_, new_n14646_,
    new_n14647_, new_n14648_, new_n14649_, new_n14650_, new_n14651_,
    new_n14652_, new_n14653_, new_n14654_, new_n14655_, new_n14656_,
    new_n14657_, new_n14658_, new_n14659_, new_n14660_, new_n14661_,
    new_n14662_, new_n14663_, new_n14664_, new_n14665_, new_n14666_,
    new_n14667_, new_n14668_, new_n14669_, new_n14670_, new_n14671_,
    new_n14672_, new_n14673_, new_n14674_, new_n14675_, new_n14676_,
    new_n14677_, new_n14678_, new_n14679_, new_n14680_, new_n14681_,
    new_n14682_, new_n14683_, new_n14684_, new_n14685_, new_n14686_,
    new_n14687_, new_n14688_, new_n14689_, new_n14690_, new_n14691_,
    new_n14692_, new_n14693_, new_n14694_, new_n14695_, new_n14696_,
    new_n14697_, new_n14698_, new_n14699_, new_n14700_, new_n14701_,
    new_n14702_, new_n14703_, new_n14704_, new_n14705_, new_n14706_,
    new_n14707_, new_n14708_, new_n14709_, new_n14710_, new_n14711_,
    new_n14712_, new_n14713_, new_n14714_, new_n14715_, new_n14716_,
    new_n14717_, new_n14718_, new_n14719_, new_n14720_, new_n14721_,
    new_n14722_, new_n14723_, new_n14724_, new_n14725_, new_n14726_,
    new_n14727_, new_n14728_, new_n14729_, new_n14730_, new_n14731_,
    new_n14732_, new_n14733_, new_n14734_, new_n14735_, new_n14736_,
    new_n14737_, new_n14738_, new_n14739_, new_n14740_, new_n14741_,
    new_n14742_, new_n14743_, new_n14744_, new_n14745_, new_n14746_,
    new_n14747_, new_n14748_, new_n14749_, new_n14750_, new_n14751_,
    new_n14752_, new_n14753_, new_n14754_, new_n14755_, new_n14756_,
    new_n14757_, new_n14758_, new_n14759_, new_n14760_, new_n14761_,
    new_n14762_, new_n14763_, new_n14764_, new_n14765_, new_n14766_,
    new_n14767_, new_n14768_, new_n14769_, new_n14770_, new_n14771_,
    new_n14772_, new_n14773_, new_n14774_, new_n14775_, new_n14776_,
    new_n14777_, new_n14778_, new_n14779_, new_n14780_, new_n14781_,
    new_n14782_, new_n14783_, new_n14784_, new_n14785_, new_n14786_,
    new_n14787_, new_n14788_, new_n14789_, new_n14790_, new_n14791_,
    new_n14792_, new_n14793_, new_n14794_, new_n14795_, new_n14796_,
    new_n14797_, new_n14798_, new_n14799_, new_n14800_, new_n14801_,
    new_n14802_, new_n14803_, new_n14804_, new_n14805_, new_n14806_,
    new_n14807_, new_n14808_, new_n14809_, new_n14810_, new_n14811_,
    new_n14812_, new_n14813_, new_n14814_, new_n14815_, new_n14816_,
    new_n14817_, new_n14818_, new_n14819_, new_n14820_, new_n14821_,
    new_n14822_, new_n14823_, new_n14824_, new_n14825_, new_n14826_,
    new_n14827_, new_n14828_, new_n14829_, new_n14830_, new_n14831_,
    new_n14832_, new_n14833_, new_n14834_, new_n14835_, new_n14836_,
    new_n14837_, new_n14838_, new_n14839_, new_n14840_, new_n14841_,
    new_n14842_, new_n14843_, new_n14844_, new_n14845_, new_n14846_,
    new_n14847_, new_n14848_, new_n14849_, new_n14850_, new_n14851_,
    new_n14852_, new_n14853_, new_n14854_, new_n14855_, new_n14856_,
    new_n14857_, new_n14858_, new_n14859_, new_n14860_, new_n14861_,
    new_n14862_, new_n14863_, new_n14864_, new_n14865_, new_n14866_,
    new_n14867_, new_n14868_, new_n14869_, new_n14870_, new_n14871_,
    new_n14872_, new_n14873_, new_n14874_, new_n14875_, new_n14876_,
    new_n14877_, new_n14878_, new_n14879_, new_n14880_, new_n14881_,
    new_n14882_, new_n14883_, new_n14884_, new_n14885_, new_n14886_,
    new_n14887_, new_n14888_, new_n14889_, new_n14890_, new_n14891_,
    new_n14892_, new_n14893_, new_n14894_, new_n14895_, new_n14896_,
    new_n14897_, new_n14898_, new_n14899_, new_n14900_, new_n14901_,
    new_n14902_, new_n14903_, new_n14904_, new_n14905_, new_n14906_,
    new_n14907_, new_n14908_, new_n14909_, new_n14910_, new_n14911_,
    new_n14912_, new_n14913_, new_n14914_, new_n14915_, new_n14916_,
    new_n14917_, new_n14918_, new_n14919_, new_n14920_, new_n14921_,
    new_n14922_, new_n14923_, new_n14924_, new_n14925_, new_n14926_,
    new_n14927_, new_n14928_, new_n14929_, new_n14930_, new_n14931_,
    new_n14932_, new_n14933_, new_n14934_, new_n14935_, new_n14936_,
    new_n14937_, new_n14938_, new_n14939_, new_n14940_, new_n14941_,
    new_n14942_, new_n14943_, new_n14944_, new_n14945_, new_n14946_,
    new_n14947_, new_n14948_, new_n14949_, new_n14950_, new_n14951_,
    new_n14952_, new_n14953_, new_n14954_, new_n14955_, new_n14956_,
    new_n14957_, new_n14958_, new_n14959_, new_n14960_, new_n14961_,
    new_n14962_, new_n14963_, new_n14964_, new_n14965_, new_n14966_,
    new_n14967_, new_n14968_, new_n14969_, new_n14970_, new_n14971_,
    new_n14972_, new_n14973_, new_n14974_, new_n14975_, new_n14976_,
    new_n14977_, new_n14978_, new_n14979_, new_n14980_, new_n14981_,
    new_n14982_, new_n14983_, new_n14984_, new_n14985_, new_n14986_,
    new_n14987_, new_n14988_, new_n14989_, new_n14990_, new_n14991_,
    new_n14992_, new_n14993_, new_n14994_, new_n14995_, new_n14996_,
    new_n14997_, new_n14998_, new_n14999_, new_n15000_, new_n15001_,
    new_n15002_, new_n15003_, new_n15004_, new_n15005_, new_n15006_,
    new_n15007_, new_n15008_, new_n15009_, new_n15010_, new_n15011_,
    new_n15012_, new_n15013_, new_n15014_, new_n15015_, new_n15016_,
    new_n15017_, new_n15018_, new_n15019_, new_n15020_, new_n15021_,
    new_n15022_, new_n15023_, new_n15024_, new_n15025_, new_n15026_,
    new_n15027_, new_n15028_, new_n15029_, new_n15030_, new_n15031_,
    new_n15032_, new_n15033_, new_n15034_, new_n15035_, new_n15036_,
    new_n15037_, new_n15038_, new_n15039_, new_n15040_, new_n15041_,
    new_n15042_, new_n15043_, new_n15044_, new_n15045_, new_n15046_,
    new_n15047_, new_n15048_, new_n15049_, new_n15050_, new_n15051_,
    new_n15052_, new_n15053_, new_n15054_, new_n15055_, new_n15056_,
    new_n15057_, new_n15058_, new_n15059_, new_n15060_, new_n15061_,
    new_n15062_, new_n15063_, new_n15064_, new_n15065_, new_n15066_,
    new_n15067_, new_n15068_, new_n15069_, new_n15070_, new_n15071_,
    new_n15072_, new_n15073_, new_n15074_, new_n15075_, new_n15076_,
    new_n15077_, new_n15078_, new_n15079_, new_n15080_, new_n15081_,
    new_n15082_, new_n15083_, new_n15084_, new_n15085_, new_n15086_,
    new_n15087_, new_n15088_, new_n15089_, new_n15090_, new_n15091_,
    new_n15092_, new_n15093_, new_n15094_, new_n15095_, new_n15096_,
    new_n15097_, new_n15098_, new_n15099_, new_n15100_, new_n15101_,
    new_n15102_, new_n15103_, new_n15104_, new_n15105_, new_n15106_,
    new_n15107_, new_n15108_, new_n15109_, new_n15110_, new_n15111_,
    new_n15112_, new_n15113_, new_n15114_, new_n15115_, new_n15116_,
    new_n15117_, new_n15118_, new_n15119_, new_n15120_, new_n15121_,
    new_n15122_, new_n15123_, new_n15124_, new_n15125_, new_n15126_,
    new_n15127_, new_n15128_, new_n15129_, new_n15130_, new_n15131_,
    new_n15132_, new_n15133_, new_n15134_, new_n15135_, new_n15136_,
    new_n15137_, new_n15138_, new_n15139_, new_n15140_, new_n15141_,
    new_n15142_, new_n15143_, new_n15144_, new_n15145_, new_n15146_,
    new_n15147_, new_n15148_, new_n15149_, new_n15150_, new_n15151_,
    new_n15152_, new_n15153_, new_n15154_, new_n15155_, new_n15156_,
    new_n15157_, new_n15158_, new_n15159_, new_n15160_, new_n15161_,
    new_n15162_, new_n15163_, new_n15164_, new_n15165_, new_n15166_,
    new_n15167_, new_n15168_, new_n15169_, new_n15170_, new_n15171_,
    new_n15172_, new_n15173_, new_n15174_, new_n15175_, new_n15176_,
    new_n15177_, new_n15178_, new_n15179_, new_n15180_, new_n15181_,
    new_n15182_, new_n15183_, new_n15184_, new_n15185_, new_n15186_,
    new_n15187_, new_n15188_, new_n15189_, new_n15190_, new_n15191_,
    new_n15192_, new_n15193_, new_n15194_, new_n15195_, new_n15196_,
    new_n15197_, new_n15198_, new_n15199_, new_n15200_, new_n15201_,
    new_n15202_, new_n15203_, new_n15204_, new_n15205_, new_n15206_,
    new_n15207_, new_n15208_, new_n15209_, new_n15210_, new_n15211_,
    new_n15212_, new_n15214_, new_n15215_, new_n15216_, new_n15217_,
    new_n15218_, new_n15219_, new_n15220_, new_n15221_, new_n15222_,
    new_n15223_, new_n15224_, new_n15225_, new_n15226_, new_n15227_,
    new_n15228_, new_n15229_, new_n15230_, new_n15231_, new_n15232_,
    new_n15233_, new_n15234_, new_n15235_, new_n15236_, new_n15237_,
    new_n15238_, new_n15239_, new_n15240_, new_n15241_, new_n15242_,
    new_n15243_, new_n15244_, new_n15245_, new_n15246_, new_n15247_,
    new_n15248_, new_n15249_, new_n15250_, new_n15251_, new_n15252_,
    new_n15253_, new_n15254_, new_n15255_, new_n15256_, new_n15257_,
    new_n15258_, new_n15259_, new_n15260_, new_n15261_, new_n15262_,
    new_n15263_, new_n15264_, new_n15265_, new_n15266_, new_n15267_,
    new_n15268_, new_n15269_, new_n15270_, new_n15271_, new_n15272_,
    new_n15273_, new_n15274_, new_n15275_, new_n15276_, new_n15277_,
    new_n15278_, new_n15279_, new_n15280_, new_n15281_, new_n15282_,
    new_n15283_, new_n15284_, new_n15285_, new_n15286_, new_n15287_,
    new_n15288_, new_n15289_, new_n15290_, new_n15291_, new_n15292_,
    new_n15293_, new_n15294_, new_n15295_, new_n15296_, new_n15297_,
    new_n15298_, new_n15299_, new_n15300_, new_n15301_, new_n15302_,
    new_n15303_, new_n15304_, new_n15305_, new_n15306_, new_n15307_,
    new_n15308_, new_n15309_, new_n15310_, new_n15311_, new_n15312_,
    new_n15313_, new_n15314_, new_n15315_, new_n15316_, new_n15317_,
    new_n15318_, new_n15319_, new_n15320_, new_n15321_, new_n15322_,
    new_n15323_, new_n15324_, new_n15325_, new_n15326_, new_n15327_,
    new_n15328_, new_n15329_, new_n15330_, new_n15331_, new_n15332_,
    new_n15333_, new_n15334_, new_n15335_, new_n15336_, new_n15337_,
    new_n15338_, new_n15339_, new_n15340_, new_n15341_, new_n15342_,
    new_n15343_, new_n15344_, new_n15345_, new_n15346_, new_n15347_,
    new_n15348_, new_n15349_, new_n15350_, new_n15351_, new_n15352_,
    new_n15353_, new_n15354_, new_n15355_, new_n15356_, new_n15357_,
    new_n15358_, new_n15359_, new_n15360_, new_n15361_, new_n15362_,
    new_n15363_, new_n15364_, new_n15365_, new_n15366_, new_n15367_,
    new_n15368_, new_n15369_, new_n15370_, new_n15371_, new_n15372_,
    new_n15373_, new_n15374_, new_n15375_, new_n15376_, new_n15377_,
    new_n15378_, new_n15379_, new_n15380_, new_n15381_, new_n15382_,
    new_n15383_, new_n15384_, new_n15385_, new_n15386_, new_n15387_,
    new_n15388_, new_n15389_, new_n15390_, new_n15391_, new_n15392_,
    new_n15393_, new_n15394_, new_n15395_, new_n15396_, new_n15397_,
    new_n15398_, new_n15399_, new_n15400_, new_n15401_, new_n15402_,
    new_n15403_, new_n15404_, new_n15405_, new_n15406_, new_n15407_,
    new_n15408_, new_n15409_, new_n15410_, new_n15411_, new_n15412_,
    new_n15413_, new_n15414_, new_n15415_, new_n15416_, new_n15417_,
    new_n15418_, new_n15419_, new_n15420_, new_n15421_, new_n15422_,
    new_n15423_, new_n15424_, new_n15425_, new_n15426_, new_n15427_,
    new_n15428_, new_n15429_, new_n15430_, new_n15431_, new_n15432_,
    new_n15433_, new_n15434_, new_n15435_, new_n15436_, new_n15437_,
    new_n15438_, new_n15439_, new_n15440_, new_n15441_, new_n15442_,
    new_n15443_, new_n15444_, new_n15445_, new_n15446_, new_n15447_,
    new_n15448_, new_n15449_, new_n15450_, new_n15451_, new_n15452_,
    new_n15453_, new_n15454_, new_n15455_, new_n15456_, new_n15457_,
    new_n15458_, new_n15459_, new_n15460_, new_n15461_, new_n15462_,
    new_n15463_, new_n15464_, new_n15465_, new_n15466_, new_n15467_,
    new_n15468_, new_n15469_, new_n15470_, new_n15471_, new_n15472_,
    new_n15473_, new_n15474_, new_n15475_, new_n15476_, new_n15477_,
    new_n15478_, new_n15479_, new_n15480_, new_n15481_, new_n15482_,
    new_n15483_, new_n15484_, new_n15485_, new_n15486_, new_n15487_,
    new_n15488_, new_n15489_, new_n15490_, new_n15491_, new_n15492_,
    new_n15493_, new_n15494_, new_n15495_, new_n15496_, new_n15497_,
    new_n15498_, new_n15499_, new_n15500_, new_n15501_, new_n15502_,
    new_n15503_, new_n15504_, new_n15505_, new_n15506_, new_n15507_,
    new_n15508_, new_n15509_, new_n15510_, new_n15511_, new_n15512_,
    new_n15513_, new_n15514_, new_n15515_, new_n15516_, new_n15517_,
    new_n15518_, new_n15519_, new_n15520_, new_n15521_, new_n15522_,
    new_n15523_, new_n15524_, new_n15525_, new_n15526_, new_n15527_,
    new_n15528_, new_n15529_, new_n15530_, new_n15531_, new_n15532_,
    new_n15533_, new_n15534_, new_n15535_, new_n15536_, new_n15537_,
    new_n15538_, new_n15539_, new_n15540_, new_n15541_, new_n15542_,
    new_n15543_, new_n15544_, new_n15545_, new_n15546_, new_n15547_,
    new_n15548_, new_n15549_, new_n15550_, new_n15551_, new_n15552_,
    new_n15553_, new_n15554_, new_n15555_, new_n15556_, new_n15557_,
    new_n15558_, new_n15559_, new_n15560_, new_n15561_, new_n15562_,
    new_n15563_, new_n15564_, new_n15565_, new_n15566_, new_n15567_,
    new_n15568_, new_n15569_, new_n15570_, new_n15571_, new_n15572_,
    new_n15573_, new_n15574_, new_n15575_, new_n15576_, new_n15577_,
    new_n15578_, new_n15579_, new_n15580_, new_n15581_, new_n15582_,
    new_n15583_, new_n15584_, new_n15585_, new_n15586_, new_n15587_,
    new_n15588_, new_n15589_, new_n15590_, new_n15591_, new_n15592_,
    new_n15593_, new_n15594_, new_n15595_, new_n15596_, new_n15597_,
    new_n15598_, new_n15599_, new_n15600_, new_n15601_, new_n15602_,
    new_n15603_, new_n15604_, new_n15605_, new_n15606_, new_n15607_,
    new_n15608_, new_n15609_, new_n15610_, new_n15611_, new_n15612_,
    new_n15613_, new_n15614_, new_n15615_, new_n15616_, new_n15617_,
    new_n15618_, new_n15619_, new_n15620_, new_n15621_, new_n15622_,
    new_n15623_, new_n15624_, new_n15625_, new_n15626_, new_n15627_,
    new_n15628_, new_n15629_, new_n15630_, new_n15631_, new_n15632_,
    new_n15633_, new_n15634_, new_n15635_, new_n15636_, new_n15637_,
    new_n15638_, new_n15639_, new_n15640_, new_n15641_, new_n15642_,
    new_n15643_, new_n15644_, new_n15645_, new_n15646_, new_n15647_,
    new_n15648_, new_n15649_, new_n15650_, new_n15651_, new_n15652_,
    new_n15653_, new_n15654_, new_n15655_, new_n15656_, new_n15657_,
    new_n15658_, new_n15659_, new_n15660_, new_n15661_, new_n15662_,
    new_n15663_, new_n15664_, new_n15665_, new_n15666_, new_n15667_,
    new_n15668_, new_n15669_, new_n15670_, new_n15671_, new_n15672_,
    new_n15673_, new_n15674_, new_n15675_, new_n15676_, new_n15677_,
    new_n15678_, new_n15679_, new_n15680_, new_n15681_, new_n15682_,
    new_n15683_, new_n15684_, new_n15685_, new_n15686_, new_n15687_,
    new_n15688_, new_n15689_, new_n15690_, new_n15691_, new_n15692_,
    new_n15693_, new_n15694_, new_n15695_, new_n15696_, new_n15697_,
    new_n15698_, new_n15699_, new_n15700_, new_n15701_, new_n15702_,
    new_n15703_, new_n15704_, new_n15705_, new_n15706_, new_n15707_,
    new_n15708_, new_n15709_, new_n15710_, new_n15711_, new_n15712_,
    new_n15713_, new_n15714_, new_n15715_, new_n15716_, new_n15717_,
    new_n15718_, new_n15719_, new_n15720_, new_n15721_, new_n15722_,
    new_n15723_, new_n15724_, new_n15725_, new_n15726_, new_n15727_,
    new_n15728_, new_n15729_, new_n15730_, new_n15731_, new_n15732_,
    new_n15733_, new_n15734_, new_n15735_, new_n15736_, new_n15737_,
    new_n15738_, new_n15739_, new_n15740_, new_n15741_, new_n15742_,
    new_n15743_, new_n15744_, new_n15745_, new_n15746_, new_n15747_,
    new_n15748_, new_n15749_, new_n15750_, new_n15751_, new_n15752_,
    new_n15753_, new_n15754_, new_n15755_, new_n15756_, new_n15757_,
    new_n15758_, new_n15759_, new_n15760_, new_n15761_, new_n15762_,
    new_n15763_, new_n15764_, new_n15765_, new_n15766_, new_n15767_,
    new_n15768_, new_n15769_, new_n15770_, new_n15771_, new_n15772_,
    new_n15773_, new_n15774_, new_n15775_, new_n15776_, new_n15777_,
    new_n15778_, new_n15779_, new_n15780_, new_n15781_, new_n15782_,
    new_n15783_, new_n15784_, new_n15785_, new_n15786_, new_n15787_,
    new_n15788_, new_n15789_, new_n15790_, new_n15791_, new_n15792_,
    new_n15793_, new_n15794_, new_n15795_, new_n15796_, new_n15797_,
    new_n15798_, new_n15799_, new_n15800_, new_n15801_, new_n15802_,
    new_n15803_, new_n15804_, new_n15805_, new_n15806_, new_n15807_,
    new_n15808_, new_n15809_, new_n15810_, new_n15811_, new_n15812_,
    new_n15813_, new_n15814_, new_n15815_, new_n15816_, new_n15817_,
    new_n15818_, new_n15819_, new_n15820_, new_n15821_, new_n15822_,
    new_n15823_, new_n15824_, new_n15825_, new_n15826_, new_n15827_,
    new_n15828_, new_n15829_, new_n15830_, new_n15831_, new_n15832_,
    new_n15833_, new_n15834_, new_n15835_, new_n15836_, new_n15837_,
    new_n15838_, new_n15839_, new_n15840_, new_n15841_, new_n15842_,
    new_n15843_, new_n15844_, new_n15845_, new_n15846_, new_n15847_,
    new_n15848_, new_n15849_, new_n15850_, new_n15851_, new_n15852_,
    new_n15853_, new_n15854_, new_n15855_, new_n15856_, new_n15857_,
    new_n15858_, new_n15859_, new_n15860_, new_n15861_, new_n15862_,
    new_n15863_, new_n15865_, new_n15866_, new_n15867_, new_n15868_,
    new_n15869_, new_n15870_, new_n15871_, new_n15872_, new_n15873_,
    new_n15874_, new_n15875_, new_n15876_, new_n15877_, new_n15878_,
    new_n15879_, new_n15880_, new_n15881_, new_n15882_, new_n15883_,
    new_n15884_, new_n15885_, new_n15886_, new_n15887_, new_n15888_,
    new_n15889_, new_n15890_, new_n15891_, new_n15892_, new_n15893_,
    new_n15894_, new_n15895_, new_n15896_, new_n15897_, new_n15898_,
    new_n15899_, new_n15900_, new_n15901_, new_n15902_, new_n15903_,
    new_n15904_, new_n15905_, new_n15906_, new_n15907_, new_n15908_,
    new_n15909_, new_n15910_, new_n15911_, new_n15912_, new_n15913_,
    new_n15914_, new_n15915_, new_n15916_, new_n15917_, new_n15918_,
    new_n15919_, new_n15920_, new_n15921_, new_n15922_, new_n15923_,
    new_n15924_, new_n15925_, new_n15926_, new_n15927_, new_n15928_,
    new_n15929_, new_n15930_, new_n15931_, new_n15932_, new_n15933_,
    new_n15934_, new_n15935_, new_n15936_, new_n15937_, new_n15938_,
    new_n15939_, new_n15940_, new_n15941_, new_n15942_, new_n15943_,
    new_n15944_, new_n15945_, new_n15946_, new_n15947_, new_n15948_,
    new_n15949_, new_n15950_, new_n15951_, new_n15952_, new_n15953_,
    new_n15954_, new_n15955_, new_n15956_, new_n15957_, new_n15958_,
    new_n15959_, new_n15960_, new_n15961_, new_n15962_, new_n15963_,
    new_n15964_, new_n15965_, new_n15966_, new_n15967_, new_n15968_,
    new_n15969_, new_n15970_, new_n15971_, new_n15972_, new_n15973_,
    new_n15974_, new_n15975_, new_n15976_, new_n15977_, new_n15978_,
    new_n15979_, new_n15980_, new_n15981_, new_n15982_, new_n15983_,
    new_n15984_, new_n15985_, new_n15986_, new_n15987_, new_n15988_,
    new_n15989_, new_n15990_, new_n15991_, new_n15992_, new_n15993_,
    new_n15994_, new_n15995_, new_n15996_, new_n15997_, new_n15998_,
    new_n15999_, new_n16000_, new_n16001_, new_n16002_, new_n16003_,
    new_n16004_, new_n16005_, new_n16006_, new_n16007_, new_n16008_,
    new_n16009_, new_n16010_, new_n16011_, new_n16012_, new_n16013_,
    new_n16014_, new_n16015_, new_n16016_, new_n16017_, new_n16018_,
    new_n16019_, new_n16020_, new_n16021_, new_n16022_, new_n16023_,
    new_n16024_, new_n16025_, new_n16026_, new_n16027_, new_n16028_,
    new_n16029_, new_n16030_, new_n16031_, new_n16032_, new_n16033_,
    new_n16034_, new_n16035_, new_n16036_, new_n16037_, new_n16038_,
    new_n16039_, new_n16040_, new_n16041_, new_n16042_, new_n16043_,
    new_n16044_, new_n16045_, new_n16046_, new_n16047_, new_n16048_,
    new_n16049_, new_n16050_, new_n16051_, new_n16052_, new_n16053_,
    new_n16054_, new_n16055_, new_n16056_, new_n16057_, new_n16058_,
    new_n16059_, new_n16060_, new_n16061_, new_n16062_, new_n16063_,
    new_n16064_, new_n16065_, new_n16066_, new_n16067_, new_n16068_,
    new_n16069_, new_n16070_, new_n16071_, new_n16072_, new_n16073_,
    new_n16074_, new_n16075_, new_n16076_, new_n16077_, new_n16078_,
    new_n16079_, new_n16080_, new_n16081_, new_n16082_, new_n16083_,
    new_n16084_, new_n16085_, new_n16086_, new_n16087_, new_n16088_,
    new_n16089_, new_n16090_, new_n16091_, new_n16092_, new_n16093_,
    new_n16094_, new_n16095_, new_n16096_, new_n16097_, new_n16098_,
    new_n16099_, new_n16100_, new_n16101_, new_n16102_, new_n16103_,
    new_n16104_, new_n16105_, new_n16106_, new_n16107_, new_n16108_,
    new_n16109_, new_n16110_, new_n16111_, new_n16112_, new_n16113_,
    new_n16114_, new_n16115_, new_n16116_, new_n16117_, new_n16118_,
    new_n16119_, new_n16120_, new_n16121_, new_n16122_, new_n16123_,
    new_n16124_, new_n16125_, new_n16126_, new_n16127_, new_n16128_,
    new_n16129_, new_n16130_, new_n16131_, new_n16132_, new_n16133_,
    new_n16134_, new_n16135_, new_n16136_, new_n16137_, new_n16138_,
    new_n16139_, new_n16140_, new_n16141_, new_n16142_, new_n16143_,
    new_n16144_, new_n16145_, new_n16146_, new_n16147_, new_n16148_,
    new_n16149_, new_n16150_, new_n16151_, new_n16152_, new_n16153_,
    new_n16154_, new_n16155_, new_n16156_, new_n16157_, new_n16158_,
    new_n16159_, new_n16160_, new_n16161_, new_n16162_, new_n16163_,
    new_n16164_, new_n16165_, new_n16166_, new_n16167_, new_n16168_,
    new_n16169_, new_n16170_, new_n16171_, new_n16172_, new_n16173_,
    new_n16174_, new_n16175_, new_n16176_, new_n16177_, new_n16178_,
    new_n16179_, new_n16180_, new_n16181_, new_n16182_, new_n16183_,
    new_n16184_, new_n16185_, new_n16186_, new_n16187_, new_n16188_,
    new_n16189_, new_n16190_, new_n16191_, new_n16192_, new_n16193_,
    new_n16194_, new_n16195_, new_n16196_, new_n16197_, new_n16198_,
    new_n16199_, new_n16200_, new_n16201_, new_n16202_, new_n16203_,
    new_n16204_, new_n16205_, new_n16206_, new_n16207_, new_n16208_,
    new_n16209_, new_n16210_, new_n16211_, new_n16212_, new_n16213_,
    new_n16214_, new_n16215_, new_n16216_, new_n16217_, new_n16218_,
    new_n16219_, new_n16220_, new_n16221_, new_n16222_, new_n16223_,
    new_n16224_, new_n16225_, new_n16226_, new_n16227_, new_n16228_,
    new_n16229_, new_n16230_, new_n16231_, new_n16232_, new_n16233_,
    new_n16234_, new_n16235_, new_n16236_, new_n16237_, new_n16238_,
    new_n16239_, new_n16240_, new_n16241_, new_n16242_, new_n16243_,
    new_n16244_, new_n16245_, new_n16246_, new_n16247_, new_n16248_,
    new_n16249_, new_n16250_, new_n16251_, new_n16252_, new_n16253_,
    new_n16254_, new_n16255_, new_n16256_, new_n16257_, new_n16258_,
    new_n16259_, new_n16260_, new_n16261_, new_n16262_, new_n16263_,
    new_n16264_, new_n16265_, new_n16266_, new_n16267_, new_n16268_,
    new_n16269_, new_n16270_, new_n16271_, new_n16272_, new_n16273_,
    new_n16274_, new_n16275_, new_n16276_, new_n16277_, new_n16278_,
    new_n16279_, new_n16280_, new_n16281_, new_n16282_, new_n16283_,
    new_n16284_, new_n16285_, new_n16286_, new_n16287_, new_n16288_,
    new_n16289_, new_n16290_, new_n16291_, new_n16292_, new_n16293_,
    new_n16294_, new_n16295_, new_n16296_, new_n16297_, new_n16298_,
    new_n16299_, new_n16300_, new_n16301_, new_n16302_, new_n16303_,
    new_n16304_, new_n16305_, new_n16306_, new_n16307_, new_n16308_,
    new_n16309_, new_n16310_, new_n16311_, new_n16312_, new_n16313_,
    new_n16314_, new_n16315_, new_n16316_, new_n16317_, new_n16318_,
    new_n16319_, new_n16320_, new_n16321_, new_n16322_, new_n16323_,
    new_n16324_, new_n16325_, new_n16326_, new_n16327_, new_n16328_,
    new_n16329_, new_n16330_, new_n16331_, new_n16332_, new_n16333_,
    new_n16334_, new_n16335_, new_n16336_, new_n16337_, new_n16338_,
    new_n16339_, new_n16340_, new_n16341_, new_n16342_, new_n16343_,
    new_n16344_, new_n16345_, new_n16346_, new_n16347_, new_n16348_,
    new_n16349_, new_n16350_, new_n16351_, new_n16352_, new_n16353_,
    new_n16354_, new_n16355_, new_n16356_, new_n16357_, new_n16358_,
    new_n16359_, new_n16360_, new_n16361_, new_n16362_, new_n16363_,
    new_n16364_, new_n16365_, new_n16366_, new_n16367_, new_n16368_,
    new_n16369_, new_n16370_, new_n16371_, new_n16372_, new_n16373_,
    new_n16374_, new_n16375_, new_n16376_, new_n16377_, new_n16378_,
    new_n16379_, new_n16380_, new_n16381_, new_n16382_, new_n16383_,
    new_n16384_, new_n16385_, new_n16386_, new_n16387_, new_n16388_,
    new_n16389_, new_n16390_, new_n16391_, new_n16392_, new_n16393_,
    new_n16394_, new_n16395_, new_n16396_, new_n16397_, new_n16398_,
    new_n16399_, new_n16400_, new_n16401_, new_n16402_, new_n16403_,
    new_n16404_, new_n16405_, new_n16406_, new_n16407_, new_n16408_,
    new_n16409_, new_n16410_, new_n16411_, new_n16412_, new_n16413_,
    new_n16414_, new_n16415_, new_n16416_, new_n16417_, new_n16418_,
    new_n16419_, new_n16420_, new_n16421_, new_n16422_, new_n16423_,
    new_n16424_, new_n16425_, new_n16426_, new_n16427_, new_n16428_,
    new_n16429_, new_n16430_, new_n16431_, new_n16432_, new_n16433_,
    new_n16434_, new_n16435_, new_n16436_, new_n16437_, new_n16438_,
    new_n16439_, new_n16440_, new_n16441_, new_n16442_, new_n16443_,
    new_n16444_, new_n16445_, new_n16446_, new_n16447_, new_n16448_,
    new_n16449_, new_n16450_, new_n16451_, new_n16452_, new_n16453_,
    new_n16454_, new_n16455_, new_n16456_, new_n16457_, new_n16458_,
    new_n16459_, new_n16460_, new_n16461_, new_n16462_, new_n16463_,
    new_n16464_, new_n16465_, new_n16466_, new_n16467_, new_n16468_,
    new_n16469_, new_n16470_, new_n16471_, new_n16472_, new_n16473_,
    new_n16474_, new_n16475_, new_n16476_, new_n16477_, new_n16478_,
    new_n16479_, new_n16480_, new_n16481_, new_n16482_, new_n16483_,
    new_n16484_, new_n16485_, new_n16486_, new_n16487_, new_n16488_,
    new_n16489_, new_n16490_, new_n16491_, new_n16492_, new_n16493_,
    new_n16494_, new_n16495_, new_n16496_, new_n16497_, new_n16498_,
    new_n16499_, new_n16500_, new_n16501_, new_n16502_, new_n16503_,
    new_n16504_, new_n16505_, new_n16506_, new_n16507_, new_n16508_,
    new_n16509_, new_n16510_, new_n16511_, new_n16512_, new_n16513_,
    new_n16514_, new_n16515_, new_n16516_, new_n16517_, new_n16518_,
    new_n16519_, new_n16520_, new_n16521_, new_n16522_, new_n16524_,
    new_n16525_, new_n16526_, new_n16527_, new_n16528_, new_n16529_,
    new_n16530_, new_n16531_, new_n16532_, new_n16533_, new_n16534_,
    new_n16535_, new_n16536_, new_n16537_, new_n16538_, new_n16539_,
    new_n16540_, new_n16541_, new_n16542_, new_n16543_, new_n16544_,
    new_n16545_, new_n16546_, new_n16547_, new_n16548_, new_n16549_,
    new_n16550_, new_n16551_, new_n16552_, new_n16553_, new_n16554_,
    new_n16555_, new_n16556_, new_n16557_, new_n16558_, new_n16559_,
    new_n16560_, new_n16561_, new_n16562_, new_n16563_, new_n16564_,
    new_n16565_, new_n16566_, new_n16567_, new_n16568_, new_n16569_,
    new_n16570_, new_n16571_, new_n16572_, new_n16573_, new_n16574_,
    new_n16575_, new_n16576_, new_n16577_, new_n16578_, new_n16579_,
    new_n16580_, new_n16581_, new_n16582_, new_n16583_, new_n16584_,
    new_n16585_, new_n16586_, new_n16587_, new_n16588_, new_n16589_,
    new_n16590_, new_n16591_, new_n16592_, new_n16593_, new_n16594_,
    new_n16595_, new_n16596_, new_n16597_, new_n16598_, new_n16599_,
    new_n16600_, new_n16601_, new_n16602_, new_n16603_, new_n16604_,
    new_n16605_, new_n16606_, new_n16607_, new_n16608_, new_n16609_,
    new_n16610_, new_n16611_, new_n16612_, new_n16613_, new_n16614_,
    new_n16615_, new_n16616_, new_n16617_, new_n16618_, new_n16619_,
    new_n16620_, new_n16621_, new_n16622_, new_n16623_, new_n16624_,
    new_n16625_, new_n16626_, new_n16627_, new_n16628_, new_n16629_,
    new_n16630_, new_n16631_, new_n16632_, new_n16633_, new_n16634_,
    new_n16635_, new_n16636_, new_n16637_, new_n16638_, new_n16639_,
    new_n16640_, new_n16641_, new_n16642_, new_n16643_, new_n16644_,
    new_n16645_, new_n16646_, new_n16647_, new_n16648_, new_n16649_,
    new_n16650_, new_n16651_, new_n16652_, new_n16653_, new_n16654_,
    new_n16655_, new_n16656_, new_n16657_, new_n16658_, new_n16659_,
    new_n16660_, new_n16661_, new_n16662_, new_n16663_, new_n16664_,
    new_n16665_, new_n16666_, new_n16667_, new_n16668_, new_n16669_,
    new_n16670_, new_n16671_, new_n16672_, new_n16673_, new_n16674_,
    new_n16675_, new_n16676_, new_n16677_, new_n16678_, new_n16679_,
    new_n16680_, new_n16681_, new_n16682_, new_n16683_, new_n16684_,
    new_n16685_, new_n16686_, new_n16687_, new_n16688_, new_n16689_,
    new_n16690_, new_n16691_, new_n16692_, new_n16693_, new_n16694_,
    new_n16695_, new_n16696_, new_n16697_, new_n16698_, new_n16699_,
    new_n16700_, new_n16701_, new_n16702_, new_n16703_, new_n16704_,
    new_n16705_, new_n16706_, new_n16707_, new_n16708_, new_n16709_,
    new_n16710_, new_n16711_, new_n16712_, new_n16713_, new_n16714_,
    new_n16715_, new_n16716_, new_n16717_, new_n16718_, new_n16719_,
    new_n16720_, new_n16721_, new_n16722_, new_n16723_, new_n16724_,
    new_n16725_, new_n16726_, new_n16727_, new_n16728_, new_n16729_,
    new_n16730_, new_n16731_, new_n16732_, new_n16733_, new_n16734_,
    new_n16735_, new_n16736_, new_n16737_, new_n16738_, new_n16739_,
    new_n16740_, new_n16741_, new_n16742_, new_n16743_, new_n16744_,
    new_n16745_, new_n16746_, new_n16747_, new_n16748_, new_n16749_,
    new_n16750_, new_n16751_, new_n16752_, new_n16753_, new_n16754_,
    new_n16755_, new_n16756_, new_n16757_, new_n16758_, new_n16759_,
    new_n16760_, new_n16761_, new_n16762_, new_n16763_, new_n16764_,
    new_n16765_, new_n16766_, new_n16767_, new_n16768_, new_n16769_,
    new_n16770_, new_n16771_, new_n16772_, new_n16773_, new_n16774_,
    new_n16775_, new_n16776_, new_n16777_, new_n16778_, new_n16779_,
    new_n16780_, new_n16781_, new_n16782_, new_n16783_, new_n16784_,
    new_n16785_, new_n16786_, new_n16787_, new_n16788_, new_n16789_,
    new_n16790_, new_n16791_, new_n16792_, new_n16793_, new_n16794_,
    new_n16795_, new_n16796_, new_n16797_, new_n16798_, new_n16799_,
    new_n16800_, new_n16801_, new_n16802_, new_n16803_, new_n16804_,
    new_n16805_, new_n16806_, new_n16807_, new_n16808_, new_n16809_,
    new_n16810_, new_n16811_, new_n16812_, new_n16813_, new_n16814_,
    new_n16815_, new_n16816_, new_n16817_, new_n16818_, new_n16819_,
    new_n16820_, new_n16821_, new_n16822_, new_n16823_, new_n16824_,
    new_n16825_, new_n16826_, new_n16827_, new_n16828_, new_n16829_,
    new_n16830_, new_n16831_, new_n16832_, new_n16833_, new_n16834_,
    new_n16835_, new_n16836_, new_n16837_, new_n16838_, new_n16839_,
    new_n16840_, new_n16841_, new_n16842_, new_n16843_, new_n16844_,
    new_n16845_, new_n16846_, new_n16847_, new_n16848_, new_n16849_,
    new_n16850_, new_n16851_, new_n16852_, new_n16853_, new_n16854_,
    new_n16855_, new_n16856_, new_n16857_, new_n16858_, new_n16859_,
    new_n16860_, new_n16861_, new_n16862_, new_n16863_, new_n16864_,
    new_n16865_, new_n16866_, new_n16867_, new_n16868_, new_n16869_,
    new_n16870_, new_n16871_, new_n16872_, new_n16873_, new_n16874_,
    new_n16875_, new_n16876_, new_n16877_, new_n16878_, new_n16879_,
    new_n16880_, new_n16881_, new_n16882_, new_n16883_, new_n16884_,
    new_n16885_, new_n16886_, new_n16887_, new_n16888_, new_n16889_,
    new_n16890_, new_n16891_, new_n16892_, new_n16893_, new_n16894_,
    new_n16895_, new_n16896_, new_n16897_, new_n16898_, new_n16899_,
    new_n16900_, new_n16901_, new_n16902_, new_n16903_, new_n16904_,
    new_n16905_, new_n16906_, new_n16907_, new_n16908_, new_n16909_,
    new_n16910_, new_n16911_, new_n16912_, new_n16913_, new_n16914_,
    new_n16915_, new_n16916_, new_n16917_, new_n16918_, new_n16919_,
    new_n16920_, new_n16921_, new_n16922_, new_n16923_, new_n16924_,
    new_n16925_, new_n16926_, new_n16927_, new_n16928_, new_n16929_,
    new_n16930_, new_n16931_, new_n16932_, new_n16933_, new_n16934_,
    new_n16935_, new_n16936_, new_n16937_, new_n16938_, new_n16939_,
    new_n16940_, new_n16941_, new_n16942_, new_n16943_, new_n16944_,
    new_n16945_, new_n16946_, new_n16947_, new_n16948_, new_n16949_,
    new_n16950_, new_n16951_, new_n16952_, new_n16953_, new_n16954_,
    new_n16955_, new_n16956_, new_n16957_, new_n16958_, new_n16959_,
    new_n16960_, new_n16961_, new_n16962_, new_n16963_, new_n16964_,
    new_n16965_, new_n16966_, new_n16967_, new_n16968_, new_n16969_,
    new_n16970_, new_n16971_, new_n16972_, new_n16973_, new_n16974_,
    new_n16975_, new_n16976_, new_n16977_, new_n16978_, new_n16979_,
    new_n16980_, new_n16981_, new_n16982_, new_n16983_, new_n16984_,
    new_n16985_, new_n16986_, new_n16987_, new_n16988_, new_n16989_,
    new_n16990_, new_n16991_, new_n16992_, new_n16993_, new_n16994_,
    new_n16995_, new_n16996_, new_n16997_, new_n16998_, new_n16999_,
    new_n17000_, new_n17001_, new_n17002_, new_n17003_, new_n17004_,
    new_n17005_, new_n17006_, new_n17007_, new_n17008_, new_n17009_,
    new_n17010_, new_n17011_, new_n17012_, new_n17013_, new_n17014_,
    new_n17015_, new_n17016_, new_n17017_, new_n17018_, new_n17019_,
    new_n17020_, new_n17021_, new_n17022_, new_n17023_, new_n17024_,
    new_n17025_, new_n17026_, new_n17027_, new_n17028_, new_n17029_,
    new_n17030_, new_n17031_, new_n17032_, new_n17033_, new_n17034_,
    new_n17035_, new_n17036_, new_n17037_, new_n17038_, new_n17039_,
    new_n17040_, new_n17041_, new_n17042_, new_n17043_, new_n17044_,
    new_n17045_, new_n17046_, new_n17047_, new_n17048_, new_n17049_,
    new_n17050_, new_n17051_, new_n17052_, new_n17053_, new_n17054_,
    new_n17055_, new_n17056_, new_n17057_, new_n17058_, new_n17059_,
    new_n17060_, new_n17061_, new_n17062_, new_n17063_, new_n17064_,
    new_n17065_, new_n17066_, new_n17067_, new_n17068_, new_n17069_,
    new_n17070_, new_n17071_, new_n17072_, new_n17073_, new_n17074_,
    new_n17075_, new_n17076_, new_n17077_, new_n17078_, new_n17079_,
    new_n17080_, new_n17081_, new_n17082_, new_n17083_, new_n17084_,
    new_n17085_, new_n17086_, new_n17087_, new_n17088_, new_n17089_,
    new_n17090_, new_n17091_, new_n17092_, new_n17093_, new_n17094_,
    new_n17095_, new_n17096_, new_n17097_, new_n17098_, new_n17099_,
    new_n17100_, new_n17101_, new_n17102_, new_n17103_, new_n17104_,
    new_n17105_, new_n17106_, new_n17107_, new_n17108_, new_n17109_,
    new_n17110_, new_n17111_, new_n17112_, new_n17113_, new_n17114_,
    new_n17115_, new_n17116_, new_n17117_, new_n17118_, new_n17119_,
    new_n17120_, new_n17121_, new_n17122_, new_n17123_, new_n17124_,
    new_n17125_, new_n17126_, new_n17127_, new_n17128_, new_n17129_,
    new_n17130_, new_n17131_, new_n17132_, new_n17133_, new_n17134_,
    new_n17135_, new_n17136_, new_n17137_, new_n17138_, new_n17139_,
    new_n17140_, new_n17141_, new_n17142_, new_n17143_, new_n17144_,
    new_n17145_, new_n17146_, new_n17147_, new_n17148_, new_n17149_,
    new_n17150_, new_n17151_, new_n17152_, new_n17153_, new_n17154_,
    new_n17155_, new_n17156_, new_n17157_, new_n17158_, new_n17159_,
    new_n17160_, new_n17161_, new_n17162_, new_n17163_, new_n17164_,
    new_n17165_, new_n17166_, new_n17167_, new_n17168_, new_n17169_,
    new_n17170_, new_n17171_, new_n17172_, new_n17173_, new_n17174_,
    new_n17175_, new_n17176_, new_n17177_, new_n17178_, new_n17179_,
    new_n17180_, new_n17181_, new_n17182_, new_n17183_, new_n17184_,
    new_n17185_, new_n17186_, new_n17187_, new_n17188_, new_n17189_,
    new_n17190_, new_n17191_, new_n17192_, new_n17193_, new_n17194_,
    new_n17196_, new_n17197_, new_n17198_, new_n17199_, new_n17200_,
    new_n17201_, new_n17202_, new_n17203_, new_n17204_, new_n17205_,
    new_n17206_, new_n17207_, new_n17208_, new_n17209_, new_n17210_,
    new_n17211_, new_n17212_, new_n17213_, new_n17214_, new_n17215_,
    new_n17216_, new_n17217_, new_n17218_, new_n17219_, new_n17220_,
    new_n17221_, new_n17222_, new_n17223_, new_n17224_, new_n17225_,
    new_n17226_, new_n17227_, new_n17228_, new_n17229_, new_n17230_,
    new_n17231_, new_n17232_, new_n17233_, new_n17234_, new_n17235_,
    new_n17236_, new_n17237_, new_n17238_, new_n17239_, new_n17240_,
    new_n17241_, new_n17242_, new_n17243_, new_n17244_, new_n17245_,
    new_n17246_, new_n17247_, new_n17248_, new_n17249_, new_n17250_,
    new_n17251_, new_n17252_, new_n17253_, new_n17254_, new_n17255_,
    new_n17256_, new_n17257_, new_n17258_, new_n17259_, new_n17260_,
    new_n17261_, new_n17262_, new_n17263_, new_n17264_, new_n17265_,
    new_n17266_, new_n17267_, new_n17268_, new_n17269_, new_n17270_,
    new_n17271_, new_n17272_, new_n17273_, new_n17274_, new_n17275_,
    new_n17276_, new_n17277_, new_n17278_, new_n17279_, new_n17280_,
    new_n17281_, new_n17282_, new_n17283_, new_n17284_, new_n17285_,
    new_n17286_, new_n17287_, new_n17288_, new_n17289_, new_n17290_,
    new_n17291_, new_n17292_, new_n17293_, new_n17294_, new_n17295_,
    new_n17296_, new_n17297_, new_n17298_, new_n17299_, new_n17300_,
    new_n17301_, new_n17302_, new_n17303_, new_n17304_, new_n17305_,
    new_n17306_, new_n17307_, new_n17308_, new_n17309_, new_n17310_,
    new_n17311_, new_n17312_, new_n17313_, new_n17314_, new_n17315_,
    new_n17316_, new_n17317_, new_n17318_, new_n17319_, new_n17320_,
    new_n17321_, new_n17322_, new_n17323_, new_n17324_, new_n17325_,
    new_n17326_, new_n17327_, new_n17328_, new_n17329_, new_n17330_,
    new_n17331_, new_n17332_, new_n17333_, new_n17334_, new_n17335_,
    new_n17336_, new_n17337_, new_n17338_, new_n17339_, new_n17340_,
    new_n17341_, new_n17342_, new_n17343_, new_n17344_, new_n17345_,
    new_n17346_, new_n17347_, new_n17348_, new_n17349_, new_n17350_,
    new_n17351_, new_n17352_, new_n17353_, new_n17354_, new_n17355_,
    new_n17356_, new_n17357_, new_n17358_, new_n17359_, new_n17360_,
    new_n17361_, new_n17362_, new_n17363_, new_n17364_, new_n17365_,
    new_n17366_, new_n17367_, new_n17368_, new_n17369_, new_n17370_,
    new_n17371_, new_n17372_, new_n17373_, new_n17374_, new_n17375_,
    new_n17376_, new_n17377_, new_n17378_, new_n17379_, new_n17380_,
    new_n17381_, new_n17382_, new_n17383_, new_n17384_, new_n17385_,
    new_n17386_, new_n17387_, new_n17388_, new_n17389_, new_n17390_,
    new_n17391_, new_n17392_, new_n17393_, new_n17394_, new_n17395_,
    new_n17396_, new_n17397_, new_n17398_, new_n17399_, new_n17400_,
    new_n17401_, new_n17402_, new_n17403_, new_n17404_, new_n17405_,
    new_n17406_, new_n17407_, new_n17408_, new_n17409_, new_n17410_,
    new_n17411_, new_n17412_, new_n17413_, new_n17414_, new_n17415_,
    new_n17416_, new_n17417_, new_n17418_, new_n17419_, new_n17420_,
    new_n17421_, new_n17422_, new_n17423_, new_n17424_, new_n17425_,
    new_n17426_, new_n17427_, new_n17428_, new_n17429_, new_n17430_,
    new_n17431_, new_n17432_, new_n17433_, new_n17434_, new_n17435_,
    new_n17436_, new_n17437_, new_n17438_, new_n17439_, new_n17440_,
    new_n17441_, new_n17442_, new_n17443_, new_n17444_, new_n17445_,
    new_n17446_, new_n17447_, new_n17448_, new_n17449_, new_n17450_,
    new_n17451_, new_n17452_, new_n17453_, new_n17454_, new_n17455_,
    new_n17456_, new_n17457_, new_n17458_, new_n17459_, new_n17460_,
    new_n17461_, new_n17462_, new_n17463_, new_n17464_, new_n17465_,
    new_n17466_, new_n17467_, new_n17468_, new_n17469_, new_n17470_,
    new_n17471_, new_n17472_, new_n17473_, new_n17474_, new_n17475_,
    new_n17476_, new_n17477_, new_n17478_, new_n17479_, new_n17480_,
    new_n17481_, new_n17482_, new_n17483_, new_n17484_, new_n17485_,
    new_n17486_, new_n17487_, new_n17488_, new_n17489_, new_n17490_,
    new_n17491_, new_n17492_, new_n17493_, new_n17494_, new_n17495_,
    new_n17496_, new_n17497_, new_n17498_, new_n17499_, new_n17500_,
    new_n17501_, new_n17502_, new_n17503_, new_n17504_, new_n17505_,
    new_n17506_, new_n17507_, new_n17508_, new_n17509_, new_n17510_,
    new_n17511_, new_n17512_, new_n17513_, new_n17514_, new_n17515_,
    new_n17516_, new_n17517_, new_n17518_, new_n17519_, new_n17520_,
    new_n17521_, new_n17522_, new_n17523_, new_n17524_, new_n17525_,
    new_n17526_, new_n17527_, new_n17528_, new_n17529_, new_n17530_,
    new_n17531_, new_n17532_, new_n17533_, new_n17534_, new_n17535_,
    new_n17536_, new_n17537_, new_n17538_, new_n17539_, new_n17540_,
    new_n17541_, new_n17542_, new_n17543_, new_n17544_, new_n17545_,
    new_n17546_, new_n17547_, new_n17548_, new_n17549_, new_n17550_,
    new_n17551_, new_n17552_, new_n17553_, new_n17554_, new_n17555_,
    new_n17556_, new_n17557_, new_n17558_, new_n17559_, new_n17560_,
    new_n17561_, new_n17562_, new_n17563_, new_n17564_, new_n17565_,
    new_n17566_, new_n17567_, new_n17568_, new_n17569_, new_n17570_,
    new_n17571_, new_n17572_, new_n17573_, new_n17574_, new_n17575_,
    new_n17576_, new_n17577_, new_n17578_, new_n17579_, new_n17580_,
    new_n17581_, new_n17582_, new_n17583_, new_n17584_, new_n17585_,
    new_n17586_, new_n17587_, new_n17588_, new_n17589_, new_n17590_,
    new_n17591_, new_n17592_, new_n17593_, new_n17594_, new_n17595_,
    new_n17596_, new_n17597_, new_n17598_, new_n17599_, new_n17600_,
    new_n17601_, new_n17602_, new_n17603_, new_n17604_, new_n17605_,
    new_n17606_, new_n17607_, new_n17608_, new_n17609_, new_n17610_,
    new_n17611_, new_n17612_, new_n17613_, new_n17614_, new_n17615_,
    new_n17616_, new_n17617_, new_n17618_, new_n17619_, new_n17620_,
    new_n17621_, new_n17622_, new_n17623_, new_n17624_, new_n17625_,
    new_n17626_, new_n17627_, new_n17628_, new_n17629_, new_n17630_,
    new_n17631_, new_n17632_, new_n17633_, new_n17634_, new_n17635_,
    new_n17636_, new_n17637_, new_n17638_, new_n17639_, new_n17640_,
    new_n17641_, new_n17642_, new_n17643_, new_n17644_, new_n17645_,
    new_n17646_, new_n17647_, new_n17648_, new_n17649_, new_n17650_,
    new_n17651_, new_n17652_, new_n17653_, new_n17654_, new_n17655_,
    new_n17656_, new_n17657_, new_n17658_, new_n17659_, new_n17660_,
    new_n17661_, new_n17662_, new_n17663_, new_n17664_, new_n17665_,
    new_n17666_, new_n17667_, new_n17668_, new_n17669_, new_n17670_,
    new_n17671_, new_n17672_, new_n17673_, new_n17674_, new_n17675_,
    new_n17676_, new_n17677_, new_n17678_, new_n17679_, new_n17680_,
    new_n17681_, new_n17682_, new_n17683_, new_n17684_, new_n17685_,
    new_n17686_, new_n17687_, new_n17688_, new_n17689_, new_n17690_,
    new_n17691_, new_n17692_, new_n17693_, new_n17694_, new_n17695_,
    new_n17696_, new_n17697_, new_n17698_, new_n17699_, new_n17700_,
    new_n17701_, new_n17702_, new_n17703_, new_n17704_, new_n17705_,
    new_n17706_, new_n17707_, new_n17708_, new_n17709_, new_n17710_,
    new_n17711_, new_n17712_, new_n17713_, new_n17714_, new_n17715_,
    new_n17716_, new_n17717_, new_n17718_, new_n17719_, new_n17720_,
    new_n17721_, new_n17722_, new_n17723_, new_n17724_, new_n17725_,
    new_n17726_, new_n17727_, new_n17728_, new_n17729_, new_n17730_,
    new_n17731_, new_n17732_, new_n17733_, new_n17734_, new_n17735_,
    new_n17736_, new_n17737_, new_n17738_, new_n17739_, new_n17740_,
    new_n17741_, new_n17742_, new_n17743_, new_n17744_, new_n17745_,
    new_n17746_, new_n17747_, new_n17748_, new_n17749_, new_n17750_,
    new_n17751_, new_n17752_, new_n17753_, new_n17754_, new_n17755_,
    new_n17756_, new_n17757_, new_n17758_, new_n17759_, new_n17760_,
    new_n17761_, new_n17762_, new_n17763_, new_n17764_, new_n17765_,
    new_n17766_, new_n17767_, new_n17768_, new_n17769_, new_n17770_,
    new_n17771_, new_n17772_, new_n17773_, new_n17774_, new_n17775_,
    new_n17776_, new_n17777_, new_n17778_, new_n17779_, new_n17780_,
    new_n17781_, new_n17782_, new_n17783_, new_n17784_, new_n17785_,
    new_n17786_, new_n17787_, new_n17788_, new_n17789_, new_n17790_,
    new_n17791_, new_n17792_, new_n17793_, new_n17794_, new_n17795_,
    new_n17796_, new_n17797_, new_n17798_, new_n17799_, new_n17800_,
    new_n17801_, new_n17802_, new_n17803_, new_n17804_, new_n17805_,
    new_n17806_, new_n17807_, new_n17808_, new_n17809_, new_n17810_,
    new_n17811_, new_n17812_, new_n17813_, new_n17814_, new_n17815_,
    new_n17816_, new_n17817_, new_n17818_, new_n17819_, new_n17820_,
    new_n17821_, new_n17822_, new_n17823_, new_n17824_, new_n17825_,
    new_n17826_, new_n17827_, new_n17828_, new_n17829_, new_n17830_,
    new_n17831_, new_n17832_, new_n17833_, new_n17834_, new_n17835_,
    new_n17836_, new_n17837_, new_n17838_, new_n17839_, new_n17840_,
    new_n17841_, new_n17842_, new_n17843_, new_n17844_, new_n17845_,
    new_n17846_, new_n17847_, new_n17848_, new_n17849_, new_n17850_,
    new_n17851_, new_n17852_, new_n17853_, new_n17854_, new_n17855_,
    new_n17856_, new_n17857_, new_n17858_, new_n17859_, new_n17860_,
    new_n17861_, new_n17862_, new_n17863_, new_n17864_, new_n17865_,
    new_n17866_, new_n17867_, new_n17868_, new_n17869_, new_n17870_,
    new_n17871_, new_n17872_, new_n17873_, new_n17874_, new_n17875_,
    new_n17876_, new_n17877_, new_n17878_, new_n17879_, new_n17880_,
    new_n17881_, new_n17882_, new_n17883_, new_n17884_, new_n17885_,
    new_n17886_, new_n17888_, new_n17889_, new_n17890_, new_n17891_,
    new_n17892_, new_n17893_, new_n17894_, new_n17895_, new_n17896_,
    new_n17897_, new_n17898_, new_n17899_, new_n17900_, new_n17901_,
    new_n17902_, new_n17903_, new_n17904_, new_n17905_, new_n17906_,
    new_n17907_, new_n17908_, new_n17909_, new_n17910_, new_n17911_,
    new_n17912_, new_n17913_, new_n17914_, new_n17915_, new_n17916_,
    new_n17917_, new_n17918_, new_n17919_, new_n17920_, new_n17921_,
    new_n17922_, new_n17923_, new_n17924_, new_n17925_, new_n17926_,
    new_n17927_, new_n17928_, new_n17929_, new_n17930_, new_n17931_,
    new_n17932_, new_n17933_, new_n17934_, new_n17935_, new_n17936_,
    new_n17937_, new_n17938_, new_n17939_, new_n17940_, new_n17941_,
    new_n17942_, new_n17943_, new_n17944_, new_n17945_, new_n17946_,
    new_n17947_, new_n17948_, new_n17949_, new_n17950_, new_n17951_,
    new_n17952_, new_n17953_, new_n17954_, new_n17955_, new_n17956_,
    new_n17957_, new_n17958_, new_n17959_, new_n17960_, new_n17961_,
    new_n17962_, new_n17963_, new_n17964_, new_n17965_, new_n17966_,
    new_n17967_, new_n17968_, new_n17969_, new_n17970_, new_n17971_,
    new_n17972_, new_n17973_, new_n17974_, new_n17975_, new_n17976_,
    new_n17977_, new_n17978_, new_n17979_, new_n17980_, new_n17981_,
    new_n17982_, new_n17983_, new_n17984_, new_n17985_, new_n17986_,
    new_n17987_, new_n17988_, new_n17989_, new_n17990_, new_n17991_,
    new_n17992_, new_n17993_, new_n17994_, new_n17995_, new_n17996_,
    new_n17997_, new_n17998_, new_n17999_, new_n18000_, new_n18001_,
    new_n18002_, new_n18003_, new_n18004_, new_n18005_, new_n18006_,
    new_n18007_, new_n18008_, new_n18009_, new_n18010_, new_n18011_,
    new_n18012_, new_n18013_, new_n18014_, new_n18015_, new_n18016_,
    new_n18017_, new_n18018_, new_n18019_, new_n18020_, new_n18021_,
    new_n18022_, new_n18023_, new_n18024_, new_n18025_, new_n18026_,
    new_n18027_, new_n18028_, new_n18029_, new_n18030_, new_n18031_,
    new_n18032_, new_n18033_, new_n18034_, new_n18035_, new_n18036_,
    new_n18037_, new_n18038_, new_n18039_, new_n18040_, new_n18041_,
    new_n18042_, new_n18043_, new_n18044_, new_n18045_, new_n18046_,
    new_n18047_, new_n18048_, new_n18049_, new_n18050_, new_n18051_,
    new_n18052_, new_n18053_, new_n18054_, new_n18055_, new_n18056_,
    new_n18057_, new_n18058_, new_n18059_, new_n18060_, new_n18061_,
    new_n18062_, new_n18063_, new_n18064_, new_n18065_, new_n18066_,
    new_n18067_, new_n18068_, new_n18069_, new_n18070_, new_n18071_,
    new_n18072_, new_n18073_, new_n18074_, new_n18075_, new_n18076_,
    new_n18077_, new_n18078_, new_n18079_, new_n18080_, new_n18081_,
    new_n18082_, new_n18083_, new_n18084_, new_n18085_, new_n18086_,
    new_n18087_, new_n18088_, new_n18089_, new_n18090_, new_n18091_,
    new_n18092_, new_n18093_, new_n18094_, new_n18095_, new_n18096_,
    new_n18097_, new_n18098_, new_n18099_, new_n18100_, new_n18101_,
    new_n18102_, new_n18103_, new_n18104_, new_n18105_, new_n18106_,
    new_n18107_, new_n18108_, new_n18109_, new_n18110_, new_n18111_,
    new_n18112_, new_n18113_, new_n18114_, new_n18115_, new_n18116_,
    new_n18117_, new_n18118_, new_n18119_, new_n18120_, new_n18121_,
    new_n18122_, new_n18123_, new_n18124_, new_n18125_, new_n18126_,
    new_n18127_, new_n18128_, new_n18129_, new_n18130_, new_n18131_,
    new_n18132_, new_n18133_, new_n18134_, new_n18135_, new_n18136_,
    new_n18137_, new_n18138_, new_n18139_, new_n18140_, new_n18141_,
    new_n18142_, new_n18143_, new_n18144_, new_n18145_, new_n18146_,
    new_n18147_, new_n18148_, new_n18149_, new_n18150_, new_n18151_,
    new_n18152_, new_n18153_, new_n18154_, new_n18155_, new_n18156_,
    new_n18157_, new_n18158_, new_n18159_, new_n18160_, new_n18161_,
    new_n18162_, new_n18163_, new_n18164_, new_n18165_, new_n18166_,
    new_n18167_, new_n18168_, new_n18169_, new_n18170_, new_n18171_,
    new_n18172_, new_n18173_, new_n18174_, new_n18175_, new_n18176_,
    new_n18177_, new_n18178_, new_n18179_, new_n18180_, new_n18181_,
    new_n18182_, new_n18183_, new_n18184_, new_n18185_, new_n18186_,
    new_n18187_, new_n18188_, new_n18189_, new_n18190_, new_n18191_,
    new_n18192_, new_n18193_, new_n18194_, new_n18195_, new_n18196_,
    new_n18197_, new_n18198_, new_n18199_, new_n18200_, new_n18201_,
    new_n18202_, new_n18203_, new_n18204_, new_n18205_, new_n18206_,
    new_n18207_, new_n18208_, new_n18209_, new_n18210_, new_n18211_,
    new_n18212_, new_n18213_, new_n18214_, new_n18215_, new_n18216_,
    new_n18217_, new_n18218_, new_n18219_, new_n18220_, new_n18221_,
    new_n18222_, new_n18223_, new_n18224_, new_n18225_, new_n18226_,
    new_n18227_, new_n18228_, new_n18229_, new_n18230_, new_n18231_,
    new_n18232_, new_n18233_, new_n18234_, new_n18235_, new_n18236_,
    new_n18237_, new_n18238_, new_n18239_, new_n18240_, new_n18241_,
    new_n18242_, new_n18243_, new_n18244_, new_n18245_, new_n18246_,
    new_n18247_, new_n18248_, new_n18249_, new_n18250_, new_n18251_,
    new_n18252_, new_n18253_, new_n18254_, new_n18255_, new_n18256_,
    new_n18257_, new_n18258_, new_n18259_, new_n18260_, new_n18261_,
    new_n18262_, new_n18263_, new_n18264_, new_n18265_, new_n18266_,
    new_n18267_, new_n18268_, new_n18269_, new_n18270_, new_n18271_,
    new_n18272_, new_n18273_, new_n18274_, new_n18275_, new_n18276_,
    new_n18277_, new_n18278_, new_n18279_, new_n18280_, new_n18281_,
    new_n18282_, new_n18283_, new_n18284_, new_n18285_, new_n18286_,
    new_n18287_, new_n18288_, new_n18289_, new_n18290_, new_n18291_,
    new_n18292_, new_n18293_, new_n18294_, new_n18295_, new_n18296_,
    new_n18297_, new_n18298_, new_n18299_, new_n18300_, new_n18301_,
    new_n18302_, new_n18303_, new_n18304_, new_n18305_, new_n18306_,
    new_n18307_, new_n18308_, new_n18309_, new_n18310_, new_n18311_,
    new_n18312_, new_n18313_, new_n18314_, new_n18315_, new_n18316_,
    new_n18317_, new_n18318_, new_n18319_, new_n18320_, new_n18321_,
    new_n18322_, new_n18323_, new_n18324_, new_n18325_, new_n18326_,
    new_n18327_, new_n18328_, new_n18329_, new_n18330_, new_n18331_,
    new_n18332_, new_n18333_, new_n18334_, new_n18335_, new_n18336_,
    new_n18337_, new_n18338_, new_n18339_, new_n18340_, new_n18341_,
    new_n18342_, new_n18343_, new_n18344_, new_n18345_, new_n18346_,
    new_n18347_, new_n18348_, new_n18349_, new_n18350_, new_n18351_,
    new_n18352_, new_n18353_, new_n18354_, new_n18355_, new_n18356_,
    new_n18357_, new_n18358_, new_n18359_, new_n18360_, new_n18361_,
    new_n18362_, new_n18363_, new_n18364_, new_n18365_, new_n18366_,
    new_n18367_, new_n18368_, new_n18369_, new_n18370_, new_n18371_,
    new_n18372_, new_n18373_, new_n18374_, new_n18375_, new_n18376_,
    new_n18377_, new_n18378_, new_n18379_, new_n18380_, new_n18381_,
    new_n18382_, new_n18383_, new_n18384_, new_n18385_, new_n18386_,
    new_n18387_, new_n18388_, new_n18389_, new_n18390_, new_n18391_,
    new_n18392_, new_n18393_, new_n18394_, new_n18395_, new_n18396_,
    new_n18397_, new_n18398_, new_n18399_, new_n18400_, new_n18401_,
    new_n18402_, new_n18403_, new_n18404_, new_n18405_, new_n18406_,
    new_n18407_, new_n18408_, new_n18409_, new_n18410_, new_n18411_,
    new_n18412_, new_n18413_, new_n18414_, new_n18415_, new_n18416_,
    new_n18417_, new_n18418_, new_n18419_, new_n18420_, new_n18421_,
    new_n18422_, new_n18423_, new_n18424_, new_n18425_, new_n18426_,
    new_n18427_, new_n18428_, new_n18429_, new_n18430_, new_n18431_,
    new_n18432_, new_n18433_, new_n18434_, new_n18435_, new_n18436_,
    new_n18437_, new_n18438_, new_n18439_, new_n18440_, new_n18441_,
    new_n18442_, new_n18443_, new_n18444_, new_n18445_, new_n18446_,
    new_n18447_, new_n18448_, new_n18449_, new_n18450_, new_n18451_,
    new_n18452_, new_n18453_, new_n18454_, new_n18455_, new_n18456_,
    new_n18457_, new_n18458_, new_n18459_, new_n18460_, new_n18461_,
    new_n18462_, new_n18463_, new_n18464_, new_n18465_, new_n18466_,
    new_n18467_, new_n18468_, new_n18469_, new_n18470_, new_n18471_,
    new_n18472_, new_n18473_, new_n18474_, new_n18475_, new_n18476_,
    new_n18477_, new_n18478_, new_n18479_, new_n18480_, new_n18481_,
    new_n18482_, new_n18483_, new_n18484_, new_n18485_, new_n18486_,
    new_n18487_, new_n18488_, new_n18489_, new_n18490_, new_n18491_,
    new_n18492_, new_n18493_, new_n18494_, new_n18495_, new_n18496_,
    new_n18497_, new_n18498_, new_n18499_, new_n18500_, new_n18501_,
    new_n18502_, new_n18503_, new_n18504_, new_n18505_, new_n18506_,
    new_n18507_, new_n18508_, new_n18509_, new_n18510_, new_n18511_,
    new_n18512_, new_n18513_, new_n18514_, new_n18515_, new_n18516_,
    new_n18517_, new_n18518_, new_n18519_, new_n18520_, new_n18521_,
    new_n18522_, new_n18523_, new_n18524_, new_n18525_, new_n18526_,
    new_n18527_, new_n18528_, new_n18529_, new_n18530_, new_n18531_,
    new_n18532_, new_n18533_, new_n18534_, new_n18535_, new_n18536_,
    new_n18537_, new_n18538_, new_n18539_, new_n18540_, new_n18541_,
    new_n18542_, new_n18543_, new_n18544_, new_n18545_, new_n18546_,
    new_n18547_, new_n18548_, new_n18549_, new_n18550_, new_n18551_,
    new_n18552_, new_n18553_, new_n18554_, new_n18555_, new_n18556_,
    new_n18557_, new_n18558_, new_n18559_, new_n18560_, new_n18561_,
    new_n18562_, new_n18563_, new_n18564_, new_n18565_, new_n18566_,
    new_n18567_, new_n18568_, new_n18569_, new_n18570_, new_n18571_,
    new_n18572_, new_n18573_, new_n18574_, new_n18575_, new_n18576_,
    new_n18577_, new_n18578_, new_n18579_, new_n18580_, new_n18581_,
    new_n18582_, new_n18583_, new_n18584_, new_n18585_, new_n18586_,
    new_n18587_, new_n18588_, new_n18589_, new_n18591_, new_n18592_,
    new_n18593_, new_n18594_, new_n18595_, new_n18596_, new_n18597_,
    new_n18598_, new_n18599_, new_n18600_, new_n18601_, new_n18602_,
    new_n18603_, new_n18604_, new_n18605_, new_n18606_, new_n18607_,
    new_n18608_, new_n18609_, new_n18610_, new_n18611_, new_n18612_,
    new_n18613_, new_n18614_, new_n18615_, new_n18616_, new_n18617_,
    new_n18618_, new_n18619_, new_n18620_, new_n18621_, new_n18622_,
    new_n18623_, new_n18624_, new_n18625_, new_n18626_, new_n18627_,
    new_n18628_, new_n18629_, new_n18630_, new_n18631_, new_n18632_,
    new_n18633_, new_n18634_, new_n18635_, new_n18636_, new_n18637_,
    new_n18638_, new_n18639_, new_n18640_, new_n18641_, new_n18642_,
    new_n18643_, new_n18644_, new_n18645_, new_n18646_, new_n18647_,
    new_n18648_, new_n18649_, new_n18650_, new_n18651_, new_n18652_,
    new_n18653_, new_n18654_, new_n18655_, new_n18656_, new_n18657_,
    new_n18658_, new_n18659_, new_n18660_, new_n18661_, new_n18662_,
    new_n18663_, new_n18664_, new_n18665_, new_n18666_, new_n18667_,
    new_n18668_, new_n18669_, new_n18670_, new_n18671_, new_n18672_,
    new_n18673_, new_n18674_, new_n18675_, new_n18676_, new_n18677_,
    new_n18678_, new_n18679_, new_n18680_, new_n18681_, new_n18682_,
    new_n18683_, new_n18684_, new_n18685_, new_n18686_, new_n18687_,
    new_n18688_, new_n18689_, new_n18690_, new_n18691_, new_n18692_,
    new_n18693_, new_n18694_, new_n18695_, new_n18696_, new_n18697_,
    new_n18698_, new_n18699_, new_n18700_, new_n18701_, new_n18702_,
    new_n18703_, new_n18704_, new_n18705_, new_n18706_, new_n18707_,
    new_n18708_, new_n18709_, new_n18710_, new_n18711_, new_n18712_,
    new_n18713_, new_n18714_, new_n18715_, new_n18716_, new_n18717_,
    new_n18718_, new_n18719_, new_n18720_, new_n18721_, new_n18722_,
    new_n18723_, new_n18724_, new_n18725_, new_n18726_, new_n18727_,
    new_n18728_, new_n18729_, new_n18730_, new_n18731_, new_n18732_,
    new_n18733_, new_n18734_, new_n18735_, new_n18736_, new_n18737_,
    new_n18738_, new_n18739_, new_n18740_, new_n18741_, new_n18742_,
    new_n18743_, new_n18744_, new_n18745_, new_n18746_, new_n18747_,
    new_n18748_, new_n18749_, new_n18750_, new_n18751_, new_n18752_,
    new_n18753_, new_n18754_, new_n18755_, new_n18756_, new_n18757_,
    new_n18758_, new_n18759_, new_n18760_, new_n18761_, new_n18762_,
    new_n18763_, new_n18764_, new_n18765_, new_n18766_, new_n18767_,
    new_n18768_, new_n18769_, new_n18770_, new_n18771_, new_n18772_,
    new_n18773_, new_n18774_, new_n18775_, new_n18776_, new_n18777_,
    new_n18778_, new_n18779_, new_n18780_, new_n18781_, new_n18782_,
    new_n18783_, new_n18784_, new_n18785_, new_n18786_, new_n18787_,
    new_n18788_, new_n18789_, new_n18790_, new_n18791_, new_n18792_,
    new_n18793_, new_n18794_, new_n18795_, new_n18796_, new_n18797_,
    new_n18798_, new_n18799_, new_n18800_, new_n18801_, new_n18802_,
    new_n18803_, new_n18804_, new_n18805_, new_n18806_, new_n18807_,
    new_n18808_, new_n18809_, new_n18810_, new_n18811_, new_n18812_,
    new_n18813_, new_n18814_, new_n18815_, new_n18816_, new_n18817_,
    new_n18818_, new_n18819_, new_n18820_, new_n18821_, new_n18822_,
    new_n18823_, new_n18824_, new_n18825_, new_n18826_, new_n18827_,
    new_n18828_, new_n18829_, new_n18830_, new_n18831_, new_n18832_,
    new_n18833_, new_n18834_, new_n18835_, new_n18836_, new_n18837_,
    new_n18838_, new_n18839_, new_n18840_, new_n18841_, new_n18842_,
    new_n18843_, new_n18844_, new_n18845_, new_n18846_, new_n18847_,
    new_n18848_, new_n18849_, new_n18850_, new_n18851_, new_n18852_,
    new_n18853_, new_n18854_, new_n18855_, new_n18856_, new_n18857_,
    new_n18858_, new_n18859_, new_n18860_, new_n18861_, new_n18862_,
    new_n18863_, new_n18864_, new_n18865_, new_n18866_, new_n18867_,
    new_n18868_, new_n18869_, new_n18870_, new_n18871_, new_n18872_,
    new_n18873_, new_n18874_, new_n18875_, new_n18876_, new_n18877_,
    new_n18878_, new_n18879_, new_n18880_, new_n18881_, new_n18882_,
    new_n18883_, new_n18884_, new_n18885_, new_n18886_, new_n18887_,
    new_n18888_, new_n18889_, new_n18890_, new_n18891_, new_n18892_,
    new_n18893_, new_n18894_, new_n18895_, new_n18896_, new_n18897_,
    new_n18898_, new_n18899_, new_n18900_, new_n18901_, new_n18902_,
    new_n18903_, new_n18904_, new_n18905_, new_n18906_, new_n18907_,
    new_n18908_, new_n18909_, new_n18910_, new_n18911_, new_n18912_,
    new_n18913_, new_n18914_, new_n18915_, new_n18916_, new_n18917_,
    new_n18918_, new_n18919_, new_n18920_, new_n18921_, new_n18922_,
    new_n18923_, new_n18924_, new_n18925_, new_n18926_, new_n18927_,
    new_n18928_, new_n18929_, new_n18930_, new_n18931_, new_n18932_,
    new_n18933_, new_n18934_, new_n18935_, new_n18936_, new_n18937_,
    new_n18938_, new_n18939_, new_n18940_, new_n18941_, new_n18942_,
    new_n18943_, new_n18944_, new_n18945_, new_n18946_, new_n18947_,
    new_n18948_, new_n18949_, new_n18950_, new_n18951_, new_n18952_,
    new_n18953_, new_n18954_, new_n18955_, new_n18956_, new_n18957_,
    new_n18958_, new_n18959_, new_n18960_, new_n18961_, new_n18962_,
    new_n18963_, new_n18964_, new_n18965_, new_n18966_, new_n18967_,
    new_n18968_, new_n18969_, new_n18970_, new_n18971_, new_n18972_,
    new_n18973_, new_n18974_, new_n18975_, new_n18976_, new_n18977_,
    new_n18978_, new_n18979_, new_n18980_, new_n18981_, new_n18982_,
    new_n18983_, new_n18984_, new_n18985_, new_n18986_, new_n18987_,
    new_n18988_, new_n18989_, new_n18990_, new_n18991_, new_n18992_,
    new_n18993_, new_n18994_, new_n18995_, new_n18996_, new_n18997_,
    new_n18998_, new_n18999_, new_n19000_, new_n19001_, new_n19002_,
    new_n19003_, new_n19004_, new_n19005_, new_n19006_, new_n19007_,
    new_n19008_, new_n19009_, new_n19010_, new_n19011_, new_n19012_,
    new_n19013_, new_n19014_, new_n19015_, new_n19016_, new_n19017_,
    new_n19018_, new_n19019_, new_n19020_, new_n19021_, new_n19022_,
    new_n19023_, new_n19024_, new_n19025_, new_n19026_, new_n19027_,
    new_n19028_, new_n19029_, new_n19030_, new_n19031_, new_n19032_,
    new_n19033_, new_n19034_, new_n19035_, new_n19036_, new_n19037_,
    new_n19038_, new_n19039_, new_n19040_, new_n19041_, new_n19042_,
    new_n19043_, new_n19044_, new_n19045_, new_n19046_, new_n19047_,
    new_n19048_, new_n19049_, new_n19050_, new_n19051_, new_n19052_,
    new_n19053_, new_n19054_, new_n19055_, new_n19056_, new_n19057_,
    new_n19058_, new_n19059_, new_n19060_, new_n19061_, new_n19062_,
    new_n19063_, new_n19064_, new_n19065_, new_n19066_, new_n19067_,
    new_n19068_, new_n19069_, new_n19070_, new_n19071_, new_n19072_,
    new_n19073_, new_n19074_, new_n19075_, new_n19076_, new_n19077_,
    new_n19078_, new_n19079_, new_n19080_, new_n19081_, new_n19082_,
    new_n19083_, new_n19084_, new_n19085_, new_n19086_, new_n19087_,
    new_n19088_, new_n19089_, new_n19090_, new_n19091_, new_n19092_,
    new_n19093_, new_n19094_, new_n19095_, new_n19096_, new_n19097_,
    new_n19098_, new_n19099_, new_n19100_, new_n19101_, new_n19102_,
    new_n19103_, new_n19104_, new_n19105_, new_n19106_, new_n19107_,
    new_n19108_, new_n19109_, new_n19110_, new_n19111_, new_n19112_,
    new_n19113_, new_n19114_, new_n19115_, new_n19116_, new_n19117_,
    new_n19118_, new_n19119_, new_n19120_, new_n19121_, new_n19122_,
    new_n19123_, new_n19124_, new_n19125_, new_n19126_, new_n19127_,
    new_n19128_, new_n19129_, new_n19130_, new_n19131_, new_n19132_,
    new_n19133_, new_n19134_, new_n19135_, new_n19136_, new_n19137_,
    new_n19138_, new_n19139_, new_n19140_, new_n19141_, new_n19142_,
    new_n19143_, new_n19144_, new_n19145_, new_n19146_, new_n19147_,
    new_n19148_, new_n19149_, new_n19150_, new_n19151_, new_n19152_,
    new_n19153_, new_n19154_, new_n19155_, new_n19156_, new_n19157_,
    new_n19158_, new_n19159_, new_n19160_, new_n19161_, new_n19162_,
    new_n19163_, new_n19164_, new_n19165_, new_n19166_, new_n19167_,
    new_n19168_, new_n19169_, new_n19170_, new_n19171_, new_n19172_,
    new_n19173_, new_n19174_, new_n19175_, new_n19176_, new_n19177_,
    new_n19178_, new_n19179_, new_n19180_, new_n19181_, new_n19182_,
    new_n19183_, new_n19184_, new_n19185_, new_n19186_, new_n19187_,
    new_n19188_, new_n19189_, new_n19190_, new_n19191_, new_n19192_,
    new_n19193_, new_n19194_, new_n19195_, new_n19196_, new_n19197_,
    new_n19198_, new_n19199_, new_n19200_, new_n19201_, new_n19202_,
    new_n19203_, new_n19204_, new_n19205_, new_n19206_, new_n19207_,
    new_n19208_, new_n19209_, new_n19210_, new_n19211_, new_n19212_,
    new_n19213_, new_n19214_, new_n19215_, new_n19216_, new_n19217_,
    new_n19218_, new_n19219_, new_n19220_, new_n19221_, new_n19222_,
    new_n19223_, new_n19224_, new_n19225_, new_n19226_, new_n19227_,
    new_n19228_, new_n19229_, new_n19230_, new_n19231_, new_n19232_,
    new_n19233_, new_n19234_, new_n19235_, new_n19236_, new_n19237_,
    new_n19238_, new_n19239_, new_n19240_, new_n19241_, new_n19242_,
    new_n19243_, new_n19244_, new_n19245_, new_n19246_, new_n19247_,
    new_n19248_, new_n19249_, new_n19250_, new_n19251_, new_n19252_,
    new_n19253_, new_n19254_, new_n19255_, new_n19256_, new_n19257_,
    new_n19258_, new_n19259_, new_n19260_, new_n19261_, new_n19262_,
    new_n19263_, new_n19264_, new_n19265_, new_n19266_, new_n19267_,
    new_n19268_, new_n19269_, new_n19270_, new_n19271_, new_n19272_,
    new_n19273_, new_n19274_, new_n19275_, new_n19276_, new_n19277_,
    new_n19278_, new_n19279_, new_n19280_, new_n19281_, new_n19282_,
    new_n19283_, new_n19284_, new_n19285_, new_n19286_, new_n19287_,
    new_n19288_, new_n19289_, new_n19290_, new_n19291_, new_n19292_,
    new_n19293_, new_n19294_, new_n19295_, new_n19296_, new_n19297_,
    new_n19298_, new_n19299_, new_n19300_, new_n19301_, new_n19302_,
    new_n19303_, new_n19305_, new_n19306_, new_n19307_, new_n19308_,
    new_n19309_, new_n19310_, new_n19311_, new_n19312_, new_n19313_,
    new_n19314_, new_n19315_, new_n19316_, new_n19317_, new_n19318_,
    new_n19319_, new_n19320_, new_n19321_, new_n19322_, new_n19323_,
    new_n19324_, new_n19325_, new_n19326_, new_n19327_, new_n19328_,
    new_n19329_, new_n19330_, new_n19331_, new_n19332_, new_n19333_,
    new_n19334_, new_n19335_, new_n19336_, new_n19337_, new_n19338_,
    new_n19339_, new_n19340_, new_n19341_, new_n19342_, new_n19343_,
    new_n19344_, new_n19345_, new_n19346_, new_n19347_, new_n19348_,
    new_n19349_, new_n19350_, new_n19351_, new_n19352_, new_n19353_,
    new_n19354_, new_n19355_, new_n19356_, new_n19357_, new_n19358_,
    new_n19359_, new_n19360_, new_n19361_, new_n19362_, new_n19363_,
    new_n19364_, new_n19365_, new_n19366_, new_n19367_, new_n19368_,
    new_n19369_, new_n19370_, new_n19371_, new_n19372_, new_n19373_,
    new_n19374_, new_n19375_, new_n19376_, new_n19377_, new_n19378_,
    new_n19379_, new_n19380_, new_n19381_, new_n19382_, new_n19383_,
    new_n19384_, new_n19385_, new_n19386_, new_n19387_, new_n19388_,
    new_n19389_, new_n19390_, new_n19391_, new_n19392_, new_n19393_,
    new_n19394_, new_n19395_, new_n19396_, new_n19397_, new_n19398_,
    new_n19399_, new_n19400_, new_n19401_, new_n19402_, new_n19403_,
    new_n19404_, new_n19405_, new_n19406_, new_n19407_, new_n19408_,
    new_n19409_, new_n19410_, new_n19411_, new_n19412_, new_n19413_,
    new_n19414_, new_n19415_, new_n19416_, new_n19417_, new_n19418_,
    new_n19419_, new_n19420_, new_n19421_, new_n19422_, new_n19423_,
    new_n19424_, new_n19425_, new_n19426_, new_n19427_, new_n19428_,
    new_n19429_, new_n19430_, new_n19431_, new_n19432_, new_n19433_,
    new_n19434_, new_n19435_, new_n19436_, new_n19437_, new_n19438_,
    new_n19439_, new_n19440_, new_n19441_, new_n19442_, new_n19443_,
    new_n19444_, new_n19445_, new_n19446_, new_n19447_, new_n19448_,
    new_n19449_, new_n19450_, new_n19451_, new_n19452_, new_n19453_,
    new_n19454_, new_n19455_, new_n19456_, new_n19457_, new_n19458_,
    new_n19459_, new_n19460_, new_n19461_, new_n19462_, new_n19463_,
    new_n19464_, new_n19465_, new_n19466_, new_n19467_, new_n19468_,
    new_n19469_, new_n19470_, new_n19471_, new_n19472_, new_n19473_,
    new_n19474_, new_n19475_, new_n19476_, new_n19477_, new_n19478_,
    new_n19479_, new_n19480_, new_n19481_, new_n19482_, new_n19483_,
    new_n19484_, new_n19485_, new_n19486_, new_n19487_, new_n19488_,
    new_n19489_, new_n19490_, new_n19491_, new_n19492_, new_n19493_,
    new_n19494_, new_n19495_, new_n19496_, new_n19497_, new_n19498_,
    new_n19499_, new_n19500_, new_n19501_, new_n19502_, new_n19503_,
    new_n19504_, new_n19505_, new_n19506_, new_n19507_, new_n19508_,
    new_n19509_, new_n19510_, new_n19511_, new_n19512_, new_n19513_,
    new_n19514_, new_n19515_, new_n19516_, new_n19517_, new_n19518_,
    new_n19519_, new_n19520_, new_n19521_, new_n19522_, new_n19523_,
    new_n19524_, new_n19525_, new_n19526_, new_n19527_, new_n19528_,
    new_n19529_, new_n19530_, new_n19531_, new_n19532_, new_n19533_,
    new_n19534_, new_n19535_, new_n19536_, new_n19537_, new_n19538_,
    new_n19539_, new_n19540_, new_n19541_, new_n19542_, new_n19543_,
    new_n19544_, new_n19545_, new_n19546_, new_n19547_, new_n19548_,
    new_n19549_, new_n19550_, new_n19551_, new_n19552_, new_n19553_,
    new_n19554_, new_n19555_, new_n19556_, new_n19557_, new_n19558_,
    new_n19559_, new_n19560_, new_n19561_, new_n19562_, new_n19563_,
    new_n19564_, new_n19565_, new_n19566_, new_n19567_, new_n19568_,
    new_n19569_, new_n19570_, new_n19571_, new_n19572_, new_n19573_,
    new_n19574_, new_n19575_, new_n19576_, new_n19577_, new_n19578_,
    new_n19579_, new_n19580_, new_n19581_, new_n19582_, new_n19583_,
    new_n19584_, new_n19585_, new_n19586_, new_n19587_, new_n19588_,
    new_n19589_, new_n19590_, new_n19591_, new_n19592_, new_n19593_,
    new_n19594_, new_n19595_, new_n19596_, new_n19597_, new_n19598_,
    new_n19599_, new_n19600_, new_n19601_, new_n19602_, new_n19603_,
    new_n19604_, new_n19605_, new_n19606_, new_n19607_, new_n19608_,
    new_n19609_, new_n19610_, new_n19611_, new_n19612_, new_n19613_,
    new_n19614_, new_n19615_, new_n19616_, new_n19617_, new_n19618_,
    new_n19619_, new_n19620_, new_n19621_, new_n19622_, new_n19623_,
    new_n19624_, new_n19625_, new_n19626_, new_n19627_, new_n19628_,
    new_n19629_, new_n19630_, new_n19631_, new_n19632_, new_n19633_,
    new_n19634_, new_n19635_, new_n19636_, new_n19637_, new_n19638_,
    new_n19639_, new_n19640_, new_n19641_, new_n19642_, new_n19643_,
    new_n19644_, new_n19645_, new_n19646_, new_n19647_, new_n19648_,
    new_n19649_, new_n19650_, new_n19651_, new_n19652_, new_n19653_,
    new_n19654_, new_n19655_, new_n19656_, new_n19657_, new_n19658_,
    new_n19659_, new_n19660_, new_n19661_, new_n19662_, new_n19663_,
    new_n19664_, new_n19665_, new_n19666_, new_n19667_, new_n19668_,
    new_n19669_, new_n19670_, new_n19671_, new_n19672_, new_n19673_,
    new_n19674_, new_n19675_, new_n19676_, new_n19677_, new_n19678_,
    new_n19679_, new_n19680_, new_n19681_, new_n19682_, new_n19683_,
    new_n19684_, new_n19685_, new_n19686_, new_n19687_, new_n19688_,
    new_n19689_, new_n19690_, new_n19691_, new_n19692_, new_n19693_,
    new_n19694_, new_n19695_, new_n19696_, new_n19697_, new_n19698_,
    new_n19699_, new_n19700_, new_n19701_, new_n19702_, new_n19703_,
    new_n19704_, new_n19705_, new_n19706_, new_n19707_, new_n19708_,
    new_n19709_, new_n19710_, new_n19711_, new_n19712_, new_n19713_,
    new_n19714_, new_n19715_, new_n19716_, new_n19717_, new_n19718_,
    new_n19719_, new_n19720_, new_n19721_, new_n19722_, new_n19723_,
    new_n19724_, new_n19725_, new_n19726_, new_n19727_, new_n19728_,
    new_n19729_, new_n19730_, new_n19731_, new_n19732_, new_n19733_,
    new_n19734_, new_n19735_, new_n19736_, new_n19737_, new_n19738_,
    new_n19739_, new_n19740_, new_n19741_, new_n19742_, new_n19743_,
    new_n19744_, new_n19745_, new_n19746_, new_n19747_, new_n19748_,
    new_n19749_, new_n19750_, new_n19751_, new_n19752_, new_n19753_,
    new_n19754_, new_n19755_, new_n19756_, new_n19757_, new_n19758_,
    new_n19759_, new_n19760_, new_n19761_, new_n19762_, new_n19763_,
    new_n19764_, new_n19765_, new_n19766_, new_n19767_, new_n19768_,
    new_n19769_, new_n19770_, new_n19771_, new_n19772_, new_n19773_,
    new_n19774_, new_n19775_, new_n19776_, new_n19777_, new_n19778_,
    new_n19779_, new_n19780_, new_n19781_, new_n19782_, new_n19783_,
    new_n19784_, new_n19785_, new_n19786_, new_n19787_, new_n19788_,
    new_n19789_, new_n19790_, new_n19791_, new_n19792_, new_n19793_,
    new_n19794_, new_n19795_, new_n19796_, new_n19797_, new_n19798_,
    new_n19799_, new_n19800_, new_n19801_, new_n19802_, new_n19803_,
    new_n19804_, new_n19805_, new_n19806_, new_n19807_, new_n19808_,
    new_n19809_, new_n19810_, new_n19811_, new_n19812_, new_n19813_,
    new_n19814_, new_n19815_, new_n19816_, new_n19817_, new_n19818_,
    new_n19819_, new_n19820_, new_n19821_, new_n19822_, new_n19823_,
    new_n19824_, new_n19825_, new_n19826_, new_n19827_, new_n19828_,
    new_n19829_, new_n19830_, new_n19831_, new_n19832_, new_n19833_,
    new_n19834_, new_n19835_, new_n19836_, new_n19837_, new_n19838_,
    new_n19839_, new_n19840_, new_n19841_, new_n19842_, new_n19843_,
    new_n19844_, new_n19845_, new_n19846_, new_n19847_, new_n19848_,
    new_n19849_, new_n19850_, new_n19851_, new_n19852_, new_n19853_,
    new_n19854_, new_n19855_, new_n19856_, new_n19857_, new_n19858_,
    new_n19859_, new_n19860_, new_n19861_, new_n19862_, new_n19863_,
    new_n19864_, new_n19865_, new_n19866_, new_n19867_, new_n19868_,
    new_n19869_, new_n19870_, new_n19871_, new_n19872_, new_n19873_,
    new_n19874_, new_n19875_, new_n19876_, new_n19877_, new_n19878_,
    new_n19879_, new_n19880_, new_n19881_, new_n19882_, new_n19883_,
    new_n19884_, new_n19885_, new_n19886_, new_n19887_, new_n19888_,
    new_n19889_, new_n19890_, new_n19891_, new_n19892_, new_n19893_,
    new_n19894_, new_n19895_, new_n19896_, new_n19897_, new_n19898_,
    new_n19899_, new_n19900_, new_n19901_, new_n19902_, new_n19903_,
    new_n19904_, new_n19905_, new_n19906_, new_n19907_, new_n19908_,
    new_n19909_, new_n19910_, new_n19911_, new_n19912_, new_n19913_,
    new_n19914_, new_n19915_, new_n19916_, new_n19917_, new_n19918_,
    new_n19919_, new_n19920_, new_n19921_, new_n19922_, new_n19923_,
    new_n19924_, new_n19925_, new_n19926_, new_n19927_, new_n19928_,
    new_n19929_, new_n19930_, new_n19931_, new_n19932_, new_n19933_,
    new_n19934_, new_n19935_, new_n19936_, new_n19937_, new_n19938_,
    new_n19939_, new_n19940_, new_n19941_, new_n19942_, new_n19943_,
    new_n19944_, new_n19945_, new_n19946_, new_n19947_, new_n19948_,
    new_n19949_, new_n19950_, new_n19951_, new_n19952_, new_n19953_,
    new_n19954_, new_n19955_, new_n19956_, new_n19957_, new_n19958_,
    new_n19959_, new_n19960_, new_n19961_, new_n19962_, new_n19963_,
    new_n19964_, new_n19965_, new_n19966_, new_n19967_, new_n19968_,
    new_n19969_, new_n19970_, new_n19971_, new_n19972_, new_n19973_,
    new_n19974_, new_n19975_, new_n19976_, new_n19977_, new_n19978_,
    new_n19979_, new_n19980_, new_n19981_, new_n19982_, new_n19983_,
    new_n19984_, new_n19985_, new_n19986_, new_n19987_, new_n19988_,
    new_n19989_, new_n19990_, new_n19991_, new_n19992_, new_n19993_,
    new_n19994_, new_n19995_, new_n19996_, new_n19997_, new_n19998_,
    new_n19999_, new_n20000_, new_n20001_, new_n20002_, new_n20003_,
    new_n20004_, new_n20005_, new_n20006_, new_n20007_, new_n20008_,
    new_n20009_, new_n20010_, new_n20011_, new_n20012_, new_n20013_,
    new_n20014_, new_n20015_, new_n20016_, new_n20017_, new_n20018_,
    new_n20019_, new_n20020_, new_n20021_, new_n20022_, new_n20023_,
    new_n20024_, new_n20025_, new_n20026_, new_n20027_, new_n20028_,
    new_n20029_, new_n20030_, new_n20031_, new_n20032_, new_n20033_,
    new_n20034_, new_n20036_, new_n20037_, new_n20038_, new_n20039_,
    new_n20040_, new_n20041_, new_n20042_, new_n20043_, new_n20044_,
    new_n20045_, new_n20046_, new_n20047_, new_n20048_, new_n20049_,
    new_n20050_, new_n20051_, new_n20052_, new_n20053_, new_n20054_,
    new_n20055_, new_n20056_, new_n20057_, new_n20058_, new_n20059_,
    new_n20060_, new_n20061_, new_n20062_, new_n20063_, new_n20064_,
    new_n20065_, new_n20066_, new_n20067_, new_n20068_, new_n20069_,
    new_n20070_, new_n20071_, new_n20072_, new_n20073_, new_n20074_,
    new_n20075_, new_n20076_, new_n20077_, new_n20078_, new_n20079_,
    new_n20080_, new_n20081_, new_n20082_, new_n20083_, new_n20084_,
    new_n20085_, new_n20086_, new_n20087_, new_n20088_, new_n20089_,
    new_n20090_, new_n20091_, new_n20092_, new_n20093_, new_n20094_,
    new_n20095_, new_n20096_, new_n20097_, new_n20098_, new_n20099_,
    new_n20100_, new_n20101_, new_n20102_, new_n20103_, new_n20104_,
    new_n20105_, new_n20106_, new_n20107_, new_n20108_, new_n20109_,
    new_n20110_, new_n20111_, new_n20112_, new_n20113_, new_n20114_,
    new_n20115_, new_n20116_, new_n20117_, new_n20118_, new_n20119_,
    new_n20120_, new_n20121_, new_n20122_, new_n20123_, new_n20124_,
    new_n20125_, new_n20126_, new_n20127_, new_n20128_, new_n20129_,
    new_n20130_, new_n20131_, new_n20132_, new_n20133_, new_n20134_,
    new_n20135_, new_n20136_, new_n20137_, new_n20138_, new_n20139_,
    new_n20140_, new_n20141_, new_n20142_, new_n20143_, new_n20144_,
    new_n20145_, new_n20146_, new_n20147_, new_n20148_, new_n20149_,
    new_n20150_, new_n20151_, new_n20152_, new_n20153_, new_n20154_,
    new_n20155_, new_n20156_, new_n20157_, new_n20158_, new_n20159_,
    new_n20160_, new_n20161_, new_n20162_, new_n20163_, new_n20164_,
    new_n20165_, new_n20166_, new_n20167_, new_n20168_, new_n20169_,
    new_n20170_, new_n20171_, new_n20172_, new_n20173_, new_n20174_,
    new_n20175_, new_n20176_, new_n20177_, new_n20178_, new_n20179_,
    new_n20180_, new_n20181_, new_n20182_, new_n20183_, new_n20184_,
    new_n20185_, new_n20186_, new_n20187_, new_n20188_, new_n20189_,
    new_n20190_, new_n20191_, new_n20192_, new_n20193_, new_n20194_,
    new_n20195_, new_n20196_, new_n20197_, new_n20198_, new_n20199_,
    new_n20200_, new_n20201_, new_n20202_, new_n20203_, new_n20204_,
    new_n20205_, new_n20206_, new_n20207_, new_n20208_, new_n20209_,
    new_n20210_, new_n20211_, new_n20212_, new_n20213_, new_n20214_,
    new_n20215_, new_n20216_, new_n20217_, new_n20218_, new_n20219_,
    new_n20220_, new_n20221_, new_n20222_, new_n20223_, new_n20224_,
    new_n20225_, new_n20226_, new_n20227_, new_n20228_, new_n20229_,
    new_n20230_, new_n20231_, new_n20232_, new_n20233_, new_n20234_,
    new_n20235_, new_n20236_, new_n20237_, new_n20238_, new_n20239_,
    new_n20240_, new_n20241_, new_n20242_, new_n20243_, new_n20244_,
    new_n20245_, new_n20246_, new_n20247_, new_n20248_, new_n20249_,
    new_n20250_, new_n20251_, new_n20252_, new_n20253_, new_n20254_,
    new_n20255_, new_n20256_, new_n20257_, new_n20258_, new_n20259_,
    new_n20260_, new_n20261_, new_n20262_, new_n20263_, new_n20264_,
    new_n20265_, new_n20266_, new_n20267_, new_n20268_, new_n20269_,
    new_n20270_, new_n20271_, new_n20272_, new_n20273_, new_n20274_,
    new_n20275_, new_n20276_, new_n20277_, new_n20278_, new_n20279_,
    new_n20280_, new_n20281_, new_n20282_, new_n20283_, new_n20284_,
    new_n20285_, new_n20286_, new_n20287_, new_n20288_, new_n20289_,
    new_n20290_, new_n20291_, new_n20292_, new_n20293_, new_n20294_,
    new_n20295_, new_n20296_, new_n20297_, new_n20298_, new_n20299_,
    new_n20300_, new_n20301_, new_n20302_, new_n20303_, new_n20304_,
    new_n20305_, new_n20306_, new_n20307_, new_n20308_, new_n20309_,
    new_n20310_, new_n20311_, new_n20312_, new_n20313_, new_n20314_,
    new_n20315_, new_n20316_, new_n20317_, new_n20318_, new_n20319_,
    new_n20320_, new_n20321_, new_n20322_, new_n20323_, new_n20324_,
    new_n20325_, new_n20326_, new_n20327_, new_n20328_, new_n20329_,
    new_n20330_, new_n20331_, new_n20332_, new_n20333_, new_n20334_,
    new_n20335_, new_n20336_, new_n20337_, new_n20338_, new_n20339_,
    new_n20340_, new_n20341_, new_n20342_, new_n20343_, new_n20344_,
    new_n20345_, new_n20346_, new_n20347_, new_n20348_, new_n20349_,
    new_n20350_, new_n20351_, new_n20352_, new_n20353_, new_n20354_,
    new_n20355_, new_n20356_, new_n20357_, new_n20358_, new_n20359_,
    new_n20360_, new_n20361_, new_n20362_, new_n20363_, new_n20364_,
    new_n20365_, new_n20366_, new_n20367_, new_n20368_, new_n20369_,
    new_n20370_, new_n20371_, new_n20372_, new_n20373_, new_n20374_,
    new_n20375_, new_n20376_, new_n20377_, new_n20378_, new_n20379_,
    new_n20380_, new_n20381_, new_n20382_, new_n20383_, new_n20384_,
    new_n20385_, new_n20386_, new_n20387_, new_n20388_, new_n20389_,
    new_n20390_, new_n20391_, new_n20392_, new_n20393_, new_n20394_,
    new_n20395_, new_n20396_, new_n20397_, new_n20398_, new_n20399_,
    new_n20400_, new_n20401_, new_n20402_, new_n20403_, new_n20404_,
    new_n20405_, new_n20406_, new_n20407_, new_n20408_, new_n20409_,
    new_n20410_, new_n20411_, new_n20412_, new_n20413_, new_n20414_,
    new_n20415_, new_n20416_, new_n20417_, new_n20418_, new_n20419_,
    new_n20420_, new_n20421_, new_n20422_, new_n20423_, new_n20424_,
    new_n20425_, new_n20426_, new_n20427_, new_n20428_, new_n20429_,
    new_n20430_, new_n20431_, new_n20432_, new_n20433_, new_n20434_,
    new_n20435_, new_n20436_, new_n20437_, new_n20438_, new_n20439_,
    new_n20440_, new_n20441_, new_n20442_, new_n20443_, new_n20444_,
    new_n20445_, new_n20446_, new_n20447_, new_n20448_, new_n20449_,
    new_n20450_, new_n20451_, new_n20452_, new_n20453_, new_n20454_,
    new_n20455_, new_n20456_, new_n20457_, new_n20458_, new_n20459_,
    new_n20460_, new_n20461_, new_n20462_, new_n20463_, new_n20464_,
    new_n20465_, new_n20466_, new_n20467_, new_n20468_, new_n20469_,
    new_n20470_, new_n20471_, new_n20472_, new_n20473_, new_n20474_,
    new_n20475_, new_n20476_, new_n20477_, new_n20478_, new_n20479_,
    new_n20480_, new_n20481_, new_n20482_, new_n20483_, new_n20484_,
    new_n20485_, new_n20486_, new_n20487_, new_n20488_, new_n20489_,
    new_n20490_, new_n20491_, new_n20492_, new_n20493_, new_n20494_,
    new_n20495_, new_n20496_, new_n20497_, new_n20498_, new_n20499_,
    new_n20500_, new_n20501_, new_n20502_, new_n20503_, new_n20504_,
    new_n20505_, new_n20506_, new_n20507_, new_n20508_, new_n20509_,
    new_n20510_, new_n20511_, new_n20512_, new_n20513_, new_n20514_,
    new_n20515_, new_n20516_, new_n20517_, new_n20518_, new_n20519_,
    new_n20520_, new_n20521_, new_n20522_, new_n20523_, new_n20524_,
    new_n20525_, new_n20526_, new_n20527_, new_n20528_, new_n20529_,
    new_n20530_, new_n20531_, new_n20532_, new_n20533_, new_n20534_,
    new_n20535_, new_n20536_, new_n20537_, new_n20538_, new_n20539_,
    new_n20540_, new_n20541_, new_n20542_, new_n20543_, new_n20544_,
    new_n20545_, new_n20546_, new_n20547_, new_n20548_, new_n20549_,
    new_n20550_, new_n20551_, new_n20552_, new_n20553_, new_n20554_,
    new_n20555_, new_n20556_, new_n20557_, new_n20558_, new_n20559_,
    new_n20560_, new_n20561_, new_n20562_, new_n20563_, new_n20564_,
    new_n20565_, new_n20566_, new_n20567_, new_n20568_, new_n20569_,
    new_n20570_, new_n20571_, new_n20572_, new_n20573_, new_n20574_,
    new_n20575_, new_n20576_, new_n20577_, new_n20578_, new_n20579_,
    new_n20580_, new_n20581_, new_n20582_, new_n20583_, new_n20584_,
    new_n20585_, new_n20586_, new_n20587_, new_n20588_, new_n20589_,
    new_n20590_, new_n20591_, new_n20592_, new_n20593_, new_n20594_,
    new_n20595_, new_n20596_, new_n20597_, new_n20598_, new_n20599_,
    new_n20600_, new_n20601_, new_n20602_, new_n20603_, new_n20604_,
    new_n20605_, new_n20606_, new_n20607_, new_n20608_, new_n20609_,
    new_n20610_, new_n20611_, new_n20612_, new_n20613_, new_n20614_,
    new_n20615_, new_n20616_, new_n20617_, new_n20618_, new_n20619_,
    new_n20620_, new_n20621_, new_n20622_, new_n20623_, new_n20624_,
    new_n20625_, new_n20626_, new_n20627_, new_n20628_, new_n20629_,
    new_n20630_, new_n20631_, new_n20632_, new_n20633_, new_n20634_,
    new_n20635_, new_n20636_, new_n20637_, new_n20638_, new_n20639_,
    new_n20640_, new_n20641_, new_n20642_, new_n20643_, new_n20644_,
    new_n20645_, new_n20646_, new_n20647_, new_n20648_, new_n20649_,
    new_n20650_, new_n20651_, new_n20652_, new_n20653_, new_n20654_,
    new_n20655_, new_n20656_, new_n20657_, new_n20658_, new_n20659_,
    new_n20660_, new_n20661_, new_n20662_, new_n20663_, new_n20664_,
    new_n20665_, new_n20666_, new_n20667_, new_n20668_, new_n20669_,
    new_n20670_, new_n20671_, new_n20672_, new_n20673_, new_n20674_,
    new_n20675_, new_n20676_, new_n20677_, new_n20678_, new_n20679_,
    new_n20680_, new_n20681_, new_n20682_, new_n20683_, new_n20684_,
    new_n20685_, new_n20686_, new_n20687_, new_n20688_, new_n20689_,
    new_n20690_, new_n20691_, new_n20692_, new_n20693_, new_n20694_,
    new_n20695_, new_n20696_, new_n20697_, new_n20698_, new_n20699_,
    new_n20700_, new_n20701_, new_n20702_, new_n20703_, new_n20704_,
    new_n20705_, new_n20706_, new_n20707_, new_n20708_, new_n20709_,
    new_n20710_, new_n20711_, new_n20712_, new_n20713_, new_n20714_,
    new_n20715_, new_n20716_, new_n20717_, new_n20718_, new_n20719_,
    new_n20720_, new_n20721_, new_n20722_, new_n20723_, new_n20724_,
    new_n20725_, new_n20726_, new_n20727_, new_n20728_, new_n20729_,
    new_n20730_, new_n20731_, new_n20732_, new_n20733_, new_n20734_,
    new_n20735_, new_n20736_, new_n20737_, new_n20738_, new_n20739_,
    new_n20740_, new_n20741_, new_n20742_, new_n20743_, new_n20744_,
    new_n20745_, new_n20746_, new_n20747_, new_n20748_, new_n20749_,
    new_n20750_, new_n20751_, new_n20752_, new_n20753_, new_n20754_,
    new_n20755_, new_n20756_, new_n20757_, new_n20758_, new_n20759_,
    new_n20760_, new_n20761_, new_n20762_, new_n20763_, new_n20764_,
    new_n20765_, new_n20766_, new_n20767_, new_n20768_, new_n20769_,
    new_n20770_, new_n20771_, new_n20772_, new_n20773_, new_n20774_,
    new_n20775_, new_n20776_, new_n20777_, new_n20778_, new_n20779_,
    new_n20781_, new_n20782_, new_n20783_, new_n20784_, new_n20785_,
    new_n20786_, new_n20787_, new_n20788_, new_n20789_, new_n20790_,
    new_n20791_, new_n20792_, new_n20793_, new_n20794_, new_n20795_,
    new_n20796_, new_n20797_, new_n20798_, new_n20799_, new_n20800_,
    new_n20801_, new_n20802_, new_n20803_, new_n20804_, new_n20805_,
    new_n20806_, new_n20807_, new_n20808_, new_n20809_, new_n20810_,
    new_n20811_, new_n20812_, new_n20813_, new_n20814_, new_n20815_,
    new_n20816_, new_n20817_, new_n20818_, new_n20819_, new_n20820_,
    new_n20821_, new_n20822_, new_n20823_, new_n20824_, new_n20825_,
    new_n20826_, new_n20827_, new_n20828_, new_n20829_, new_n20830_,
    new_n20831_, new_n20832_, new_n20833_, new_n20834_, new_n20835_,
    new_n20836_, new_n20837_, new_n20838_, new_n20839_, new_n20840_,
    new_n20841_, new_n20842_, new_n20843_, new_n20844_, new_n20845_,
    new_n20846_, new_n20847_, new_n20848_, new_n20849_, new_n20850_,
    new_n20851_, new_n20852_, new_n20853_, new_n20854_, new_n20855_,
    new_n20856_, new_n20857_, new_n20858_, new_n20859_, new_n20860_,
    new_n20861_, new_n20862_, new_n20863_, new_n20864_, new_n20865_,
    new_n20866_, new_n20867_, new_n20868_, new_n20869_, new_n20870_,
    new_n20871_, new_n20872_, new_n20873_, new_n20874_, new_n20875_,
    new_n20876_, new_n20877_, new_n20878_, new_n20879_, new_n20880_,
    new_n20881_, new_n20882_, new_n20883_, new_n20884_, new_n20885_,
    new_n20886_, new_n20887_, new_n20888_, new_n20889_, new_n20890_,
    new_n20891_, new_n20892_, new_n20893_, new_n20894_, new_n20895_,
    new_n20896_, new_n20897_, new_n20898_, new_n20899_, new_n20900_,
    new_n20901_, new_n20902_, new_n20903_, new_n20904_, new_n20905_,
    new_n20906_, new_n20907_, new_n20908_, new_n20909_, new_n20910_,
    new_n20911_, new_n20912_, new_n20913_, new_n20914_, new_n20915_,
    new_n20916_, new_n20917_, new_n20918_, new_n20919_, new_n20920_,
    new_n20921_, new_n20922_, new_n20923_, new_n20924_, new_n20925_,
    new_n20926_, new_n20927_, new_n20928_, new_n20929_, new_n20930_,
    new_n20931_, new_n20932_, new_n20933_, new_n20934_, new_n20935_,
    new_n20936_, new_n20937_, new_n20938_, new_n20939_, new_n20940_,
    new_n20941_, new_n20942_, new_n20943_, new_n20944_, new_n20945_,
    new_n20946_, new_n20947_, new_n20948_, new_n20949_, new_n20950_,
    new_n20951_, new_n20952_, new_n20953_, new_n20954_, new_n20955_,
    new_n20956_, new_n20957_, new_n20958_, new_n20959_, new_n20960_,
    new_n20961_, new_n20962_, new_n20963_, new_n20964_, new_n20965_,
    new_n20966_, new_n20967_, new_n20968_, new_n20969_, new_n20970_,
    new_n20971_, new_n20972_, new_n20973_, new_n20974_, new_n20975_,
    new_n20976_, new_n20977_, new_n20978_, new_n20979_, new_n20980_,
    new_n20981_, new_n20982_, new_n20983_, new_n20984_, new_n20985_,
    new_n20986_, new_n20987_, new_n20988_, new_n20989_, new_n20990_,
    new_n20991_, new_n20992_, new_n20993_, new_n20994_, new_n20995_,
    new_n20996_, new_n20997_, new_n20998_, new_n20999_, new_n21000_,
    new_n21001_, new_n21002_, new_n21003_, new_n21004_, new_n21005_,
    new_n21006_, new_n21007_, new_n21008_, new_n21009_, new_n21010_,
    new_n21011_, new_n21012_, new_n21013_, new_n21014_, new_n21015_,
    new_n21016_, new_n21017_, new_n21018_, new_n21019_, new_n21020_,
    new_n21021_, new_n21022_, new_n21023_, new_n21024_, new_n21025_,
    new_n21026_, new_n21027_, new_n21028_, new_n21029_, new_n21030_,
    new_n21031_, new_n21032_, new_n21033_, new_n21034_, new_n21035_,
    new_n21036_, new_n21037_, new_n21038_, new_n21039_, new_n21040_,
    new_n21041_, new_n21042_, new_n21043_, new_n21044_, new_n21045_,
    new_n21046_, new_n21047_, new_n21048_, new_n21049_, new_n21050_,
    new_n21051_, new_n21052_, new_n21053_, new_n21054_, new_n21055_,
    new_n21056_, new_n21057_, new_n21058_, new_n21059_, new_n21060_,
    new_n21061_, new_n21062_, new_n21063_, new_n21064_, new_n21065_,
    new_n21066_, new_n21067_, new_n21068_, new_n21069_, new_n21070_,
    new_n21071_, new_n21072_, new_n21073_, new_n21074_, new_n21075_,
    new_n21076_, new_n21077_, new_n21078_, new_n21079_, new_n21080_,
    new_n21081_, new_n21082_, new_n21083_, new_n21084_, new_n21085_,
    new_n21086_, new_n21087_, new_n21088_, new_n21089_, new_n21090_,
    new_n21091_, new_n21092_, new_n21093_, new_n21094_, new_n21095_,
    new_n21096_, new_n21097_, new_n21098_, new_n21099_, new_n21100_,
    new_n21101_, new_n21102_, new_n21103_, new_n21104_, new_n21105_,
    new_n21106_, new_n21107_, new_n21108_, new_n21109_, new_n21110_,
    new_n21111_, new_n21112_, new_n21113_, new_n21114_, new_n21115_,
    new_n21116_, new_n21117_, new_n21118_, new_n21119_, new_n21120_,
    new_n21121_, new_n21122_, new_n21123_, new_n21124_, new_n21125_,
    new_n21126_, new_n21127_, new_n21128_, new_n21129_, new_n21130_,
    new_n21131_, new_n21132_, new_n21133_, new_n21134_, new_n21135_,
    new_n21136_, new_n21137_, new_n21138_, new_n21139_, new_n21140_,
    new_n21141_, new_n21142_, new_n21143_, new_n21144_, new_n21145_,
    new_n21146_, new_n21147_, new_n21148_, new_n21149_, new_n21150_,
    new_n21151_, new_n21152_, new_n21153_, new_n21154_, new_n21155_,
    new_n21156_, new_n21157_, new_n21158_, new_n21159_, new_n21160_,
    new_n21161_, new_n21162_, new_n21163_, new_n21164_, new_n21165_,
    new_n21166_, new_n21167_, new_n21168_, new_n21169_, new_n21170_,
    new_n21171_, new_n21172_, new_n21173_, new_n21174_, new_n21175_,
    new_n21176_, new_n21177_, new_n21178_, new_n21179_, new_n21180_,
    new_n21181_, new_n21182_, new_n21183_, new_n21184_, new_n21185_,
    new_n21186_, new_n21187_, new_n21188_, new_n21189_, new_n21190_,
    new_n21191_, new_n21192_, new_n21193_, new_n21194_, new_n21195_,
    new_n21196_, new_n21197_, new_n21198_, new_n21199_, new_n21200_,
    new_n21201_, new_n21202_, new_n21203_, new_n21204_, new_n21205_,
    new_n21206_, new_n21207_, new_n21208_, new_n21209_, new_n21210_,
    new_n21211_, new_n21212_, new_n21213_, new_n21214_, new_n21215_,
    new_n21216_, new_n21217_, new_n21218_, new_n21219_, new_n21220_,
    new_n21221_, new_n21222_, new_n21223_, new_n21224_, new_n21225_,
    new_n21226_, new_n21227_, new_n21228_, new_n21229_, new_n21230_,
    new_n21231_, new_n21232_, new_n21233_, new_n21234_, new_n21235_,
    new_n21236_, new_n21237_, new_n21238_, new_n21239_, new_n21240_,
    new_n21241_, new_n21242_, new_n21243_, new_n21244_, new_n21245_,
    new_n21246_, new_n21247_, new_n21248_, new_n21249_, new_n21250_,
    new_n21251_, new_n21252_, new_n21253_, new_n21254_, new_n21255_,
    new_n21256_, new_n21257_, new_n21258_, new_n21259_, new_n21260_,
    new_n21261_, new_n21262_, new_n21263_, new_n21264_, new_n21265_,
    new_n21266_, new_n21267_, new_n21268_, new_n21269_, new_n21270_,
    new_n21271_, new_n21272_, new_n21273_, new_n21274_, new_n21275_,
    new_n21276_, new_n21277_, new_n21278_, new_n21279_, new_n21280_,
    new_n21281_, new_n21282_, new_n21283_, new_n21284_, new_n21285_,
    new_n21286_, new_n21287_, new_n21288_, new_n21289_, new_n21290_,
    new_n21291_, new_n21292_, new_n21293_, new_n21294_, new_n21295_,
    new_n21296_, new_n21297_, new_n21298_, new_n21299_, new_n21300_,
    new_n21301_, new_n21302_, new_n21303_, new_n21304_, new_n21305_,
    new_n21306_, new_n21307_, new_n21308_, new_n21309_, new_n21310_,
    new_n21311_, new_n21312_, new_n21313_, new_n21314_, new_n21315_,
    new_n21316_, new_n21317_, new_n21318_, new_n21319_, new_n21320_,
    new_n21321_, new_n21322_, new_n21323_, new_n21324_, new_n21325_,
    new_n21326_, new_n21327_, new_n21328_, new_n21329_, new_n21330_,
    new_n21331_, new_n21332_, new_n21333_, new_n21334_, new_n21335_,
    new_n21336_, new_n21337_, new_n21338_, new_n21339_, new_n21340_,
    new_n21341_, new_n21342_, new_n21343_, new_n21344_, new_n21345_,
    new_n21346_, new_n21347_, new_n21348_, new_n21349_, new_n21350_,
    new_n21351_, new_n21352_, new_n21353_, new_n21354_, new_n21355_,
    new_n21356_, new_n21357_, new_n21358_, new_n21359_, new_n21360_,
    new_n21361_, new_n21362_, new_n21363_, new_n21364_, new_n21365_,
    new_n21366_, new_n21367_, new_n21368_, new_n21369_, new_n21370_,
    new_n21371_, new_n21372_, new_n21373_, new_n21374_, new_n21375_,
    new_n21376_, new_n21377_, new_n21378_, new_n21379_, new_n21380_,
    new_n21381_, new_n21382_, new_n21383_, new_n21384_, new_n21385_,
    new_n21386_, new_n21387_, new_n21388_, new_n21389_, new_n21390_,
    new_n21391_, new_n21392_, new_n21393_, new_n21394_, new_n21395_,
    new_n21396_, new_n21397_, new_n21398_, new_n21399_, new_n21400_,
    new_n21401_, new_n21402_, new_n21403_, new_n21404_, new_n21405_,
    new_n21406_, new_n21407_, new_n21408_, new_n21409_, new_n21410_,
    new_n21411_, new_n21412_, new_n21413_, new_n21414_, new_n21415_,
    new_n21416_, new_n21417_, new_n21418_, new_n21419_, new_n21420_,
    new_n21421_, new_n21422_, new_n21423_, new_n21424_, new_n21425_,
    new_n21426_, new_n21427_, new_n21428_, new_n21429_, new_n21430_,
    new_n21431_, new_n21432_, new_n21433_, new_n21434_, new_n21435_,
    new_n21436_, new_n21437_, new_n21438_, new_n21439_, new_n21440_,
    new_n21441_, new_n21442_, new_n21443_, new_n21444_, new_n21445_,
    new_n21446_, new_n21447_, new_n21448_, new_n21449_, new_n21450_,
    new_n21451_, new_n21452_, new_n21453_, new_n21454_, new_n21455_,
    new_n21456_, new_n21457_, new_n21458_, new_n21459_, new_n21460_,
    new_n21461_, new_n21462_, new_n21463_, new_n21464_, new_n21465_,
    new_n21466_, new_n21467_, new_n21468_, new_n21469_, new_n21470_,
    new_n21471_, new_n21472_, new_n21473_, new_n21474_, new_n21475_,
    new_n21476_, new_n21477_, new_n21478_, new_n21479_, new_n21480_,
    new_n21481_, new_n21482_, new_n21483_, new_n21484_, new_n21485_,
    new_n21486_, new_n21487_, new_n21488_, new_n21489_, new_n21490_,
    new_n21491_, new_n21492_, new_n21493_, new_n21494_, new_n21495_,
    new_n21496_, new_n21497_, new_n21498_, new_n21499_, new_n21500_,
    new_n21501_, new_n21502_, new_n21503_, new_n21504_, new_n21505_,
    new_n21506_, new_n21507_, new_n21508_, new_n21509_, new_n21510_,
    new_n21511_, new_n21512_, new_n21513_, new_n21514_, new_n21515_,
    new_n21516_, new_n21517_, new_n21518_, new_n21519_, new_n21520_,
    new_n21521_, new_n21522_, new_n21523_, new_n21524_, new_n21525_,
    new_n21526_, new_n21527_, new_n21528_, new_n21529_, new_n21530_,
    new_n21531_, new_n21532_, new_n21533_, new_n21534_, new_n21535_,
    new_n21536_, new_n21537_, new_n21539_, new_n21540_, new_n21541_,
    new_n21542_, new_n21543_, new_n21544_, new_n21545_, new_n21546_,
    new_n21547_, new_n21548_, new_n21549_, new_n21550_, new_n21551_,
    new_n21552_, new_n21553_, new_n21554_, new_n21555_, new_n21556_,
    new_n21557_, new_n21558_, new_n21559_, new_n21560_, new_n21561_,
    new_n21562_, new_n21563_, new_n21564_, new_n21565_, new_n21566_,
    new_n21567_, new_n21568_, new_n21569_, new_n21570_, new_n21571_,
    new_n21572_, new_n21573_, new_n21574_, new_n21575_, new_n21576_,
    new_n21577_, new_n21578_, new_n21579_, new_n21580_, new_n21581_,
    new_n21582_, new_n21583_, new_n21584_, new_n21585_, new_n21586_,
    new_n21587_, new_n21588_, new_n21589_, new_n21590_, new_n21591_,
    new_n21592_, new_n21593_, new_n21594_, new_n21595_, new_n21596_,
    new_n21597_, new_n21598_, new_n21599_, new_n21600_, new_n21601_,
    new_n21602_, new_n21603_, new_n21604_, new_n21605_, new_n21606_,
    new_n21607_, new_n21608_, new_n21609_, new_n21610_, new_n21611_,
    new_n21612_, new_n21613_, new_n21614_, new_n21615_, new_n21616_,
    new_n21617_, new_n21618_, new_n21619_, new_n21620_, new_n21621_,
    new_n21622_, new_n21623_, new_n21624_, new_n21625_, new_n21626_,
    new_n21627_, new_n21628_, new_n21629_, new_n21630_, new_n21631_,
    new_n21632_, new_n21633_, new_n21634_, new_n21635_, new_n21636_,
    new_n21637_, new_n21638_, new_n21639_, new_n21640_, new_n21641_,
    new_n21642_, new_n21643_, new_n21644_, new_n21645_, new_n21646_,
    new_n21647_, new_n21648_, new_n21649_, new_n21650_, new_n21651_,
    new_n21652_, new_n21653_, new_n21654_, new_n21655_, new_n21656_,
    new_n21657_, new_n21658_, new_n21659_, new_n21660_, new_n21661_,
    new_n21662_, new_n21663_, new_n21664_, new_n21665_, new_n21666_,
    new_n21667_, new_n21668_, new_n21669_, new_n21670_, new_n21671_,
    new_n21672_, new_n21673_, new_n21674_, new_n21675_, new_n21676_,
    new_n21677_, new_n21678_, new_n21679_, new_n21680_, new_n21681_,
    new_n21682_, new_n21683_, new_n21684_, new_n21685_, new_n21686_,
    new_n21687_, new_n21688_, new_n21689_, new_n21690_, new_n21691_,
    new_n21692_, new_n21693_, new_n21694_, new_n21695_, new_n21696_,
    new_n21697_, new_n21698_, new_n21699_, new_n21700_, new_n21701_,
    new_n21702_, new_n21703_, new_n21704_, new_n21705_, new_n21706_,
    new_n21707_, new_n21708_, new_n21709_, new_n21710_, new_n21711_,
    new_n21712_, new_n21713_, new_n21714_, new_n21715_, new_n21716_,
    new_n21717_, new_n21718_, new_n21719_, new_n21720_, new_n21721_,
    new_n21722_, new_n21723_, new_n21724_, new_n21725_, new_n21726_,
    new_n21727_, new_n21728_, new_n21729_, new_n21730_, new_n21731_,
    new_n21732_, new_n21733_, new_n21734_, new_n21735_, new_n21736_,
    new_n21737_, new_n21738_, new_n21739_, new_n21740_, new_n21741_,
    new_n21742_, new_n21743_, new_n21744_, new_n21745_, new_n21746_,
    new_n21747_, new_n21748_, new_n21749_, new_n21750_, new_n21751_,
    new_n21752_, new_n21753_, new_n21754_, new_n21755_, new_n21756_,
    new_n21757_, new_n21758_, new_n21759_, new_n21760_, new_n21761_,
    new_n21762_, new_n21763_, new_n21764_, new_n21765_, new_n21766_,
    new_n21767_, new_n21768_, new_n21769_, new_n21770_, new_n21771_,
    new_n21772_, new_n21773_, new_n21774_, new_n21775_, new_n21776_,
    new_n21777_, new_n21778_, new_n21779_, new_n21780_, new_n21781_,
    new_n21782_, new_n21783_, new_n21784_, new_n21785_, new_n21786_,
    new_n21787_, new_n21788_, new_n21789_, new_n21790_, new_n21791_,
    new_n21792_, new_n21793_, new_n21794_, new_n21795_, new_n21796_,
    new_n21797_, new_n21798_, new_n21799_, new_n21800_, new_n21801_,
    new_n21802_, new_n21803_, new_n21804_, new_n21805_, new_n21806_,
    new_n21807_, new_n21808_, new_n21809_, new_n21810_, new_n21811_,
    new_n21812_, new_n21813_, new_n21814_, new_n21815_, new_n21816_,
    new_n21817_, new_n21818_, new_n21819_, new_n21820_, new_n21821_,
    new_n21822_, new_n21823_, new_n21824_, new_n21825_, new_n21826_,
    new_n21827_, new_n21828_, new_n21829_, new_n21830_, new_n21831_,
    new_n21832_, new_n21833_, new_n21834_, new_n21835_, new_n21836_,
    new_n21837_, new_n21838_, new_n21839_, new_n21840_, new_n21841_,
    new_n21842_, new_n21843_, new_n21844_, new_n21845_, new_n21846_,
    new_n21847_, new_n21848_, new_n21849_, new_n21850_, new_n21851_,
    new_n21852_, new_n21853_, new_n21854_, new_n21855_, new_n21856_,
    new_n21857_, new_n21858_, new_n21859_, new_n21860_, new_n21861_,
    new_n21862_, new_n21863_, new_n21864_, new_n21865_, new_n21866_,
    new_n21867_, new_n21868_, new_n21869_, new_n21870_, new_n21871_,
    new_n21872_, new_n21873_, new_n21874_, new_n21875_, new_n21876_,
    new_n21877_, new_n21878_, new_n21879_, new_n21880_, new_n21881_,
    new_n21882_, new_n21883_, new_n21884_, new_n21885_, new_n21886_,
    new_n21887_, new_n21888_, new_n21889_, new_n21890_, new_n21891_,
    new_n21892_, new_n21893_, new_n21894_, new_n21895_, new_n21896_,
    new_n21897_, new_n21898_, new_n21899_, new_n21900_, new_n21901_,
    new_n21902_, new_n21903_, new_n21904_, new_n21905_, new_n21906_,
    new_n21907_, new_n21908_, new_n21909_, new_n21910_, new_n21911_,
    new_n21912_, new_n21913_, new_n21914_, new_n21915_, new_n21916_,
    new_n21917_, new_n21918_, new_n21919_, new_n21920_, new_n21921_,
    new_n21922_, new_n21923_, new_n21924_, new_n21925_, new_n21926_,
    new_n21927_, new_n21928_, new_n21929_, new_n21930_, new_n21931_,
    new_n21932_, new_n21933_, new_n21934_, new_n21935_, new_n21936_,
    new_n21937_, new_n21938_, new_n21939_, new_n21940_, new_n21941_,
    new_n21942_, new_n21943_, new_n21944_, new_n21945_, new_n21946_,
    new_n21947_, new_n21948_, new_n21949_, new_n21950_, new_n21951_,
    new_n21952_, new_n21953_, new_n21954_, new_n21955_, new_n21956_,
    new_n21957_, new_n21958_, new_n21959_, new_n21960_, new_n21961_,
    new_n21962_, new_n21963_, new_n21964_, new_n21965_, new_n21966_,
    new_n21967_, new_n21968_, new_n21969_, new_n21970_, new_n21971_,
    new_n21972_, new_n21973_, new_n21974_, new_n21975_, new_n21976_,
    new_n21977_, new_n21978_, new_n21979_, new_n21980_, new_n21981_,
    new_n21982_, new_n21983_, new_n21984_, new_n21985_, new_n21986_,
    new_n21987_, new_n21988_, new_n21989_, new_n21990_, new_n21991_,
    new_n21992_, new_n21993_, new_n21994_, new_n21995_, new_n21996_,
    new_n21997_, new_n21998_, new_n21999_, new_n22000_, new_n22001_,
    new_n22002_, new_n22003_, new_n22004_, new_n22005_, new_n22006_,
    new_n22007_, new_n22008_, new_n22009_, new_n22010_, new_n22011_,
    new_n22012_, new_n22013_, new_n22014_, new_n22015_, new_n22016_,
    new_n22017_, new_n22018_, new_n22019_, new_n22020_, new_n22021_,
    new_n22022_, new_n22023_, new_n22024_, new_n22025_, new_n22026_,
    new_n22027_, new_n22028_, new_n22029_, new_n22030_, new_n22031_,
    new_n22032_, new_n22033_, new_n22034_, new_n22035_, new_n22036_,
    new_n22037_, new_n22038_, new_n22039_, new_n22040_, new_n22041_,
    new_n22042_, new_n22043_, new_n22044_, new_n22045_, new_n22046_,
    new_n22047_, new_n22048_, new_n22049_, new_n22050_, new_n22051_,
    new_n22052_, new_n22053_, new_n22054_, new_n22055_, new_n22056_,
    new_n22057_, new_n22058_, new_n22059_, new_n22060_, new_n22061_,
    new_n22062_, new_n22063_, new_n22064_, new_n22065_, new_n22066_,
    new_n22067_, new_n22068_, new_n22069_, new_n22070_, new_n22071_,
    new_n22072_, new_n22073_, new_n22074_, new_n22075_, new_n22076_,
    new_n22077_, new_n22078_, new_n22079_, new_n22080_, new_n22081_,
    new_n22082_, new_n22083_, new_n22084_, new_n22085_, new_n22086_,
    new_n22087_, new_n22088_, new_n22089_, new_n22090_, new_n22091_,
    new_n22092_, new_n22093_, new_n22094_, new_n22095_, new_n22096_,
    new_n22097_, new_n22098_, new_n22099_, new_n22100_, new_n22101_,
    new_n22102_, new_n22103_, new_n22104_, new_n22105_, new_n22106_,
    new_n22107_, new_n22108_, new_n22109_, new_n22110_, new_n22111_,
    new_n22112_, new_n22113_, new_n22114_, new_n22115_, new_n22116_,
    new_n22117_, new_n22118_, new_n22119_, new_n22120_, new_n22121_,
    new_n22122_, new_n22123_, new_n22124_, new_n22125_, new_n22126_,
    new_n22127_, new_n22128_, new_n22129_, new_n22130_, new_n22131_,
    new_n22132_, new_n22133_, new_n22134_, new_n22135_, new_n22136_,
    new_n22137_, new_n22138_, new_n22139_, new_n22140_, new_n22141_,
    new_n22142_, new_n22143_, new_n22144_, new_n22145_, new_n22146_,
    new_n22147_, new_n22148_, new_n22149_, new_n22150_, new_n22151_,
    new_n22152_, new_n22153_, new_n22154_, new_n22155_, new_n22156_,
    new_n22157_, new_n22158_, new_n22159_, new_n22160_, new_n22161_,
    new_n22162_, new_n22163_, new_n22164_, new_n22165_, new_n22166_,
    new_n22167_, new_n22168_, new_n22169_, new_n22170_, new_n22171_,
    new_n22172_, new_n22173_, new_n22174_, new_n22175_, new_n22176_,
    new_n22177_, new_n22178_, new_n22179_, new_n22180_, new_n22181_,
    new_n22182_, new_n22183_, new_n22184_, new_n22185_, new_n22186_,
    new_n22187_, new_n22188_, new_n22189_, new_n22190_, new_n22191_,
    new_n22192_, new_n22193_, new_n22194_, new_n22195_, new_n22196_,
    new_n22197_, new_n22198_, new_n22199_, new_n22200_, new_n22201_,
    new_n22202_, new_n22203_, new_n22204_, new_n22205_, new_n22206_,
    new_n22207_, new_n22208_, new_n22209_, new_n22210_, new_n22211_,
    new_n22212_, new_n22213_, new_n22214_, new_n22215_, new_n22216_,
    new_n22217_, new_n22218_, new_n22219_, new_n22220_, new_n22221_,
    new_n22222_, new_n22223_, new_n22224_, new_n22225_, new_n22226_,
    new_n22227_, new_n22228_, new_n22229_, new_n22230_, new_n22231_,
    new_n22232_, new_n22233_, new_n22234_, new_n22235_, new_n22236_,
    new_n22237_, new_n22238_, new_n22239_, new_n22240_, new_n22241_,
    new_n22242_, new_n22243_, new_n22244_, new_n22245_, new_n22246_,
    new_n22247_, new_n22248_, new_n22249_, new_n22250_, new_n22251_,
    new_n22252_, new_n22253_, new_n22254_, new_n22255_, new_n22256_,
    new_n22257_, new_n22258_, new_n22259_, new_n22260_, new_n22261_,
    new_n22262_, new_n22263_, new_n22264_, new_n22265_, new_n22266_,
    new_n22267_, new_n22268_, new_n22269_, new_n22270_, new_n22271_,
    new_n22272_, new_n22273_, new_n22274_, new_n22275_, new_n22276_,
    new_n22277_, new_n22278_, new_n22279_, new_n22280_, new_n22281_,
    new_n22282_, new_n22283_, new_n22284_, new_n22285_, new_n22286_,
    new_n22287_, new_n22288_, new_n22289_, new_n22290_, new_n22291_,
    new_n22292_, new_n22293_, new_n22294_, new_n22295_, new_n22296_,
    new_n22297_, new_n22298_, new_n22299_, new_n22300_, new_n22301_,
    new_n22302_, new_n22303_, new_n22304_, new_n22305_, new_n22306_,
    new_n22307_, new_n22308_, new_n22309_, new_n22310_, new_n22311_,
    new_n22313_, new_n22314_, new_n22315_, new_n22316_, new_n22317_,
    new_n22318_, new_n22319_, new_n22320_, new_n22321_, new_n22322_,
    new_n22323_, new_n22324_, new_n22325_, new_n22326_, new_n22327_,
    new_n22328_, new_n22329_, new_n22330_, new_n22331_, new_n22332_,
    new_n22333_, new_n22334_, new_n22335_, new_n22336_, new_n22337_,
    new_n22338_, new_n22339_, new_n22340_, new_n22341_, new_n22342_,
    new_n22343_, new_n22344_, new_n22345_, new_n22346_, new_n22347_,
    new_n22348_, new_n22349_, new_n22350_, new_n22351_, new_n22352_,
    new_n22353_, new_n22354_, new_n22355_, new_n22356_, new_n22357_,
    new_n22358_, new_n22359_, new_n22360_, new_n22361_, new_n22362_,
    new_n22363_, new_n22364_, new_n22365_, new_n22366_, new_n22367_,
    new_n22368_, new_n22369_, new_n22370_, new_n22371_, new_n22372_,
    new_n22373_, new_n22374_, new_n22375_, new_n22376_, new_n22377_,
    new_n22378_, new_n22379_, new_n22380_, new_n22381_, new_n22382_,
    new_n22383_, new_n22384_, new_n22385_, new_n22386_, new_n22387_,
    new_n22388_, new_n22389_, new_n22390_, new_n22391_, new_n22392_,
    new_n22393_, new_n22394_, new_n22395_, new_n22396_, new_n22397_,
    new_n22398_, new_n22399_, new_n22400_, new_n22401_, new_n22402_,
    new_n22403_, new_n22404_, new_n22405_, new_n22406_, new_n22407_,
    new_n22408_, new_n22409_, new_n22410_, new_n22411_, new_n22412_,
    new_n22413_, new_n22414_, new_n22415_, new_n22416_, new_n22417_,
    new_n22418_, new_n22419_, new_n22420_, new_n22421_, new_n22422_,
    new_n22423_, new_n22424_, new_n22425_, new_n22426_, new_n22427_,
    new_n22428_, new_n22429_, new_n22430_, new_n22431_, new_n22432_,
    new_n22433_, new_n22434_, new_n22435_, new_n22436_, new_n22437_,
    new_n22438_, new_n22439_, new_n22440_, new_n22441_, new_n22442_,
    new_n22443_, new_n22444_, new_n22445_, new_n22446_, new_n22447_,
    new_n22448_, new_n22449_, new_n22450_, new_n22451_, new_n22452_,
    new_n22453_, new_n22454_, new_n22455_, new_n22456_, new_n22457_,
    new_n22458_, new_n22459_, new_n22460_, new_n22461_, new_n22462_,
    new_n22463_, new_n22464_, new_n22465_, new_n22466_, new_n22467_,
    new_n22468_, new_n22469_, new_n22470_, new_n22471_, new_n22472_,
    new_n22473_, new_n22474_, new_n22475_, new_n22476_, new_n22477_,
    new_n22478_, new_n22479_, new_n22480_, new_n22481_, new_n22482_,
    new_n22483_, new_n22484_, new_n22485_, new_n22486_, new_n22487_,
    new_n22488_, new_n22489_, new_n22490_, new_n22491_, new_n22492_,
    new_n22493_, new_n22494_, new_n22495_, new_n22496_, new_n22497_,
    new_n22498_, new_n22499_, new_n22500_, new_n22501_, new_n22502_,
    new_n22503_, new_n22504_, new_n22505_, new_n22506_, new_n22507_,
    new_n22508_, new_n22509_, new_n22510_, new_n22511_, new_n22512_,
    new_n22513_, new_n22514_, new_n22515_, new_n22516_, new_n22517_,
    new_n22518_, new_n22519_, new_n22520_, new_n22521_, new_n22522_,
    new_n22523_, new_n22524_, new_n22525_, new_n22526_, new_n22527_,
    new_n22528_, new_n22529_, new_n22530_, new_n22531_, new_n22532_,
    new_n22533_, new_n22534_, new_n22535_, new_n22536_, new_n22537_,
    new_n22538_, new_n22539_, new_n22540_, new_n22541_, new_n22542_,
    new_n22543_, new_n22544_, new_n22545_, new_n22546_, new_n22547_,
    new_n22548_, new_n22549_, new_n22550_, new_n22551_, new_n22552_,
    new_n22553_, new_n22554_, new_n22555_, new_n22556_, new_n22557_,
    new_n22558_, new_n22559_, new_n22560_, new_n22561_, new_n22562_,
    new_n22563_, new_n22564_, new_n22565_, new_n22566_, new_n22567_,
    new_n22568_, new_n22569_, new_n22570_, new_n22571_, new_n22572_,
    new_n22573_, new_n22574_, new_n22575_, new_n22576_, new_n22577_,
    new_n22578_, new_n22579_, new_n22580_, new_n22581_, new_n22582_,
    new_n22583_, new_n22584_, new_n22585_, new_n22586_, new_n22587_,
    new_n22588_, new_n22589_, new_n22590_, new_n22591_, new_n22592_,
    new_n22593_, new_n22594_, new_n22595_, new_n22596_, new_n22597_,
    new_n22598_, new_n22599_, new_n22600_, new_n22601_, new_n22602_,
    new_n22603_, new_n22604_, new_n22605_, new_n22606_, new_n22607_,
    new_n22608_, new_n22609_, new_n22610_, new_n22611_, new_n22612_,
    new_n22613_, new_n22614_, new_n22615_, new_n22616_, new_n22617_,
    new_n22618_, new_n22619_, new_n22620_, new_n22621_, new_n22622_,
    new_n22623_, new_n22624_, new_n22625_, new_n22626_, new_n22627_,
    new_n22628_, new_n22629_, new_n22630_, new_n22631_, new_n22632_,
    new_n22633_, new_n22634_, new_n22635_, new_n22636_, new_n22637_,
    new_n22638_, new_n22639_, new_n22640_, new_n22641_, new_n22642_,
    new_n22643_, new_n22644_, new_n22645_, new_n22646_, new_n22647_,
    new_n22648_, new_n22649_, new_n22650_, new_n22651_, new_n22652_,
    new_n22653_, new_n22654_, new_n22655_, new_n22656_, new_n22657_,
    new_n22658_, new_n22659_, new_n22660_, new_n22661_, new_n22662_,
    new_n22663_, new_n22664_, new_n22665_, new_n22666_, new_n22667_,
    new_n22668_, new_n22669_, new_n22670_, new_n22671_, new_n22672_,
    new_n22673_, new_n22674_, new_n22675_, new_n22676_, new_n22677_,
    new_n22678_, new_n22679_, new_n22680_, new_n22681_, new_n22682_,
    new_n22683_, new_n22684_, new_n22685_, new_n22686_, new_n22687_,
    new_n22688_, new_n22689_, new_n22690_, new_n22691_, new_n22692_,
    new_n22693_, new_n22694_, new_n22695_, new_n22696_, new_n22697_,
    new_n22698_, new_n22699_, new_n22700_, new_n22701_, new_n22702_,
    new_n22703_, new_n22704_, new_n22705_, new_n22706_, new_n22707_,
    new_n22708_, new_n22709_, new_n22710_, new_n22711_, new_n22712_,
    new_n22713_, new_n22714_, new_n22715_, new_n22716_, new_n22717_,
    new_n22718_, new_n22719_, new_n22720_, new_n22721_, new_n22722_,
    new_n22723_, new_n22724_, new_n22725_, new_n22726_, new_n22727_,
    new_n22728_, new_n22729_, new_n22730_, new_n22731_, new_n22732_,
    new_n22733_, new_n22734_, new_n22735_, new_n22736_, new_n22737_,
    new_n22738_, new_n22739_, new_n22740_, new_n22741_, new_n22742_,
    new_n22743_, new_n22744_, new_n22745_, new_n22746_, new_n22747_,
    new_n22748_, new_n22749_, new_n22750_, new_n22751_, new_n22752_,
    new_n22753_, new_n22754_, new_n22755_, new_n22756_, new_n22757_,
    new_n22758_, new_n22759_, new_n22760_, new_n22761_, new_n22762_,
    new_n22763_, new_n22764_, new_n22765_, new_n22766_, new_n22767_,
    new_n22768_, new_n22769_, new_n22770_, new_n22771_, new_n22772_,
    new_n22773_, new_n22774_, new_n22775_, new_n22776_, new_n22777_,
    new_n22778_, new_n22779_, new_n22780_, new_n22781_, new_n22782_,
    new_n22783_, new_n22784_, new_n22785_, new_n22786_, new_n22787_,
    new_n22788_, new_n22789_, new_n22790_, new_n22791_, new_n22792_,
    new_n22793_, new_n22794_, new_n22795_, new_n22796_, new_n22797_,
    new_n22798_, new_n22799_, new_n22800_, new_n22801_, new_n22802_,
    new_n22803_, new_n22804_, new_n22805_, new_n22806_, new_n22807_,
    new_n22808_, new_n22809_, new_n22810_, new_n22811_, new_n22812_,
    new_n22813_, new_n22814_, new_n22815_, new_n22816_, new_n22817_,
    new_n22818_, new_n22819_, new_n22820_, new_n22821_, new_n22822_,
    new_n22823_, new_n22824_, new_n22825_, new_n22826_, new_n22827_,
    new_n22828_, new_n22829_, new_n22830_, new_n22831_, new_n22832_,
    new_n22833_, new_n22834_, new_n22835_, new_n22836_, new_n22837_,
    new_n22838_, new_n22839_, new_n22840_, new_n22841_, new_n22842_,
    new_n22843_, new_n22844_, new_n22845_, new_n22846_, new_n22847_,
    new_n22848_, new_n22849_, new_n22850_, new_n22851_, new_n22852_,
    new_n22853_, new_n22854_, new_n22855_, new_n22856_, new_n22857_,
    new_n22858_, new_n22859_, new_n22860_, new_n22861_, new_n22862_,
    new_n22863_, new_n22864_, new_n22865_, new_n22866_, new_n22867_,
    new_n22868_, new_n22869_, new_n22870_, new_n22871_, new_n22872_,
    new_n22873_, new_n22874_, new_n22875_, new_n22876_, new_n22877_,
    new_n22878_, new_n22879_, new_n22880_, new_n22881_, new_n22882_,
    new_n22883_, new_n22884_, new_n22885_, new_n22886_, new_n22887_,
    new_n22888_, new_n22889_, new_n22890_, new_n22891_, new_n22892_,
    new_n22893_, new_n22894_, new_n22895_, new_n22896_, new_n22897_,
    new_n22898_, new_n22899_, new_n22900_, new_n22901_, new_n22902_,
    new_n22903_, new_n22904_, new_n22905_, new_n22906_, new_n22907_,
    new_n22908_, new_n22909_, new_n22910_, new_n22911_, new_n22912_,
    new_n22913_, new_n22914_, new_n22915_, new_n22916_, new_n22917_,
    new_n22918_, new_n22919_, new_n22920_, new_n22921_, new_n22922_,
    new_n22923_, new_n22924_, new_n22925_, new_n22926_, new_n22927_,
    new_n22928_, new_n22929_, new_n22930_, new_n22931_, new_n22932_,
    new_n22933_, new_n22934_, new_n22935_, new_n22936_, new_n22937_,
    new_n22938_, new_n22939_, new_n22940_, new_n22941_, new_n22942_,
    new_n22943_, new_n22944_, new_n22945_, new_n22946_, new_n22947_,
    new_n22948_, new_n22949_, new_n22950_, new_n22951_, new_n22952_,
    new_n22953_, new_n22954_, new_n22955_, new_n22956_, new_n22957_,
    new_n22958_, new_n22959_, new_n22960_, new_n22961_, new_n22962_,
    new_n22963_, new_n22964_, new_n22965_, new_n22966_, new_n22967_,
    new_n22968_, new_n22969_, new_n22970_, new_n22971_, new_n22972_,
    new_n22973_, new_n22974_, new_n22975_, new_n22976_, new_n22977_,
    new_n22978_, new_n22979_, new_n22980_, new_n22981_, new_n22982_,
    new_n22983_, new_n22984_, new_n22985_, new_n22986_, new_n22987_,
    new_n22988_, new_n22989_, new_n22990_, new_n22991_, new_n22992_,
    new_n22993_, new_n22994_, new_n22995_, new_n22996_, new_n22997_,
    new_n22998_, new_n22999_, new_n23000_, new_n23001_, new_n23002_,
    new_n23003_, new_n23004_, new_n23005_, new_n23006_, new_n23007_,
    new_n23008_, new_n23009_, new_n23010_, new_n23011_, new_n23012_,
    new_n23013_, new_n23014_, new_n23015_, new_n23016_, new_n23017_,
    new_n23018_, new_n23019_, new_n23020_, new_n23021_, new_n23022_,
    new_n23023_, new_n23024_, new_n23025_, new_n23026_, new_n23027_,
    new_n23028_, new_n23029_, new_n23030_, new_n23031_, new_n23032_,
    new_n23033_, new_n23034_, new_n23035_, new_n23036_, new_n23037_,
    new_n23038_, new_n23039_, new_n23040_, new_n23041_, new_n23042_,
    new_n23043_, new_n23044_, new_n23045_, new_n23046_, new_n23047_,
    new_n23048_, new_n23049_, new_n23050_, new_n23051_, new_n23052_,
    new_n23053_, new_n23054_, new_n23055_, new_n23056_, new_n23057_,
    new_n23058_, new_n23059_, new_n23060_, new_n23061_, new_n23062_,
    new_n23063_, new_n23064_, new_n23065_, new_n23066_, new_n23067_,
    new_n23068_, new_n23069_, new_n23070_, new_n23071_, new_n23072_,
    new_n23073_, new_n23074_, new_n23075_, new_n23076_, new_n23077_,
    new_n23078_, new_n23079_, new_n23080_, new_n23081_, new_n23082_,
    new_n23083_, new_n23084_, new_n23085_, new_n23086_, new_n23087_,
    new_n23088_, new_n23089_, new_n23090_, new_n23091_, new_n23092_,
    new_n23093_, new_n23094_, new_n23095_, new_n23096_, new_n23098_,
    new_n23099_, new_n23100_, new_n23101_, new_n23102_, new_n23103_,
    new_n23104_, new_n23105_, new_n23106_, new_n23107_, new_n23108_,
    new_n23109_, new_n23110_, new_n23111_, new_n23112_, new_n23113_,
    new_n23114_, new_n23115_, new_n23116_, new_n23117_, new_n23118_,
    new_n23119_, new_n23120_, new_n23121_, new_n23122_, new_n23123_,
    new_n23124_, new_n23125_, new_n23126_, new_n23127_, new_n23128_,
    new_n23129_, new_n23130_, new_n23131_, new_n23132_, new_n23133_,
    new_n23134_, new_n23135_, new_n23136_, new_n23137_, new_n23138_,
    new_n23139_, new_n23140_, new_n23141_, new_n23142_, new_n23143_,
    new_n23144_, new_n23145_, new_n23146_, new_n23147_, new_n23148_,
    new_n23149_, new_n23150_, new_n23151_, new_n23152_, new_n23153_,
    new_n23154_, new_n23155_, new_n23156_, new_n23157_, new_n23158_,
    new_n23159_, new_n23160_, new_n23161_, new_n23162_, new_n23163_,
    new_n23164_, new_n23165_, new_n23166_, new_n23167_, new_n23168_,
    new_n23169_, new_n23170_, new_n23171_, new_n23172_, new_n23173_,
    new_n23174_, new_n23175_, new_n23176_, new_n23177_, new_n23178_,
    new_n23179_, new_n23180_, new_n23181_, new_n23182_, new_n23183_,
    new_n23184_, new_n23185_, new_n23186_, new_n23187_, new_n23188_,
    new_n23189_, new_n23190_, new_n23191_, new_n23192_, new_n23193_,
    new_n23194_, new_n23195_, new_n23196_, new_n23197_, new_n23198_,
    new_n23199_, new_n23200_, new_n23201_, new_n23202_, new_n23203_,
    new_n23204_, new_n23205_, new_n23206_, new_n23207_, new_n23208_,
    new_n23209_, new_n23210_, new_n23211_, new_n23212_, new_n23213_,
    new_n23214_, new_n23215_, new_n23216_, new_n23217_, new_n23218_,
    new_n23219_, new_n23220_, new_n23221_, new_n23222_, new_n23223_,
    new_n23224_, new_n23225_, new_n23226_, new_n23227_, new_n23228_,
    new_n23229_, new_n23230_, new_n23231_, new_n23232_, new_n23233_,
    new_n23234_, new_n23235_, new_n23236_, new_n23237_, new_n23238_,
    new_n23239_, new_n23240_, new_n23241_, new_n23242_, new_n23243_,
    new_n23244_, new_n23245_, new_n23246_, new_n23247_, new_n23248_,
    new_n23249_, new_n23250_, new_n23251_, new_n23252_, new_n23253_,
    new_n23254_, new_n23255_, new_n23256_, new_n23257_, new_n23258_,
    new_n23259_, new_n23260_, new_n23261_, new_n23262_, new_n23263_,
    new_n23264_, new_n23265_, new_n23266_, new_n23267_, new_n23268_,
    new_n23269_, new_n23270_, new_n23271_, new_n23272_, new_n23273_,
    new_n23274_, new_n23275_, new_n23276_, new_n23277_, new_n23278_,
    new_n23279_, new_n23280_, new_n23281_, new_n23282_, new_n23283_,
    new_n23284_, new_n23285_, new_n23286_, new_n23287_, new_n23288_,
    new_n23289_, new_n23290_, new_n23291_, new_n23292_, new_n23293_,
    new_n23294_, new_n23295_, new_n23296_, new_n23297_, new_n23298_,
    new_n23299_, new_n23300_, new_n23301_, new_n23302_, new_n23303_,
    new_n23304_, new_n23305_, new_n23306_, new_n23307_, new_n23308_,
    new_n23309_, new_n23310_, new_n23311_, new_n23312_, new_n23313_,
    new_n23314_, new_n23315_, new_n23316_, new_n23317_, new_n23318_,
    new_n23319_, new_n23320_, new_n23321_, new_n23322_, new_n23323_,
    new_n23324_, new_n23325_, new_n23326_, new_n23327_, new_n23328_,
    new_n23329_, new_n23330_, new_n23331_, new_n23332_, new_n23333_,
    new_n23334_, new_n23335_, new_n23336_, new_n23337_, new_n23338_,
    new_n23339_, new_n23340_, new_n23341_, new_n23342_, new_n23343_,
    new_n23344_, new_n23345_, new_n23346_, new_n23347_, new_n23348_,
    new_n23349_, new_n23350_, new_n23351_, new_n23352_, new_n23353_,
    new_n23354_, new_n23355_, new_n23356_, new_n23357_, new_n23358_,
    new_n23359_, new_n23360_, new_n23361_, new_n23362_, new_n23363_,
    new_n23364_, new_n23365_, new_n23366_, new_n23367_, new_n23368_,
    new_n23369_, new_n23370_, new_n23371_, new_n23372_, new_n23373_,
    new_n23374_, new_n23375_, new_n23376_, new_n23377_, new_n23378_,
    new_n23379_, new_n23380_, new_n23381_, new_n23382_, new_n23383_,
    new_n23384_, new_n23385_, new_n23386_, new_n23387_, new_n23388_,
    new_n23389_, new_n23390_, new_n23391_, new_n23392_, new_n23393_,
    new_n23394_, new_n23395_, new_n23396_, new_n23397_, new_n23398_,
    new_n23399_, new_n23400_, new_n23401_, new_n23402_, new_n23403_,
    new_n23404_, new_n23405_, new_n23406_, new_n23407_, new_n23408_,
    new_n23409_, new_n23410_, new_n23411_, new_n23412_, new_n23413_,
    new_n23414_, new_n23415_, new_n23416_, new_n23417_, new_n23418_,
    new_n23419_, new_n23420_, new_n23421_, new_n23422_, new_n23423_,
    new_n23424_, new_n23425_, new_n23426_, new_n23427_, new_n23428_,
    new_n23429_, new_n23430_, new_n23431_, new_n23432_, new_n23433_,
    new_n23434_, new_n23435_, new_n23436_, new_n23437_, new_n23438_,
    new_n23439_, new_n23440_, new_n23441_, new_n23442_, new_n23443_,
    new_n23444_, new_n23445_, new_n23446_, new_n23447_, new_n23448_,
    new_n23449_, new_n23450_, new_n23451_, new_n23452_, new_n23453_,
    new_n23454_, new_n23455_, new_n23456_, new_n23457_, new_n23458_,
    new_n23459_, new_n23460_, new_n23461_, new_n23462_, new_n23463_,
    new_n23464_, new_n23465_, new_n23466_, new_n23467_, new_n23468_,
    new_n23469_, new_n23470_, new_n23471_, new_n23472_, new_n23473_,
    new_n23474_, new_n23475_, new_n23476_, new_n23477_, new_n23478_,
    new_n23479_, new_n23480_, new_n23481_, new_n23482_, new_n23483_,
    new_n23484_, new_n23485_, new_n23486_, new_n23487_, new_n23488_,
    new_n23489_, new_n23490_, new_n23491_, new_n23492_, new_n23493_,
    new_n23494_, new_n23495_, new_n23496_, new_n23497_, new_n23498_,
    new_n23499_, new_n23500_, new_n23501_, new_n23502_, new_n23503_,
    new_n23504_, new_n23505_, new_n23506_, new_n23507_, new_n23508_,
    new_n23509_, new_n23510_, new_n23511_, new_n23512_, new_n23513_,
    new_n23514_, new_n23515_, new_n23516_, new_n23517_, new_n23518_,
    new_n23519_, new_n23520_, new_n23521_, new_n23522_, new_n23523_,
    new_n23524_, new_n23525_, new_n23526_, new_n23527_, new_n23528_,
    new_n23529_, new_n23530_, new_n23531_, new_n23532_, new_n23533_,
    new_n23534_, new_n23535_, new_n23536_, new_n23537_, new_n23538_,
    new_n23539_, new_n23540_, new_n23541_, new_n23542_, new_n23543_,
    new_n23544_, new_n23545_, new_n23546_, new_n23547_, new_n23548_,
    new_n23549_, new_n23550_, new_n23551_, new_n23552_, new_n23553_,
    new_n23554_, new_n23555_, new_n23556_, new_n23557_, new_n23558_,
    new_n23559_, new_n23560_, new_n23561_, new_n23562_, new_n23563_,
    new_n23564_, new_n23565_, new_n23566_, new_n23567_, new_n23568_,
    new_n23569_, new_n23570_, new_n23571_, new_n23572_, new_n23573_,
    new_n23574_, new_n23575_, new_n23576_, new_n23577_, new_n23578_,
    new_n23579_, new_n23580_, new_n23581_, new_n23582_, new_n23583_,
    new_n23584_, new_n23585_, new_n23586_, new_n23587_, new_n23588_,
    new_n23589_, new_n23590_, new_n23591_, new_n23592_, new_n23593_,
    new_n23594_, new_n23595_, new_n23596_, new_n23597_, new_n23598_,
    new_n23599_, new_n23600_, new_n23601_, new_n23602_, new_n23603_,
    new_n23604_, new_n23605_, new_n23606_, new_n23607_, new_n23608_,
    new_n23609_, new_n23610_, new_n23611_, new_n23612_, new_n23613_,
    new_n23614_, new_n23615_, new_n23616_, new_n23617_, new_n23618_,
    new_n23619_, new_n23620_, new_n23621_, new_n23622_, new_n23623_,
    new_n23624_, new_n23625_, new_n23626_, new_n23627_, new_n23628_,
    new_n23629_, new_n23630_, new_n23631_, new_n23632_, new_n23633_,
    new_n23634_, new_n23635_, new_n23636_, new_n23637_, new_n23638_,
    new_n23639_, new_n23640_, new_n23641_, new_n23642_, new_n23643_,
    new_n23644_, new_n23645_, new_n23646_, new_n23647_, new_n23648_,
    new_n23649_, new_n23650_, new_n23651_, new_n23652_, new_n23653_,
    new_n23654_, new_n23655_, new_n23656_, new_n23657_, new_n23658_,
    new_n23659_, new_n23660_, new_n23661_, new_n23662_, new_n23663_,
    new_n23664_, new_n23665_, new_n23666_, new_n23667_, new_n23668_,
    new_n23669_, new_n23670_, new_n23671_, new_n23672_, new_n23673_,
    new_n23674_, new_n23675_, new_n23676_, new_n23677_, new_n23678_,
    new_n23679_, new_n23680_, new_n23681_, new_n23682_, new_n23683_,
    new_n23684_, new_n23685_, new_n23686_, new_n23687_, new_n23688_,
    new_n23689_, new_n23690_, new_n23691_, new_n23692_, new_n23693_,
    new_n23694_, new_n23695_, new_n23696_, new_n23697_, new_n23698_,
    new_n23699_, new_n23700_, new_n23701_, new_n23702_, new_n23703_,
    new_n23704_, new_n23705_, new_n23706_, new_n23707_, new_n23708_,
    new_n23709_, new_n23710_, new_n23711_, new_n23712_, new_n23713_,
    new_n23714_, new_n23715_, new_n23716_, new_n23717_, new_n23718_,
    new_n23719_, new_n23720_, new_n23721_, new_n23722_, new_n23723_,
    new_n23724_, new_n23725_, new_n23726_, new_n23727_, new_n23728_,
    new_n23729_, new_n23730_, new_n23731_, new_n23732_, new_n23733_,
    new_n23734_, new_n23735_, new_n23736_, new_n23737_, new_n23738_,
    new_n23739_, new_n23740_, new_n23741_, new_n23742_, new_n23743_,
    new_n23744_, new_n23745_, new_n23746_, new_n23747_, new_n23748_,
    new_n23749_, new_n23750_, new_n23751_, new_n23752_, new_n23753_,
    new_n23754_, new_n23755_, new_n23756_, new_n23757_, new_n23758_,
    new_n23759_, new_n23760_, new_n23761_, new_n23762_, new_n23763_,
    new_n23764_, new_n23765_, new_n23766_, new_n23767_, new_n23768_,
    new_n23769_, new_n23770_, new_n23771_, new_n23772_, new_n23773_,
    new_n23774_, new_n23775_, new_n23776_, new_n23777_, new_n23778_,
    new_n23779_, new_n23780_, new_n23781_, new_n23782_, new_n23783_,
    new_n23784_, new_n23785_, new_n23786_, new_n23787_, new_n23788_,
    new_n23789_, new_n23790_, new_n23791_, new_n23792_, new_n23793_,
    new_n23794_, new_n23795_, new_n23796_, new_n23797_, new_n23798_,
    new_n23799_, new_n23800_, new_n23801_, new_n23802_, new_n23803_,
    new_n23804_, new_n23805_, new_n23806_, new_n23807_, new_n23808_,
    new_n23809_, new_n23810_, new_n23811_, new_n23812_, new_n23813_,
    new_n23814_, new_n23815_, new_n23816_, new_n23817_, new_n23818_,
    new_n23819_, new_n23820_, new_n23821_, new_n23822_, new_n23823_,
    new_n23824_, new_n23825_, new_n23826_, new_n23827_, new_n23828_,
    new_n23829_, new_n23830_, new_n23831_, new_n23832_, new_n23833_,
    new_n23834_, new_n23835_, new_n23836_, new_n23837_, new_n23838_,
    new_n23839_, new_n23840_, new_n23841_, new_n23842_, new_n23843_,
    new_n23844_, new_n23845_, new_n23846_, new_n23847_, new_n23848_,
    new_n23849_, new_n23850_, new_n23851_, new_n23852_, new_n23853_,
    new_n23854_, new_n23855_, new_n23856_, new_n23857_, new_n23858_,
    new_n23859_, new_n23860_, new_n23861_, new_n23862_, new_n23863_,
    new_n23864_, new_n23865_, new_n23866_, new_n23867_, new_n23868_,
    new_n23869_, new_n23870_, new_n23871_, new_n23872_, new_n23873_,
    new_n23874_, new_n23875_, new_n23876_, new_n23877_, new_n23878_,
    new_n23879_, new_n23880_, new_n23881_, new_n23882_, new_n23883_,
    new_n23884_, new_n23885_, new_n23886_, new_n23887_, new_n23888_,
    new_n23889_, new_n23890_, new_n23891_, new_n23892_, new_n23893_,
    new_n23894_, new_n23895_, new_n23897_, new_n23898_, new_n23899_,
    new_n23900_, new_n23901_, new_n23902_, new_n23903_, new_n23904_,
    new_n23905_, new_n23906_, new_n23907_, new_n23908_, new_n23909_,
    new_n23910_, new_n23911_, new_n23912_, new_n23913_, new_n23914_,
    new_n23915_, new_n23916_, new_n23917_, new_n23918_, new_n23919_,
    new_n23920_, new_n23921_, new_n23922_, new_n23923_, new_n23924_,
    new_n23925_, new_n23926_, new_n23927_, new_n23928_, new_n23929_,
    new_n23930_, new_n23931_, new_n23932_, new_n23933_, new_n23934_,
    new_n23935_, new_n23936_, new_n23937_, new_n23938_, new_n23939_,
    new_n23940_, new_n23941_, new_n23942_, new_n23943_, new_n23944_,
    new_n23945_, new_n23946_, new_n23947_, new_n23948_, new_n23949_,
    new_n23950_, new_n23951_, new_n23952_, new_n23953_, new_n23954_,
    new_n23955_, new_n23956_, new_n23957_, new_n23958_, new_n23959_,
    new_n23960_, new_n23961_, new_n23962_, new_n23963_, new_n23964_,
    new_n23965_, new_n23966_, new_n23967_, new_n23968_, new_n23969_,
    new_n23970_, new_n23971_, new_n23972_, new_n23973_, new_n23974_,
    new_n23975_, new_n23976_, new_n23977_, new_n23978_, new_n23979_,
    new_n23980_, new_n23981_, new_n23982_, new_n23983_, new_n23984_,
    new_n23985_, new_n23986_, new_n23987_, new_n23988_, new_n23989_,
    new_n23990_, new_n23991_, new_n23992_, new_n23993_, new_n23994_,
    new_n23995_, new_n23996_, new_n23997_, new_n23998_, new_n23999_,
    new_n24000_, new_n24001_, new_n24002_, new_n24003_, new_n24004_,
    new_n24005_, new_n24006_, new_n24007_, new_n24008_, new_n24009_,
    new_n24010_, new_n24011_, new_n24012_, new_n24013_, new_n24014_,
    new_n24015_, new_n24016_, new_n24017_, new_n24018_, new_n24019_,
    new_n24020_, new_n24021_, new_n24022_, new_n24023_, new_n24024_,
    new_n24025_, new_n24026_, new_n24027_, new_n24028_, new_n24029_,
    new_n24030_, new_n24031_, new_n24032_, new_n24033_, new_n24034_,
    new_n24035_, new_n24036_, new_n24037_, new_n24038_, new_n24039_,
    new_n24040_, new_n24041_, new_n24042_, new_n24043_, new_n24044_,
    new_n24045_, new_n24046_, new_n24047_, new_n24048_, new_n24049_,
    new_n24050_, new_n24051_, new_n24052_, new_n24053_, new_n24054_,
    new_n24055_, new_n24056_, new_n24057_, new_n24058_, new_n24059_,
    new_n24060_, new_n24061_, new_n24062_, new_n24063_, new_n24064_,
    new_n24065_, new_n24066_, new_n24067_, new_n24068_, new_n24069_,
    new_n24070_, new_n24071_, new_n24072_, new_n24073_, new_n24074_,
    new_n24075_, new_n24076_, new_n24077_, new_n24078_, new_n24079_,
    new_n24080_, new_n24081_, new_n24082_, new_n24083_, new_n24084_,
    new_n24085_, new_n24086_, new_n24087_, new_n24088_, new_n24089_,
    new_n24090_, new_n24091_, new_n24092_, new_n24093_, new_n24094_,
    new_n24095_, new_n24096_, new_n24097_, new_n24098_, new_n24099_,
    new_n24100_, new_n24101_, new_n24102_, new_n24103_, new_n24104_,
    new_n24105_, new_n24106_, new_n24107_, new_n24108_, new_n24109_,
    new_n24110_, new_n24111_, new_n24112_, new_n24113_, new_n24114_,
    new_n24115_, new_n24116_, new_n24117_, new_n24118_, new_n24119_,
    new_n24120_, new_n24121_, new_n24122_, new_n24123_, new_n24124_,
    new_n24125_, new_n24126_, new_n24127_, new_n24128_, new_n24129_,
    new_n24130_, new_n24131_, new_n24132_, new_n24133_, new_n24134_,
    new_n24135_, new_n24136_, new_n24137_, new_n24138_, new_n24139_,
    new_n24140_, new_n24141_, new_n24142_, new_n24143_, new_n24144_,
    new_n24145_, new_n24146_, new_n24147_, new_n24148_, new_n24149_,
    new_n24150_, new_n24151_, new_n24152_, new_n24153_, new_n24154_,
    new_n24155_, new_n24156_, new_n24157_, new_n24158_, new_n24159_,
    new_n24160_, new_n24161_, new_n24162_, new_n24163_, new_n24164_,
    new_n24165_, new_n24166_, new_n24167_, new_n24168_, new_n24169_,
    new_n24170_, new_n24171_, new_n24172_, new_n24173_, new_n24174_,
    new_n24175_, new_n24176_, new_n24177_, new_n24178_, new_n24179_,
    new_n24180_, new_n24181_, new_n24182_, new_n24183_, new_n24184_,
    new_n24185_, new_n24186_, new_n24187_, new_n24188_, new_n24189_,
    new_n24190_, new_n24191_, new_n24192_, new_n24193_, new_n24194_,
    new_n24195_, new_n24196_, new_n24197_, new_n24198_, new_n24199_,
    new_n24200_, new_n24201_, new_n24202_, new_n24203_, new_n24204_,
    new_n24205_, new_n24206_, new_n24207_, new_n24208_, new_n24209_,
    new_n24210_, new_n24211_, new_n24212_, new_n24213_, new_n24214_,
    new_n24215_, new_n24216_, new_n24217_, new_n24218_, new_n24219_,
    new_n24220_, new_n24221_, new_n24222_, new_n24223_, new_n24224_,
    new_n24225_, new_n24226_, new_n24227_, new_n24228_, new_n24229_,
    new_n24230_, new_n24231_, new_n24232_, new_n24233_, new_n24234_,
    new_n24235_, new_n24236_, new_n24237_, new_n24238_, new_n24239_,
    new_n24240_, new_n24241_, new_n24242_, new_n24243_, new_n24244_,
    new_n24245_, new_n24246_, new_n24247_, new_n24248_, new_n24249_,
    new_n24250_, new_n24251_, new_n24252_, new_n24253_, new_n24254_,
    new_n24255_, new_n24256_, new_n24257_, new_n24258_, new_n24259_,
    new_n24260_, new_n24261_, new_n24262_, new_n24263_, new_n24264_,
    new_n24265_, new_n24266_, new_n24267_, new_n24268_, new_n24269_,
    new_n24270_, new_n24271_, new_n24272_, new_n24273_, new_n24274_,
    new_n24275_, new_n24276_, new_n24277_, new_n24278_, new_n24279_,
    new_n24280_, new_n24281_, new_n24282_, new_n24283_, new_n24284_,
    new_n24285_, new_n24286_, new_n24287_, new_n24288_, new_n24289_,
    new_n24290_, new_n24291_, new_n24292_, new_n24293_, new_n24294_,
    new_n24295_, new_n24296_, new_n24297_, new_n24298_, new_n24299_,
    new_n24300_, new_n24301_, new_n24302_, new_n24303_, new_n24304_,
    new_n24305_, new_n24306_, new_n24307_, new_n24308_, new_n24309_,
    new_n24310_, new_n24311_, new_n24312_, new_n24313_, new_n24314_,
    new_n24315_, new_n24316_, new_n24317_, new_n24318_, new_n24319_,
    new_n24320_, new_n24321_, new_n24322_, new_n24323_, new_n24324_,
    new_n24325_, new_n24326_, new_n24327_, new_n24328_, new_n24329_,
    new_n24330_, new_n24331_, new_n24332_, new_n24333_, new_n24334_,
    new_n24335_, new_n24336_, new_n24337_, new_n24338_, new_n24339_,
    new_n24340_, new_n24341_, new_n24342_, new_n24343_, new_n24344_,
    new_n24345_, new_n24346_, new_n24347_, new_n24348_, new_n24349_,
    new_n24350_, new_n24351_, new_n24352_, new_n24353_, new_n24354_,
    new_n24355_, new_n24356_, new_n24357_, new_n24358_, new_n24359_,
    new_n24360_, new_n24361_, new_n24362_, new_n24363_, new_n24364_,
    new_n24365_, new_n24366_, new_n24367_, new_n24368_, new_n24369_,
    new_n24370_, new_n24371_, new_n24372_, new_n24373_, new_n24374_,
    new_n24375_, new_n24376_, new_n24377_, new_n24378_, new_n24379_,
    new_n24380_, new_n24381_, new_n24382_, new_n24383_, new_n24384_,
    new_n24385_, new_n24386_, new_n24387_, new_n24388_, new_n24389_,
    new_n24390_, new_n24391_, new_n24392_, new_n24393_, new_n24394_,
    new_n24395_, new_n24396_, new_n24397_, new_n24398_, new_n24399_,
    new_n24400_, new_n24401_, new_n24402_, new_n24403_, new_n24404_,
    new_n24405_, new_n24406_, new_n24407_, new_n24408_, new_n24409_,
    new_n24410_, new_n24411_, new_n24412_, new_n24413_, new_n24414_,
    new_n24415_, new_n24416_, new_n24417_, new_n24418_, new_n24419_,
    new_n24420_, new_n24421_, new_n24422_, new_n24423_, new_n24424_,
    new_n24425_, new_n24426_, new_n24427_, new_n24428_, new_n24429_,
    new_n24430_, new_n24431_, new_n24432_, new_n24433_, new_n24434_,
    new_n24435_, new_n24436_, new_n24437_, new_n24438_, new_n24439_,
    new_n24440_, new_n24441_, new_n24442_, new_n24443_, new_n24444_,
    new_n24445_, new_n24446_, new_n24447_, new_n24448_, new_n24449_,
    new_n24450_, new_n24451_, new_n24452_, new_n24453_, new_n24454_,
    new_n24455_, new_n24456_, new_n24457_, new_n24458_, new_n24459_,
    new_n24460_, new_n24461_, new_n24462_, new_n24463_, new_n24464_,
    new_n24465_, new_n24466_, new_n24467_, new_n24468_, new_n24469_,
    new_n24470_, new_n24471_, new_n24472_, new_n24473_, new_n24474_,
    new_n24475_, new_n24476_, new_n24477_, new_n24478_, new_n24479_,
    new_n24480_, new_n24481_, new_n24482_, new_n24483_, new_n24484_,
    new_n24485_, new_n24486_, new_n24487_, new_n24488_, new_n24489_,
    new_n24490_, new_n24491_, new_n24492_, new_n24493_, new_n24494_,
    new_n24495_, new_n24496_, new_n24497_, new_n24498_, new_n24499_,
    new_n24500_, new_n24501_, new_n24502_, new_n24503_, new_n24504_,
    new_n24505_, new_n24506_, new_n24507_, new_n24508_, new_n24509_,
    new_n24510_, new_n24511_, new_n24512_, new_n24513_, new_n24514_,
    new_n24515_, new_n24516_, new_n24517_, new_n24518_, new_n24519_,
    new_n24520_, new_n24521_, new_n24522_, new_n24523_, new_n24524_,
    new_n24525_, new_n24526_, new_n24527_, new_n24528_, new_n24529_,
    new_n24530_, new_n24531_, new_n24532_, new_n24533_, new_n24534_,
    new_n24535_, new_n24536_, new_n24537_, new_n24538_, new_n24539_,
    new_n24540_, new_n24541_, new_n24542_, new_n24543_, new_n24544_,
    new_n24545_, new_n24546_, new_n24547_, new_n24548_, new_n24549_,
    new_n24550_, new_n24551_, new_n24552_, new_n24553_, new_n24554_,
    new_n24555_, new_n24556_, new_n24557_, new_n24558_, new_n24559_,
    new_n24560_, new_n24561_, new_n24562_, new_n24563_, new_n24564_,
    new_n24565_, new_n24566_, new_n24567_, new_n24568_, new_n24569_,
    new_n24570_, new_n24571_, new_n24572_, new_n24573_, new_n24574_,
    new_n24575_, new_n24576_, new_n24577_, new_n24578_, new_n24579_,
    new_n24580_, new_n24581_, new_n24582_, new_n24583_, new_n24584_,
    new_n24585_, new_n24586_, new_n24587_, new_n24588_, new_n24589_,
    new_n24590_, new_n24591_, new_n24592_, new_n24593_, new_n24594_,
    new_n24595_, new_n24596_, new_n24597_, new_n24598_, new_n24599_,
    new_n24600_, new_n24601_, new_n24602_, new_n24603_, new_n24604_,
    new_n24605_, new_n24606_, new_n24607_, new_n24608_, new_n24609_,
    new_n24610_, new_n24611_, new_n24612_, new_n24613_, new_n24614_,
    new_n24615_, new_n24616_, new_n24617_, new_n24618_, new_n24619_,
    new_n24620_, new_n24621_, new_n24622_, new_n24623_, new_n24624_,
    new_n24625_, new_n24626_, new_n24627_, new_n24628_, new_n24629_,
    new_n24630_, new_n24631_, new_n24632_, new_n24633_, new_n24634_,
    new_n24635_, new_n24636_, new_n24637_, new_n24638_, new_n24639_,
    new_n24640_, new_n24641_, new_n24642_, new_n24643_, new_n24644_,
    new_n24645_, new_n24646_, new_n24647_, new_n24648_, new_n24649_,
    new_n24650_, new_n24651_, new_n24652_, new_n24653_, new_n24654_,
    new_n24655_, new_n24656_, new_n24657_, new_n24658_, new_n24659_,
    new_n24660_, new_n24661_, new_n24662_, new_n24663_, new_n24664_,
    new_n24665_, new_n24666_, new_n24667_, new_n24668_, new_n24669_,
    new_n24670_, new_n24671_, new_n24672_, new_n24673_, new_n24674_,
    new_n24675_, new_n24676_, new_n24677_, new_n24678_, new_n24679_,
    new_n24680_, new_n24681_, new_n24682_, new_n24683_, new_n24684_,
    new_n24685_, new_n24686_, new_n24687_, new_n24688_, new_n24689_,
    new_n24690_, new_n24691_, new_n24692_, new_n24693_, new_n24694_,
    new_n24695_, new_n24696_, new_n24697_, new_n24698_, new_n24699_,
    new_n24700_, new_n24701_, new_n24702_, new_n24703_, new_n24704_,
    new_n24705_, new_n24706_, new_n24707_, new_n24708_, new_n24709_,
    new_n24710_, new_n24711_, new_n24713_, new_n24714_, new_n24715_,
    new_n24716_, new_n24717_, new_n24718_, new_n24719_, new_n24720_,
    new_n24721_, new_n24722_, new_n24723_, new_n24724_, new_n24725_,
    new_n24726_, new_n24727_, new_n24728_, new_n24729_, new_n24730_,
    new_n24731_, new_n24732_, new_n24733_, new_n24734_, new_n24735_,
    new_n24736_, new_n24737_, new_n24738_, new_n24739_, new_n24740_,
    new_n24741_, new_n24742_, new_n24743_, new_n24744_, new_n24745_,
    new_n24746_, new_n24747_, new_n24748_, new_n24749_, new_n24750_,
    new_n24751_, new_n24752_, new_n24753_, new_n24754_, new_n24755_,
    new_n24756_, new_n24757_, new_n24758_, new_n24759_, new_n24760_,
    new_n24761_, new_n24762_, new_n24763_, new_n24764_, new_n24765_,
    new_n24766_, new_n24767_, new_n24768_, new_n24769_, new_n24770_,
    new_n24771_, new_n24772_, new_n24773_, new_n24774_, new_n24775_,
    new_n24776_, new_n24777_, new_n24778_, new_n24779_, new_n24780_,
    new_n24781_, new_n24782_, new_n24783_, new_n24784_, new_n24785_,
    new_n24786_, new_n24787_, new_n24788_, new_n24789_, new_n24790_,
    new_n24791_, new_n24792_, new_n24793_, new_n24794_, new_n24795_,
    new_n24796_, new_n24797_, new_n24798_, new_n24799_, new_n24800_,
    new_n24801_, new_n24802_, new_n24803_, new_n24804_, new_n24805_,
    new_n24806_, new_n24807_, new_n24808_, new_n24809_, new_n24810_,
    new_n24811_, new_n24812_, new_n24813_, new_n24814_, new_n24815_,
    new_n24816_, new_n24817_, new_n24818_, new_n24819_, new_n24820_,
    new_n24821_, new_n24822_, new_n24823_, new_n24824_, new_n24825_,
    new_n24826_, new_n24827_, new_n24828_, new_n24829_, new_n24830_,
    new_n24831_, new_n24832_, new_n24833_, new_n24834_, new_n24835_,
    new_n24836_, new_n24837_, new_n24838_, new_n24839_, new_n24840_,
    new_n24841_, new_n24842_, new_n24843_, new_n24844_, new_n24845_,
    new_n24846_, new_n24847_, new_n24848_, new_n24849_, new_n24850_,
    new_n24851_, new_n24852_, new_n24853_, new_n24854_, new_n24855_,
    new_n24856_, new_n24857_, new_n24858_, new_n24859_, new_n24860_,
    new_n24861_, new_n24862_, new_n24863_, new_n24864_, new_n24865_,
    new_n24866_, new_n24867_, new_n24868_, new_n24869_, new_n24870_,
    new_n24871_, new_n24872_, new_n24873_, new_n24874_, new_n24875_,
    new_n24876_, new_n24877_, new_n24878_, new_n24879_, new_n24880_,
    new_n24881_, new_n24882_, new_n24883_, new_n24884_, new_n24885_,
    new_n24886_, new_n24887_, new_n24888_, new_n24889_, new_n24890_,
    new_n24891_, new_n24892_, new_n24893_, new_n24894_, new_n24895_,
    new_n24896_, new_n24897_, new_n24898_, new_n24899_, new_n24900_,
    new_n24901_, new_n24902_, new_n24903_, new_n24904_, new_n24905_,
    new_n24906_, new_n24907_, new_n24908_, new_n24909_, new_n24910_,
    new_n24911_, new_n24912_, new_n24913_, new_n24914_, new_n24915_,
    new_n24916_, new_n24917_, new_n24918_, new_n24919_, new_n24920_,
    new_n24921_, new_n24922_, new_n24923_, new_n24924_, new_n24925_,
    new_n24926_, new_n24927_, new_n24928_, new_n24929_, new_n24930_,
    new_n24931_, new_n24932_, new_n24933_, new_n24934_, new_n24935_,
    new_n24936_, new_n24937_, new_n24938_, new_n24939_, new_n24940_,
    new_n24941_, new_n24942_, new_n24943_, new_n24944_, new_n24945_,
    new_n24946_, new_n24947_, new_n24948_, new_n24949_, new_n24950_,
    new_n24951_, new_n24952_, new_n24953_, new_n24954_, new_n24955_,
    new_n24956_, new_n24957_, new_n24958_, new_n24959_, new_n24960_,
    new_n24961_, new_n24962_, new_n24963_, new_n24964_, new_n24965_,
    new_n24966_, new_n24967_, new_n24968_, new_n24969_, new_n24970_,
    new_n24971_, new_n24972_, new_n24973_, new_n24974_, new_n24975_,
    new_n24976_, new_n24977_, new_n24978_, new_n24979_, new_n24980_,
    new_n24981_, new_n24982_, new_n24983_, new_n24984_, new_n24985_,
    new_n24986_, new_n24987_, new_n24988_, new_n24989_, new_n24990_,
    new_n24991_, new_n24992_, new_n24993_, new_n24994_, new_n24995_,
    new_n24996_, new_n24997_, new_n24998_, new_n24999_, new_n25000_,
    new_n25001_, new_n25002_, new_n25003_, new_n25004_, new_n25005_,
    new_n25006_, new_n25007_, new_n25008_, new_n25009_, new_n25010_,
    new_n25011_, new_n25012_, new_n25013_, new_n25014_, new_n25015_,
    new_n25016_, new_n25017_, new_n25018_, new_n25019_, new_n25020_,
    new_n25021_, new_n25022_, new_n25023_, new_n25024_, new_n25025_,
    new_n25026_, new_n25027_, new_n25028_, new_n25029_, new_n25030_,
    new_n25031_, new_n25032_, new_n25033_, new_n25034_, new_n25035_,
    new_n25036_, new_n25037_, new_n25038_, new_n25039_, new_n25040_,
    new_n25041_, new_n25042_, new_n25043_, new_n25044_, new_n25045_,
    new_n25046_, new_n25047_, new_n25048_, new_n25049_, new_n25050_,
    new_n25051_, new_n25052_, new_n25053_, new_n25054_, new_n25055_,
    new_n25056_, new_n25057_, new_n25058_, new_n25059_, new_n25060_,
    new_n25061_, new_n25062_, new_n25063_, new_n25064_, new_n25065_,
    new_n25066_, new_n25067_, new_n25068_, new_n25069_, new_n25070_,
    new_n25071_, new_n25072_, new_n25073_, new_n25074_, new_n25075_,
    new_n25076_, new_n25077_, new_n25078_, new_n25079_, new_n25080_,
    new_n25081_, new_n25082_, new_n25083_, new_n25084_, new_n25085_,
    new_n25086_, new_n25087_, new_n25088_, new_n25089_, new_n25090_,
    new_n25091_, new_n25092_, new_n25093_, new_n25094_, new_n25095_,
    new_n25096_, new_n25097_, new_n25098_, new_n25099_, new_n25100_,
    new_n25101_, new_n25102_, new_n25103_, new_n25104_, new_n25105_,
    new_n25106_, new_n25107_, new_n25108_, new_n25109_, new_n25110_,
    new_n25111_, new_n25112_, new_n25113_, new_n25114_, new_n25115_,
    new_n25116_, new_n25117_, new_n25118_, new_n25119_, new_n25120_,
    new_n25121_, new_n25122_, new_n25123_, new_n25124_, new_n25125_,
    new_n25126_, new_n25127_, new_n25128_, new_n25129_, new_n25130_,
    new_n25131_, new_n25132_, new_n25133_, new_n25134_, new_n25135_,
    new_n25136_, new_n25137_, new_n25138_, new_n25139_, new_n25140_,
    new_n25141_, new_n25142_, new_n25143_, new_n25144_, new_n25145_,
    new_n25146_, new_n25147_, new_n25148_, new_n25149_, new_n25150_,
    new_n25151_, new_n25152_, new_n25153_, new_n25154_, new_n25155_,
    new_n25156_, new_n25157_, new_n25158_, new_n25159_, new_n25160_,
    new_n25161_, new_n25162_, new_n25163_, new_n25164_, new_n25165_,
    new_n25166_, new_n25167_, new_n25168_, new_n25169_, new_n25170_,
    new_n25171_, new_n25172_, new_n25173_, new_n25174_, new_n25175_,
    new_n25176_, new_n25177_, new_n25178_, new_n25179_, new_n25180_,
    new_n25181_, new_n25182_, new_n25183_, new_n25184_, new_n25185_,
    new_n25186_, new_n25187_, new_n25188_, new_n25189_, new_n25190_,
    new_n25191_, new_n25192_, new_n25193_, new_n25194_, new_n25195_,
    new_n25196_, new_n25197_, new_n25198_, new_n25199_, new_n25200_,
    new_n25201_, new_n25202_, new_n25203_, new_n25204_, new_n25205_,
    new_n25206_, new_n25207_, new_n25208_, new_n25209_, new_n25210_,
    new_n25211_, new_n25212_, new_n25213_, new_n25214_, new_n25215_,
    new_n25216_, new_n25217_, new_n25218_, new_n25219_, new_n25220_,
    new_n25221_, new_n25222_, new_n25223_, new_n25224_, new_n25225_,
    new_n25226_, new_n25227_, new_n25228_, new_n25229_, new_n25230_,
    new_n25231_, new_n25232_, new_n25233_, new_n25234_, new_n25235_,
    new_n25236_, new_n25237_, new_n25238_, new_n25239_, new_n25240_,
    new_n25241_, new_n25242_, new_n25243_, new_n25244_, new_n25245_,
    new_n25246_, new_n25247_, new_n25248_, new_n25249_, new_n25250_,
    new_n25251_, new_n25252_, new_n25253_, new_n25254_, new_n25255_,
    new_n25256_, new_n25257_, new_n25258_, new_n25259_, new_n25260_,
    new_n25261_, new_n25262_, new_n25263_, new_n25264_, new_n25265_,
    new_n25266_, new_n25267_, new_n25268_, new_n25269_, new_n25270_,
    new_n25271_, new_n25272_, new_n25273_, new_n25274_, new_n25275_,
    new_n25276_, new_n25277_, new_n25278_, new_n25279_, new_n25280_,
    new_n25281_, new_n25282_, new_n25283_, new_n25284_, new_n25285_,
    new_n25286_, new_n25287_, new_n25288_, new_n25289_, new_n25290_,
    new_n25291_, new_n25292_, new_n25293_, new_n25294_, new_n25295_,
    new_n25296_, new_n25297_, new_n25298_, new_n25299_, new_n25300_,
    new_n25301_, new_n25302_, new_n25303_, new_n25304_, new_n25305_,
    new_n25306_, new_n25307_, new_n25308_, new_n25309_, new_n25310_,
    new_n25311_, new_n25312_, new_n25313_, new_n25314_, new_n25315_,
    new_n25316_, new_n25317_, new_n25318_, new_n25319_, new_n25320_,
    new_n25321_, new_n25322_, new_n25323_, new_n25324_, new_n25325_,
    new_n25326_, new_n25327_, new_n25328_, new_n25329_, new_n25330_,
    new_n25331_, new_n25332_, new_n25333_, new_n25334_, new_n25335_,
    new_n25336_, new_n25337_, new_n25338_, new_n25339_, new_n25340_,
    new_n25341_, new_n25342_, new_n25343_, new_n25344_, new_n25345_,
    new_n25346_, new_n25347_, new_n25348_, new_n25349_, new_n25350_,
    new_n25351_, new_n25352_, new_n25353_, new_n25354_, new_n25355_,
    new_n25356_, new_n25357_, new_n25358_, new_n25359_, new_n25360_,
    new_n25361_, new_n25362_, new_n25363_, new_n25364_, new_n25365_,
    new_n25366_, new_n25367_, new_n25368_, new_n25369_, new_n25370_,
    new_n25371_, new_n25372_, new_n25373_, new_n25374_, new_n25375_,
    new_n25376_, new_n25377_, new_n25378_, new_n25379_, new_n25380_,
    new_n25381_, new_n25382_, new_n25383_, new_n25384_, new_n25385_,
    new_n25386_, new_n25387_, new_n25388_, new_n25389_, new_n25390_,
    new_n25391_, new_n25392_, new_n25393_, new_n25394_, new_n25395_,
    new_n25396_, new_n25397_, new_n25398_, new_n25399_, new_n25400_,
    new_n25401_, new_n25402_, new_n25403_, new_n25404_, new_n25405_,
    new_n25406_, new_n25407_, new_n25408_, new_n25409_, new_n25410_,
    new_n25411_, new_n25412_, new_n25413_, new_n25414_, new_n25415_,
    new_n25416_, new_n25417_, new_n25418_, new_n25419_, new_n25420_,
    new_n25421_, new_n25422_, new_n25423_, new_n25424_, new_n25425_,
    new_n25426_, new_n25427_, new_n25428_, new_n25429_, new_n25430_,
    new_n25431_, new_n25432_, new_n25433_, new_n25434_, new_n25435_,
    new_n25436_, new_n25437_, new_n25438_, new_n25439_, new_n25440_,
    new_n25441_, new_n25442_, new_n25443_, new_n25444_, new_n25445_,
    new_n25446_, new_n25447_, new_n25448_, new_n25449_, new_n25450_,
    new_n25451_, new_n25452_, new_n25453_, new_n25454_, new_n25455_,
    new_n25456_, new_n25457_, new_n25458_, new_n25459_, new_n25460_,
    new_n25461_, new_n25462_, new_n25463_, new_n25464_, new_n25465_,
    new_n25466_, new_n25467_, new_n25468_, new_n25469_, new_n25470_,
    new_n25471_, new_n25472_, new_n25473_, new_n25474_, new_n25475_,
    new_n25476_, new_n25477_, new_n25478_, new_n25479_, new_n25480_,
    new_n25481_, new_n25482_, new_n25483_, new_n25484_, new_n25485_,
    new_n25486_, new_n25487_, new_n25488_, new_n25489_, new_n25490_,
    new_n25491_, new_n25492_, new_n25493_, new_n25494_, new_n25495_,
    new_n25496_, new_n25497_, new_n25498_, new_n25499_, new_n25500_,
    new_n25501_, new_n25502_, new_n25503_, new_n25504_, new_n25505_,
    new_n25506_, new_n25507_, new_n25508_, new_n25509_, new_n25510_,
    new_n25511_, new_n25512_, new_n25513_, new_n25514_, new_n25515_,
    new_n25516_, new_n25517_, new_n25518_, new_n25519_, new_n25520_,
    new_n25521_, new_n25522_, new_n25523_, new_n25524_, new_n25525_,
    new_n25526_, new_n25527_, new_n25528_, new_n25529_, new_n25530_,
    new_n25531_, new_n25532_, new_n25533_, new_n25534_, new_n25535_,
    new_n25536_, new_n25537_, new_n25538_, new_n25540_, new_n25541_,
    new_n25542_, new_n25543_, new_n25544_, new_n25545_, new_n25546_,
    new_n25547_, new_n25548_, new_n25549_, new_n25550_, new_n25551_,
    new_n25552_, new_n25553_, new_n25554_, new_n25555_, new_n25556_,
    new_n25557_, new_n25558_, new_n25559_, new_n25560_, new_n25561_,
    new_n25562_, new_n25563_, new_n25564_, new_n25565_, new_n25566_,
    new_n25567_, new_n25568_, new_n25569_, new_n25570_, new_n25571_,
    new_n25572_, new_n25573_, new_n25574_, new_n25575_, new_n25576_,
    new_n25577_, new_n25578_, new_n25579_, new_n25580_, new_n25581_,
    new_n25582_, new_n25583_, new_n25584_, new_n25585_, new_n25586_,
    new_n25587_, new_n25588_, new_n25589_, new_n25590_, new_n25591_,
    new_n25592_, new_n25593_, new_n25594_, new_n25595_, new_n25596_,
    new_n25597_, new_n25598_, new_n25599_, new_n25600_, new_n25601_,
    new_n25602_, new_n25603_, new_n25604_, new_n25605_, new_n25606_,
    new_n25607_, new_n25608_, new_n25609_, new_n25610_, new_n25611_,
    new_n25612_, new_n25613_, new_n25614_, new_n25615_, new_n25616_,
    new_n25617_, new_n25618_, new_n25619_, new_n25620_, new_n25621_,
    new_n25622_, new_n25623_, new_n25624_, new_n25625_, new_n25626_,
    new_n25627_, new_n25628_, new_n25629_, new_n25630_, new_n25631_,
    new_n25632_, new_n25633_, new_n25634_, new_n25635_, new_n25636_,
    new_n25637_, new_n25638_, new_n25639_, new_n25640_, new_n25641_,
    new_n25642_, new_n25643_, new_n25644_, new_n25645_, new_n25646_,
    new_n25647_, new_n25648_, new_n25649_, new_n25650_, new_n25651_,
    new_n25652_, new_n25653_, new_n25654_, new_n25655_, new_n25656_,
    new_n25657_, new_n25658_, new_n25659_, new_n25660_, new_n25661_,
    new_n25662_, new_n25663_, new_n25664_, new_n25665_, new_n25666_,
    new_n25667_, new_n25668_, new_n25669_, new_n25670_, new_n25671_,
    new_n25672_, new_n25673_, new_n25674_, new_n25675_, new_n25676_,
    new_n25677_, new_n25678_, new_n25679_, new_n25680_, new_n25681_,
    new_n25682_, new_n25683_, new_n25684_, new_n25685_, new_n25686_,
    new_n25687_, new_n25688_, new_n25689_, new_n25690_, new_n25691_,
    new_n25692_, new_n25693_, new_n25694_, new_n25695_, new_n25696_,
    new_n25697_, new_n25698_, new_n25699_, new_n25700_, new_n25701_,
    new_n25702_, new_n25703_, new_n25704_, new_n25705_, new_n25706_,
    new_n25707_, new_n25708_, new_n25709_, new_n25710_, new_n25711_,
    new_n25712_, new_n25713_, new_n25714_, new_n25715_, new_n25716_,
    new_n25717_, new_n25718_, new_n25719_, new_n25720_, new_n25721_,
    new_n25722_, new_n25723_, new_n25724_, new_n25725_, new_n25726_,
    new_n25727_, new_n25728_, new_n25729_, new_n25730_, new_n25731_,
    new_n25732_, new_n25733_, new_n25734_, new_n25735_, new_n25736_,
    new_n25737_, new_n25738_, new_n25739_, new_n25740_, new_n25741_,
    new_n25742_, new_n25743_, new_n25744_, new_n25745_, new_n25746_,
    new_n25747_, new_n25748_, new_n25749_, new_n25750_, new_n25751_,
    new_n25752_, new_n25753_, new_n25754_, new_n25755_, new_n25756_,
    new_n25757_, new_n25758_, new_n25759_, new_n25760_, new_n25761_,
    new_n25762_, new_n25763_, new_n25764_, new_n25765_, new_n25766_,
    new_n25767_, new_n25768_, new_n25769_, new_n25770_, new_n25771_,
    new_n25772_, new_n25773_, new_n25774_, new_n25775_, new_n25776_,
    new_n25777_, new_n25778_, new_n25779_, new_n25780_, new_n25781_,
    new_n25782_, new_n25783_, new_n25784_, new_n25785_, new_n25786_,
    new_n25787_, new_n25788_, new_n25789_, new_n25790_, new_n25791_,
    new_n25792_, new_n25793_, new_n25794_, new_n25795_, new_n25796_,
    new_n25797_, new_n25798_, new_n25799_, new_n25800_, new_n25801_,
    new_n25802_, new_n25803_, new_n25804_, new_n25805_, new_n25806_,
    new_n25807_, new_n25808_, new_n25809_, new_n25810_, new_n25811_,
    new_n25812_, new_n25813_, new_n25814_, new_n25815_, new_n25816_,
    new_n25817_, new_n25818_, new_n25819_, new_n25820_, new_n25821_,
    new_n25822_, new_n25823_, new_n25824_, new_n25825_, new_n25826_,
    new_n25827_, new_n25828_, new_n25829_, new_n25830_, new_n25831_,
    new_n25832_, new_n25833_, new_n25834_, new_n25835_, new_n25836_,
    new_n25837_, new_n25838_, new_n25839_, new_n25840_, new_n25841_,
    new_n25842_, new_n25843_, new_n25844_, new_n25845_, new_n25846_,
    new_n25847_, new_n25848_, new_n25849_, new_n25850_, new_n25851_,
    new_n25852_, new_n25853_, new_n25854_, new_n25855_, new_n25856_,
    new_n25857_, new_n25858_, new_n25859_, new_n25860_, new_n25861_,
    new_n25862_, new_n25863_, new_n25864_, new_n25865_, new_n25866_,
    new_n25867_, new_n25868_, new_n25869_, new_n25870_, new_n25871_,
    new_n25872_, new_n25873_, new_n25874_, new_n25875_, new_n25876_,
    new_n25877_, new_n25878_, new_n25879_, new_n25880_, new_n25881_,
    new_n25882_, new_n25883_, new_n25884_, new_n25885_, new_n25886_,
    new_n25887_, new_n25888_, new_n25889_, new_n25890_, new_n25891_,
    new_n25892_, new_n25893_, new_n25894_, new_n25895_, new_n25896_,
    new_n25897_, new_n25898_, new_n25899_, new_n25900_, new_n25901_,
    new_n25902_, new_n25903_, new_n25904_, new_n25905_, new_n25906_,
    new_n25907_, new_n25908_, new_n25909_, new_n25910_, new_n25911_,
    new_n25912_, new_n25913_, new_n25914_, new_n25915_, new_n25916_,
    new_n25917_, new_n25918_, new_n25919_, new_n25920_, new_n25921_,
    new_n25922_, new_n25923_, new_n25924_, new_n25925_, new_n25926_,
    new_n25927_, new_n25928_, new_n25929_, new_n25930_, new_n25931_,
    new_n25932_, new_n25933_, new_n25934_, new_n25935_, new_n25936_,
    new_n25937_, new_n25938_, new_n25939_, new_n25940_, new_n25941_,
    new_n25942_, new_n25943_, new_n25944_, new_n25945_, new_n25946_,
    new_n25947_, new_n25948_, new_n25949_, new_n25950_, new_n25951_,
    new_n25952_, new_n25953_, new_n25954_, new_n25955_, new_n25956_,
    new_n25957_, new_n25958_, new_n25959_, new_n25960_, new_n25961_,
    new_n25962_, new_n25963_, new_n25964_, new_n25965_, new_n25966_,
    new_n25967_, new_n25968_, new_n25969_, new_n25970_, new_n25971_,
    new_n25972_, new_n25973_, new_n25974_, new_n25975_, new_n25976_,
    new_n25977_, new_n25978_, new_n25979_, new_n25980_, new_n25981_,
    new_n25982_, new_n25983_, new_n25984_, new_n25985_, new_n25986_,
    new_n25987_, new_n25988_, new_n25989_, new_n25990_, new_n25991_,
    new_n25992_, new_n25993_, new_n25994_, new_n25995_, new_n25996_,
    new_n25997_, new_n25998_, new_n25999_, new_n26000_, new_n26001_,
    new_n26002_, new_n26003_, new_n26004_, new_n26005_, new_n26006_,
    new_n26007_, new_n26008_, new_n26009_, new_n26010_, new_n26011_,
    new_n26012_, new_n26013_, new_n26014_, new_n26015_, new_n26016_,
    new_n26017_, new_n26018_, new_n26019_, new_n26020_, new_n26021_,
    new_n26022_, new_n26023_, new_n26024_, new_n26025_, new_n26026_,
    new_n26027_, new_n26028_, new_n26029_, new_n26030_, new_n26031_,
    new_n26032_, new_n26033_, new_n26034_, new_n26035_, new_n26036_,
    new_n26037_, new_n26038_, new_n26039_, new_n26040_, new_n26041_,
    new_n26042_, new_n26043_, new_n26044_, new_n26045_, new_n26046_,
    new_n26047_, new_n26048_, new_n26049_, new_n26050_, new_n26051_,
    new_n26052_, new_n26053_, new_n26054_, new_n26055_, new_n26056_,
    new_n26057_, new_n26058_, new_n26059_, new_n26060_, new_n26061_,
    new_n26062_, new_n26063_, new_n26064_, new_n26065_, new_n26066_,
    new_n26067_, new_n26068_, new_n26069_, new_n26070_, new_n26071_,
    new_n26072_, new_n26073_, new_n26074_, new_n26075_, new_n26076_,
    new_n26077_, new_n26078_, new_n26079_, new_n26080_, new_n26081_,
    new_n26082_, new_n26083_, new_n26084_, new_n26085_, new_n26086_,
    new_n26087_, new_n26088_, new_n26089_, new_n26090_, new_n26091_,
    new_n26092_, new_n26093_, new_n26094_, new_n26095_, new_n26096_,
    new_n26097_, new_n26098_, new_n26099_, new_n26100_, new_n26101_,
    new_n26102_, new_n26103_, new_n26104_, new_n26105_, new_n26106_,
    new_n26107_, new_n26108_, new_n26109_, new_n26110_, new_n26111_,
    new_n26112_, new_n26113_, new_n26114_, new_n26115_, new_n26116_,
    new_n26117_, new_n26118_, new_n26119_, new_n26120_, new_n26121_,
    new_n26122_, new_n26123_, new_n26124_, new_n26125_, new_n26126_,
    new_n26127_, new_n26128_, new_n26129_, new_n26130_, new_n26131_,
    new_n26132_, new_n26133_, new_n26134_, new_n26135_, new_n26136_,
    new_n26137_, new_n26138_, new_n26139_, new_n26140_, new_n26141_,
    new_n26142_, new_n26143_, new_n26144_, new_n26145_, new_n26146_,
    new_n26147_, new_n26148_, new_n26149_, new_n26150_, new_n26151_,
    new_n26152_, new_n26153_, new_n26154_, new_n26155_, new_n26156_,
    new_n26157_, new_n26158_, new_n26159_, new_n26160_, new_n26161_,
    new_n26162_, new_n26163_, new_n26164_, new_n26165_, new_n26166_,
    new_n26167_, new_n26168_, new_n26169_, new_n26170_, new_n26171_,
    new_n26172_, new_n26173_, new_n26174_, new_n26175_, new_n26176_,
    new_n26177_, new_n26178_, new_n26179_, new_n26180_, new_n26181_,
    new_n26182_, new_n26183_, new_n26184_, new_n26185_, new_n26186_,
    new_n26187_, new_n26188_, new_n26189_, new_n26190_, new_n26191_,
    new_n26192_, new_n26193_, new_n26194_, new_n26195_, new_n26196_,
    new_n26197_, new_n26198_, new_n26199_, new_n26200_, new_n26201_,
    new_n26202_, new_n26203_, new_n26204_, new_n26205_, new_n26206_,
    new_n26207_, new_n26208_, new_n26209_, new_n26210_, new_n26211_,
    new_n26212_, new_n26213_, new_n26214_, new_n26215_, new_n26216_,
    new_n26217_, new_n26218_, new_n26219_, new_n26220_, new_n26221_,
    new_n26222_, new_n26223_, new_n26224_, new_n26225_, new_n26226_,
    new_n26227_, new_n26228_, new_n26229_, new_n26230_, new_n26231_,
    new_n26232_, new_n26233_, new_n26234_, new_n26235_, new_n26236_,
    new_n26237_, new_n26238_, new_n26239_, new_n26240_, new_n26241_,
    new_n26242_, new_n26243_, new_n26244_, new_n26245_, new_n26246_,
    new_n26247_, new_n26248_, new_n26249_, new_n26250_, new_n26251_,
    new_n26252_, new_n26253_, new_n26254_, new_n26255_, new_n26256_,
    new_n26257_, new_n26258_, new_n26259_, new_n26260_, new_n26261_,
    new_n26262_, new_n26263_, new_n26264_, new_n26265_, new_n26266_,
    new_n26267_, new_n26268_, new_n26269_, new_n26270_, new_n26271_,
    new_n26272_, new_n26273_, new_n26274_, new_n26275_, new_n26276_,
    new_n26277_, new_n26278_, new_n26279_, new_n26280_, new_n26281_,
    new_n26282_, new_n26283_, new_n26284_, new_n26285_, new_n26286_,
    new_n26287_, new_n26288_, new_n26289_, new_n26290_, new_n26291_,
    new_n26292_, new_n26293_, new_n26294_, new_n26295_, new_n26296_,
    new_n26297_, new_n26298_, new_n26299_, new_n26300_, new_n26301_,
    new_n26302_, new_n26303_, new_n26304_, new_n26305_, new_n26306_,
    new_n26307_, new_n26308_, new_n26309_, new_n26310_, new_n26311_,
    new_n26312_, new_n26313_, new_n26314_, new_n26315_, new_n26316_,
    new_n26317_, new_n26318_, new_n26319_, new_n26320_, new_n26321_,
    new_n26322_, new_n26323_, new_n26324_, new_n26325_, new_n26326_,
    new_n26327_, new_n26328_, new_n26329_, new_n26330_, new_n26331_,
    new_n26332_, new_n26333_, new_n26334_, new_n26335_, new_n26336_,
    new_n26337_, new_n26338_, new_n26339_, new_n26340_, new_n26341_,
    new_n26342_, new_n26343_, new_n26344_, new_n26345_, new_n26346_,
    new_n26347_, new_n26348_, new_n26349_, new_n26350_, new_n26351_,
    new_n26352_, new_n26353_, new_n26354_, new_n26355_, new_n26356_,
    new_n26357_, new_n26358_, new_n26359_, new_n26360_, new_n26361_,
    new_n26362_, new_n26363_, new_n26364_, new_n26365_, new_n26366_,
    new_n26367_, new_n26368_, new_n26369_, new_n26370_, new_n26371_,
    new_n26372_, new_n26373_, new_n26374_, new_n26375_, new_n26376_,
    new_n26377_, new_n26378_, new_n26379_, new_n26381_, new_n26382_,
    new_n26383_, new_n26384_, new_n26385_, new_n26386_, new_n26387_,
    new_n26388_, new_n26389_, new_n26390_, new_n26391_, new_n26392_,
    new_n26393_, new_n26394_, new_n26395_, new_n26396_, new_n26397_,
    new_n26398_, new_n26399_, new_n26400_, new_n26401_, new_n26402_,
    new_n26403_, new_n26404_, new_n26405_, new_n26406_, new_n26407_,
    new_n26408_, new_n26409_, new_n26410_, new_n26411_, new_n26412_,
    new_n26413_, new_n26414_, new_n26415_, new_n26416_, new_n26417_,
    new_n26418_, new_n26419_, new_n26420_, new_n26421_, new_n26422_,
    new_n26423_, new_n26424_, new_n26425_, new_n26426_, new_n26427_,
    new_n26428_, new_n26429_, new_n26430_, new_n26431_, new_n26432_,
    new_n26433_, new_n26434_, new_n26435_, new_n26436_, new_n26437_,
    new_n26438_, new_n26439_, new_n26440_, new_n26441_, new_n26442_,
    new_n26443_, new_n26444_, new_n26445_, new_n26446_, new_n26447_,
    new_n26448_, new_n26449_, new_n26450_, new_n26451_, new_n26452_,
    new_n26453_, new_n26454_, new_n26455_, new_n26456_, new_n26457_,
    new_n26458_, new_n26459_, new_n26460_, new_n26461_, new_n26462_,
    new_n26463_, new_n26464_, new_n26465_, new_n26466_, new_n26467_,
    new_n26468_, new_n26469_, new_n26470_, new_n26471_, new_n26472_,
    new_n26473_, new_n26474_, new_n26475_, new_n26476_, new_n26477_,
    new_n26478_, new_n26479_, new_n26480_, new_n26481_, new_n26482_,
    new_n26483_, new_n26484_, new_n26485_, new_n26486_, new_n26487_,
    new_n26488_, new_n26489_, new_n26490_, new_n26491_, new_n26492_,
    new_n26493_, new_n26494_, new_n26495_, new_n26496_, new_n26497_,
    new_n26498_, new_n26499_, new_n26500_, new_n26501_, new_n26502_,
    new_n26503_, new_n26504_, new_n26505_, new_n26506_, new_n26507_,
    new_n26508_, new_n26509_, new_n26510_, new_n26511_, new_n26512_,
    new_n26513_, new_n26514_, new_n26515_, new_n26516_, new_n26517_,
    new_n26518_, new_n26519_, new_n26520_, new_n26521_, new_n26522_,
    new_n26523_, new_n26524_, new_n26525_, new_n26526_, new_n26527_,
    new_n26528_, new_n26529_, new_n26530_, new_n26531_, new_n26532_,
    new_n26533_, new_n26534_, new_n26535_, new_n26536_, new_n26537_,
    new_n26538_, new_n26539_, new_n26540_, new_n26541_, new_n26542_,
    new_n26543_, new_n26544_, new_n26545_, new_n26546_, new_n26547_,
    new_n26548_, new_n26549_, new_n26550_, new_n26551_, new_n26552_,
    new_n26553_, new_n26554_, new_n26555_, new_n26556_, new_n26557_,
    new_n26558_, new_n26559_, new_n26560_, new_n26561_, new_n26562_,
    new_n26563_, new_n26564_, new_n26565_, new_n26566_, new_n26567_,
    new_n26568_, new_n26569_, new_n26570_, new_n26571_, new_n26572_,
    new_n26573_, new_n26574_, new_n26575_, new_n26576_, new_n26577_,
    new_n26578_, new_n26579_, new_n26580_, new_n26581_, new_n26582_,
    new_n26583_, new_n26584_, new_n26585_, new_n26586_, new_n26587_,
    new_n26588_, new_n26589_, new_n26590_, new_n26591_, new_n26592_,
    new_n26593_, new_n26594_, new_n26595_, new_n26596_, new_n26597_,
    new_n26598_, new_n26599_, new_n26600_, new_n26601_, new_n26602_,
    new_n26603_, new_n26604_, new_n26605_, new_n26606_, new_n26607_,
    new_n26608_, new_n26609_, new_n26610_, new_n26611_, new_n26612_,
    new_n26613_, new_n26614_, new_n26615_, new_n26616_, new_n26617_,
    new_n26618_, new_n26619_, new_n26620_, new_n26621_, new_n26622_,
    new_n26623_, new_n26624_, new_n26625_, new_n26626_, new_n26627_,
    new_n26628_, new_n26629_, new_n26630_, new_n26631_, new_n26632_,
    new_n26633_, new_n26634_, new_n26635_, new_n26636_, new_n26637_,
    new_n26638_, new_n26639_, new_n26640_, new_n26641_, new_n26642_,
    new_n26643_, new_n26644_, new_n26645_, new_n26646_, new_n26647_,
    new_n26648_, new_n26649_, new_n26650_, new_n26651_, new_n26652_,
    new_n26653_, new_n26654_, new_n26655_, new_n26656_, new_n26657_,
    new_n26658_, new_n26659_, new_n26660_, new_n26661_, new_n26662_,
    new_n26663_, new_n26664_, new_n26665_, new_n26666_, new_n26667_,
    new_n26668_, new_n26669_, new_n26670_, new_n26671_, new_n26672_,
    new_n26673_, new_n26674_, new_n26675_, new_n26676_, new_n26677_,
    new_n26678_, new_n26679_, new_n26680_, new_n26681_, new_n26682_,
    new_n26683_, new_n26684_, new_n26685_, new_n26686_, new_n26687_,
    new_n26688_, new_n26689_, new_n26690_, new_n26691_, new_n26692_,
    new_n26693_, new_n26694_, new_n26695_, new_n26696_, new_n26697_,
    new_n26698_, new_n26699_, new_n26700_, new_n26701_, new_n26702_,
    new_n26703_, new_n26704_, new_n26705_, new_n26706_, new_n26707_,
    new_n26708_, new_n26709_, new_n26710_, new_n26711_, new_n26712_,
    new_n26713_, new_n26714_, new_n26715_, new_n26716_, new_n26717_,
    new_n26718_, new_n26719_, new_n26720_, new_n26721_, new_n26722_,
    new_n26723_, new_n26724_, new_n26725_, new_n26726_, new_n26727_,
    new_n26728_, new_n26729_, new_n26730_, new_n26731_, new_n26732_,
    new_n26733_, new_n26734_, new_n26735_, new_n26736_, new_n26737_,
    new_n26738_, new_n26739_, new_n26740_, new_n26741_, new_n26742_,
    new_n26743_, new_n26744_, new_n26745_, new_n26746_, new_n26747_,
    new_n26748_, new_n26749_, new_n26750_, new_n26751_, new_n26752_,
    new_n26753_, new_n26754_, new_n26755_, new_n26756_, new_n26757_,
    new_n26758_, new_n26759_, new_n26760_, new_n26761_, new_n26762_,
    new_n26763_, new_n26764_, new_n26765_, new_n26766_, new_n26767_,
    new_n26768_, new_n26769_, new_n26770_, new_n26771_, new_n26772_,
    new_n26773_, new_n26774_, new_n26775_, new_n26776_, new_n26777_,
    new_n26778_, new_n26779_, new_n26780_, new_n26781_, new_n26782_,
    new_n26783_, new_n26784_, new_n26785_, new_n26786_, new_n26787_,
    new_n26788_, new_n26789_, new_n26790_, new_n26791_, new_n26792_,
    new_n26793_, new_n26794_, new_n26795_, new_n26796_, new_n26797_,
    new_n26798_, new_n26799_, new_n26800_, new_n26801_, new_n26802_,
    new_n26803_, new_n26804_, new_n26805_, new_n26806_, new_n26807_,
    new_n26808_, new_n26809_, new_n26810_, new_n26811_, new_n26812_,
    new_n26813_, new_n26814_, new_n26815_, new_n26816_, new_n26817_,
    new_n26818_, new_n26819_, new_n26820_, new_n26821_, new_n26822_,
    new_n26823_, new_n26824_, new_n26825_, new_n26826_, new_n26827_,
    new_n26828_, new_n26829_, new_n26830_, new_n26831_, new_n26832_,
    new_n26833_, new_n26834_, new_n26835_, new_n26836_, new_n26837_,
    new_n26838_, new_n26839_, new_n26840_, new_n26841_, new_n26842_,
    new_n26843_, new_n26844_, new_n26845_, new_n26846_, new_n26847_,
    new_n26848_, new_n26849_, new_n26850_, new_n26851_, new_n26852_,
    new_n26853_, new_n26854_, new_n26855_, new_n26856_, new_n26857_,
    new_n26858_, new_n26859_, new_n26860_, new_n26861_, new_n26862_,
    new_n26863_, new_n26864_, new_n26865_, new_n26866_, new_n26867_,
    new_n26868_, new_n26869_, new_n26870_, new_n26871_, new_n26872_,
    new_n26873_, new_n26874_, new_n26875_, new_n26876_, new_n26877_,
    new_n26878_, new_n26879_, new_n26880_, new_n26881_, new_n26882_,
    new_n26883_, new_n26884_, new_n26885_, new_n26886_, new_n26887_,
    new_n26888_, new_n26889_, new_n26890_, new_n26891_, new_n26892_,
    new_n26893_, new_n26894_, new_n26895_, new_n26896_, new_n26897_,
    new_n26898_, new_n26899_, new_n26900_, new_n26901_, new_n26902_,
    new_n26903_, new_n26904_, new_n26905_, new_n26906_, new_n26907_,
    new_n26908_, new_n26909_, new_n26910_, new_n26911_, new_n26912_,
    new_n26913_, new_n26914_, new_n26915_, new_n26916_, new_n26917_,
    new_n26918_, new_n26919_, new_n26920_, new_n26921_, new_n26922_,
    new_n26923_, new_n26924_, new_n26925_, new_n26926_, new_n26927_,
    new_n26928_, new_n26929_, new_n26930_, new_n26931_, new_n26932_,
    new_n26933_, new_n26934_, new_n26935_, new_n26936_, new_n26937_,
    new_n26938_, new_n26939_, new_n26940_, new_n26941_, new_n26942_,
    new_n26943_, new_n26944_, new_n26945_, new_n26946_, new_n26947_,
    new_n26948_, new_n26949_, new_n26950_, new_n26951_, new_n26952_,
    new_n26953_, new_n26954_, new_n26955_, new_n26956_, new_n26957_,
    new_n26958_, new_n26959_, new_n26960_, new_n26961_, new_n26962_,
    new_n26963_, new_n26964_, new_n26965_, new_n26966_, new_n26967_,
    new_n26968_, new_n26969_, new_n26970_, new_n26971_, new_n26972_,
    new_n26973_, new_n26974_, new_n26975_, new_n26976_, new_n26977_,
    new_n26978_, new_n26979_, new_n26980_, new_n26981_, new_n26982_,
    new_n26983_, new_n26984_, new_n26985_, new_n26986_, new_n26987_,
    new_n26988_, new_n26989_, new_n26990_, new_n26991_, new_n26992_,
    new_n26993_, new_n26994_, new_n26995_, new_n26996_, new_n26997_,
    new_n26998_, new_n26999_, new_n27000_, new_n27001_, new_n27002_,
    new_n27003_, new_n27004_, new_n27005_, new_n27006_, new_n27007_,
    new_n27008_, new_n27009_, new_n27010_, new_n27011_, new_n27012_,
    new_n27013_, new_n27014_, new_n27015_, new_n27016_, new_n27017_,
    new_n27018_, new_n27019_, new_n27020_, new_n27021_, new_n27022_,
    new_n27023_, new_n27024_, new_n27025_, new_n27026_, new_n27027_,
    new_n27028_, new_n27029_, new_n27030_, new_n27031_, new_n27032_,
    new_n27033_, new_n27034_, new_n27035_, new_n27036_, new_n27037_,
    new_n27038_, new_n27039_, new_n27040_, new_n27041_, new_n27042_,
    new_n27043_, new_n27044_, new_n27045_, new_n27046_, new_n27047_,
    new_n27048_, new_n27049_, new_n27050_, new_n27051_, new_n27052_,
    new_n27053_, new_n27054_, new_n27055_, new_n27056_, new_n27057_,
    new_n27058_, new_n27059_, new_n27060_, new_n27061_, new_n27062_,
    new_n27063_, new_n27064_, new_n27065_, new_n27066_, new_n27067_,
    new_n27068_, new_n27069_, new_n27070_, new_n27071_, new_n27072_,
    new_n27073_, new_n27074_, new_n27075_, new_n27076_, new_n27077_,
    new_n27078_, new_n27079_, new_n27080_, new_n27081_, new_n27082_,
    new_n27083_, new_n27084_, new_n27085_, new_n27086_, new_n27087_,
    new_n27088_, new_n27089_, new_n27090_, new_n27091_, new_n27092_,
    new_n27093_, new_n27094_, new_n27095_, new_n27096_, new_n27097_,
    new_n27098_, new_n27099_, new_n27100_, new_n27101_, new_n27102_,
    new_n27103_, new_n27104_, new_n27105_, new_n27106_, new_n27107_,
    new_n27108_, new_n27109_, new_n27110_, new_n27111_, new_n27112_,
    new_n27113_, new_n27114_, new_n27115_, new_n27116_, new_n27117_,
    new_n27118_, new_n27119_, new_n27120_, new_n27121_, new_n27122_,
    new_n27123_, new_n27124_, new_n27125_, new_n27126_, new_n27127_,
    new_n27128_, new_n27129_, new_n27130_, new_n27131_, new_n27132_,
    new_n27133_, new_n27134_, new_n27135_, new_n27136_, new_n27137_,
    new_n27138_, new_n27139_, new_n27140_, new_n27141_, new_n27142_,
    new_n27143_, new_n27144_, new_n27145_, new_n27146_, new_n27147_,
    new_n27148_, new_n27149_, new_n27150_, new_n27151_, new_n27152_,
    new_n27153_, new_n27154_, new_n27155_, new_n27156_, new_n27157_,
    new_n27158_, new_n27159_, new_n27160_, new_n27161_, new_n27162_,
    new_n27163_, new_n27164_, new_n27165_, new_n27166_, new_n27167_,
    new_n27168_, new_n27169_, new_n27170_, new_n27171_, new_n27172_,
    new_n27173_, new_n27174_, new_n27175_, new_n27176_, new_n27177_,
    new_n27178_, new_n27179_, new_n27180_, new_n27181_, new_n27182_,
    new_n27183_, new_n27184_, new_n27185_, new_n27186_, new_n27187_,
    new_n27188_, new_n27189_, new_n27190_, new_n27191_, new_n27192_,
    new_n27193_, new_n27194_, new_n27195_, new_n27196_, new_n27197_,
    new_n27198_, new_n27199_, new_n27200_, new_n27201_, new_n27202_,
    new_n27203_, new_n27204_, new_n27205_, new_n27206_, new_n27207_,
    new_n27208_, new_n27209_, new_n27210_, new_n27211_, new_n27212_,
    new_n27213_, new_n27214_, new_n27215_, new_n27216_, new_n27217_,
    new_n27218_, new_n27219_, new_n27220_, new_n27221_, new_n27222_,
    new_n27223_, new_n27224_, new_n27225_, new_n27226_, new_n27227_,
    new_n27228_, new_n27229_, new_n27230_, new_n27231_, new_n27232_,
    new_n27233_, new_n27234_, new_n27236_, new_n27237_, new_n27238_,
    new_n27239_, new_n27240_, new_n27241_, new_n27242_, new_n27243_,
    new_n27244_, new_n27245_, new_n27246_, new_n27247_, new_n27248_,
    new_n27249_, new_n27250_, new_n27251_, new_n27252_, new_n27253_,
    new_n27254_, new_n27255_, new_n27256_, new_n27257_, new_n27258_,
    new_n27259_, new_n27260_, new_n27261_, new_n27262_, new_n27263_,
    new_n27264_, new_n27265_, new_n27266_, new_n27267_, new_n27268_,
    new_n27269_, new_n27270_, new_n27271_, new_n27272_, new_n27273_,
    new_n27274_, new_n27275_, new_n27276_, new_n27277_, new_n27278_,
    new_n27279_, new_n27280_, new_n27281_, new_n27282_, new_n27283_,
    new_n27284_, new_n27285_, new_n27286_, new_n27287_, new_n27288_,
    new_n27289_, new_n27290_, new_n27291_, new_n27292_, new_n27293_,
    new_n27294_, new_n27295_, new_n27296_, new_n27297_, new_n27298_,
    new_n27299_, new_n27300_, new_n27301_, new_n27302_, new_n27303_,
    new_n27304_, new_n27305_, new_n27306_, new_n27307_, new_n27308_,
    new_n27309_, new_n27310_, new_n27311_, new_n27312_, new_n27313_,
    new_n27314_, new_n27315_, new_n27316_, new_n27317_, new_n27318_,
    new_n27319_, new_n27320_, new_n27321_, new_n27322_, new_n27323_,
    new_n27324_, new_n27325_, new_n27326_, new_n27327_, new_n27328_,
    new_n27329_, new_n27330_, new_n27331_, new_n27332_, new_n27333_,
    new_n27334_, new_n27335_, new_n27336_, new_n27337_, new_n27338_,
    new_n27339_, new_n27340_, new_n27341_, new_n27342_, new_n27343_,
    new_n27344_, new_n27345_, new_n27346_, new_n27347_, new_n27348_,
    new_n27349_, new_n27350_, new_n27351_, new_n27352_, new_n27353_,
    new_n27354_, new_n27355_, new_n27356_, new_n27357_, new_n27358_,
    new_n27359_, new_n27360_, new_n27361_, new_n27362_, new_n27363_,
    new_n27364_, new_n27365_, new_n27366_, new_n27367_, new_n27368_,
    new_n27369_, new_n27370_, new_n27371_, new_n27372_, new_n27373_,
    new_n27374_, new_n27375_, new_n27376_, new_n27377_, new_n27378_,
    new_n27379_, new_n27380_, new_n27381_, new_n27382_, new_n27383_,
    new_n27384_, new_n27385_, new_n27386_, new_n27387_, new_n27388_,
    new_n27389_, new_n27390_, new_n27391_, new_n27392_, new_n27393_,
    new_n27394_, new_n27395_, new_n27396_, new_n27397_, new_n27398_,
    new_n27399_, new_n27400_, new_n27401_, new_n27402_, new_n27403_,
    new_n27404_, new_n27405_, new_n27406_, new_n27407_, new_n27408_,
    new_n27409_, new_n27410_, new_n27411_, new_n27412_, new_n27413_,
    new_n27414_, new_n27415_, new_n27416_, new_n27417_, new_n27418_,
    new_n27419_, new_n27420_, new_n27421_, new_n27422_, new_n27423_,
    new_n27424_, new_n27425_, new_n27426_, new_n27427_, new_n27428_,
    new_n27429_, new_n27430_, new_n27431_, new_n27432_, new_n27433_,
    new_n27434_, new_n27435_, new_n27436_, new_n27437_, new_n27438_,
    new_n27439_, new_n27440_, new_n27441_, new_n27442_, new_n27443_,
    new_n27444_, new_n27445_, new_n27446_, new_n27447_, new_n27448_,
    new_n27449_, new_n27450_, new_n27451_, new_n27452_, new_n27453_,
    new_n27454_, new_n27455_, new_n27456_, new_n27457_, new_n27458_,
    new_n27459_, new_n27460_, new_n27461_, new_n27462_, new_n27463_,
    new_n27464_, new_n27465_, new_n27466_, new_n27467_, new_n27468_,
    new_n27469_, new_n27470_, new_n27471_, new_n27472_, new_n27473_,
    new_n27474_, new_n27475_, new_n27476_, new_n27477_, new_n27478_,
    new_n27479_, new_n27480_, new_n27481_, new_n27482_, new_n27483_,
    new_n27484_, new_n27485_, new_n27486_, new_n27487_, new_n27488_,
    new_n27489_, new_n27490_, new_n27491_, new_n27492_, new_n27493_,
    new_n27494_, new_n27495_, new_n27496_, new_n27497_, new_n27498_,
    new_n27499_, new_n27500_, new_n27501_, new_n27502_, new_n27503_,
    new_n27504_, new_n27505_, new_n27506_, new_n27507_, new_n27508_,
    new_n27509_, new_n27510_, new_n27511_, new_n27512_, new_n27513_,
    new_n27514_, new_n27515_, new_n27516_, new_n27517_, new_n27518_,
    new_n27519_, new_n27520_, new_n27521_, new_n27522_, new_n27523_,
    new_n27524_, new_n27525_, new_n27526_, new_n27527_, new_n27528_,
    new_n27529_, new_n27530_, new_n27531_, new_n27532_, new_n27533_,
    new_n27534_, new_n27535_, new_n27536_, new_n27537_, new_n27538_,
    new_n27539_, new_n27540_, new_n27541_, new_n27542_, new_n27543_,
    new_n27544_, new_n27545_, new_n27546_, new_n27547_, new_n27548_,
    new_n27549_, new_n27550_, new_n27551_, new_n27552_, new_n27553_,
    new_n27554_, new_n27555_, new_n27556_, new_n27557_, new_n27558_,
    new_n27559_, new_n27560_, new_n27561_, new_n27562_, new_n27563_,
    new_n27564_, new_n27565_, new_n27566_, new_n27567_, new_n27568_,
    new_n27569_, new_n27570_, new_n27571_, new_n27572_, new_n27573_,
    new_n27574_, new_n27575_, new_n27576_, new_n27577_, new_n27578_,
    new_n27579_, new_n27580_, new_n27581_, new_n27582_, new_n27583_,
    new_n27584_, new_n27585_, new_n27586_, new_n27587_, new_n27588_,
    new_n27589_, new_n27590_, new_n27591_, new_n27592_, new_n27593_,
    new_n27594_, new_n27595_, new_n27596_, new_n27597_, new_n27598_,
    new_n27599_, new_n27600_, new_n27601_, new_n27602_, new_n27603_,
    new_n27604_, new_n27605_, new_n27606_, new_n27607_, new_n27608_,
    new_n27609_, new_n27610_, new_n27611_, new_n27612_, new_n27613_,
    new_n27614_, new_n27615_, new_n27616_, new_n27617_, new_n27618_,
    new_n27619_, new_n27620_, new_n27621_, new_n27622_, new_n27623_,
    new_n27624_, new_n27625_, new_n27626_, new_n27627_, new_n27628_,
    new_n27629_, new_n27630_, new_n27631_, new_n27632_, new_n27633_,
    new_n27634_, new_n27635_, new_n27636_, new_n27637_, new_n27638_,
    new_n27639_, new_n27640_, new_n27641_, new_n27642_, new_n27643_,
    new_n27644_, new_n27645_, new_n27646_, new_n27647_, new_n27648_,
    new_n27649_, new_n27650_, new_n27651_, new_n27652_, new_n27653_,
    new_n27654_, new_n27655_, new_n27656_, new_n27657_, new_n27658_,
    new_n27659_, new_n27660_, new_n27661_, new_n27662_, new_n27663_,
    new_n27664_, new_n27665_, new_n27666_, new_n27667_, new_n27668_,
    new_n27669_, new_n27670_, new_n27671_, new_n27672_, new_n27673_,
    new_n27674_, new_n27675_, new_n27676_, new_n27677_, new_n27678_,
    new_n27679_, new_n27680_, new_n27681_, new_n27682_, new_n27683_,
    new_n27684_, new_n27685_, new_n27686_, new_n27687_, new_n27688_,
    new_n27689_, new_n27690_, new_n27691_, new_n27692_, new_n27693_,
    new_n27694_, new_n27695_, new_n27696_, new_n27697_, new_n27698_,
    new_n27699_, new_n27700_, new_n27701_, new_n27702_, new_n27703_,
    new_n27704_, new_n27705_, new_n27706_, new_n27707_, new_n27708_,
    new_n27709_, new_n27710_, new_n27711_, new_n27712_, new_n27713_,
    new_n27714_, new_n27715_, new_n27716_, new_n27717_, new_n27718_,
    new_n27719_, new_n27720_, new_n27721_, new_n27722_, new_n27723_,
    new_n27724_, new_n27725_, new_n27726_, new_n27727_, new_n27728_,
    new_n27729_, new_n27730_, new_n27731_, new_n27732_, new_n27733_,
    new_n27734_, new_n27735_, new_n27736_, new_n27737_, new_n27738_,
    new_n27739_, new_n27740_, new_n27741_, new_n27742_, new_n27743_,
    new_n27744_, new_n27745_, new_n27746_, new_n27747_, new_n27748_,
    new_n27749_, new_n27750_, new_n27751_, new_n27752_, new_n27753_,
    new_n27754_, new_n27755_, new_n27756_, new_n27757_, new_n27758_,
    new_n27759_, new_n27760_, new_n27761_, new_n27762_, new_n27763_,
    new_n27764_, new_n27765_, new_n27766_, new_n27767_, new_n27768_,
    new_n27769_, new_n27770_, new_n27771_, new_n27772_, new_n27773_,
    new_n27774_, new_n27775_, new_n27776_, new_n27777_, new_n27778_,
    new_n27779_, new_n27780_, new_n27781_, new_n27782_, new_n27783_,
    new_n27784_, new_n27785_, new_n27786_, new_n27787_, new_n27788_,
    new_n27789_, new_n27790_, new_n27791_, new_n27792_, new_n27793_,
    new_n27794_, new_n27795_, new_n27796_, new_n27797_, new_n27798_,
    new_n27799_, new_n27800_, new_n27801_, new_n27802_, new_n27803_,
    new_n27804_, new_n27805_, new_n27806_, new_n27807_, new_n27808_,
    new_n27809_, new_n27810_, new_n27811_, new_n27812_, new_n27813_,
    new_n27814_, new_n27815_, new_n27816_, new_n27817_, new_n27818_,
    new_n27819_, new_n27820_, new_n27821_, new_n27822_, new_n27823_,
    new_n27824_, new_n27825_, new_n27826_, new_n27827_, new_n27828_,
    new_n27829_, new_n27830_, new_n27831_, new_n27832_, new_n27833_,
    new_n27834_, new_n27835_, new_n27836_, new_n27837_, new_n27838_,
    new_n27839_, new_n27840_, new_n27841_, new_n27842_, new_n27843_,
    new_n27844_, new_n27845_, new_n27846_, new_n27847_, new_n27848_,
    new_n27849_, new_n27850_, new_n27851_, new_n27852_, new_n27853_,
    new_n27854_, new_n27855_, new_n27856_, new_n27857_, new_n27858_,
    new_n27859_, new_n27860_, new_n27861_, new_n27862_, new_n27863_,
    new_n27864_, new_n27865_, new_n27866_, new_n27867_, new_n27868_,
    new_n27869_, new_n27870_, new_n27871_, new_n27872_, new_n27873_,
    new_n27874_, new_n27875_, new_n27876_, new_n27877_, new_n27878_,
    new_n27879_, new_n27880_, new_n27881_, new_n27882_, new_n27883_,
    new_n27884_, new_n27885_, new_n27886_, new_n27887_, new_n27888_,
    new_n27889_, new_n27890_, new_n27891_, new_n27892_, new_n27893_,
    new_n27894_, new_n27895_, new_n27896_, new_n27897_, new_n27898_,
    new_n27899_, new_n27900_, new_n27901_, new_n27902_, new_n27903_,
    new_n27904_, new_n27905_, new_n27906_, new_n27907_, new_n27908_,
    new_n27909_, new_n27910_, new_n27911_, new_n27912_, new_n27913_,
    new_n27914_, new_n27915_, new_n27916_, new_n27917_, new_n27918_,
    new_n27919_, new_n27920_, new_n27921_, new_n27922_, new_n27923_,
    new_n27924_, new_n27925_, new_n27926_, new_n27927_, new_n27928_,
    new_n27929_, new_n27930_, new_n27931_, new_n27932_, new_n27933_,
    new_n27934_, new_n27935_, new_n27936_, new_n27937_, new_n27938_,
    new_n27939_, new_n27940_, new_n27941_, new_n27942_, new_n27943_,
    new_n27944_, new_n27945_, new_n27946_, new_n27947_, new_n27948_,
    new_n27949_, new_n27950_, new_n27951_, new_n27952_, new_n27953_,
    new_n27954_, new_n27955_, new_n27956_, new_n27957_, new_n27958_,
    new_n27959_, new_n27960_, new_n27961_, new_n27962_, new_n27963_,
    new_n27964_, new_n27965_, new_n27966_, new_n27967_, new_n27968_,
    new_n27969_, new_n27970_, new_n27971_, new_n27972_, new_n27973_,
    new_n27974_, new_n27975_, new_n27976_, new_n27977_, new_n27978_,
    new_n27979_, new_n27980_, new_n27981_, new_n27982_, new_n27983_,
    new_n27984_, new_n27985_, new_n27986_, new_n27987_, new_n27988_,
    new_n27989_, new_n27990_, new_n27991_, new_n27992_, new_n27993_,
    new_n27994_, new_n27995_, new_n27996_, new_n27997_, new_n27998_,
    new_n27999_, new_n28000_, new_n28001_, new_n28002_, new_n28003_,
    new_n28004_, new_n28005_, new_n28006_, new_n28007_, new_n28008_,
    new_n28009_, new_n28010_, new_n28011_, new_n28012_, new_n28013_,
    new_n28014_, new_n28015_, new_n28016_, new_n28017_, new_n28018_,
    new_n28019_, new_n28020_, new_n28021_, new_n28022_, new_n28023_,
    new_n28024_, new_n28025_, new_n28026_, new_n28027_, new_n28028_,
    new_n28029_, new_n28030_, new_n28031_, new_n28032_, new_n28033_,
    new_n28034_, new_n28035_, new_n28036_, new_n28037_, new_n28038_,
    new_n28039_, new_n28040_, new_n28041_, new_n28042_, new_n28043_,
    new_n28044_, new_n28045_, new_n28046_, new_n28047_, new_n28048_,
    new_n28049_, new_n28050_, new_n28051_, new_n28052_, new_n28053_,
    new_n28054_, new_n28055_, new_n28056_, new_n28057_, new_n28058_,
    new_n28059_, new_n28060_, new_n28061_, new_n28062_, new_n28063_,
    new_n28064_, new_n28065_, new_n28066_, new_n28067_, new_n28068_,
    new_n28069_, new_n28070_, new_n28071_, new_n28072_, new_n28073_,
    new_n28074_, new_n28075_, new_n28076_, new_n28077_, new_n28078_,
    new_n28079_, new_n28080_, new_n28081_, new_n28082_, new_n28083_,
    new_n28084_, new_n28085_, new_n28086_, new_n28087_, new_n28088_,
    new_n28089_, new_n28090_, new_n28091_, new_n28092_, new_n28093_,
    new_n28094_, new_n28095_, new_n28096_, new_n28097_, new_n28098_,
    new_n28099_, new_n28100_, new_n28101_, new_n28102_, new_n28103_,
    new_n28105_, new_n28106_, new_n28107_, new_n28108_, new_n28109_,
    new_n28110_, new_n28111_, new_n28112_, new_n28113_, new_n28114_,
    new_n28115_, new_n28116_, new_n28117_, new_n28118_, new_n28119_,
    new_n28120_, new_n28121_, new_n28122_, new_n28123_, new_n28124_,
    new_n28125_, new_n28126_, new_n28127_, new_n28128_, new_n28129_,
    new_n28130_, new_n28131_, new_n28132_, new_n28133_, new_n28134_,
    new_n28135_, new_n28136_, new_n28137_, new_n28138_, new_n28139_,
    new_n28140_, new_n28141_, new_n28142_, new_n28143_, new_n28144_,
    new_n28145_, new_n28146_, new_n28147_, new_n28148_, new_n28149_,
    new_n28150_, new_n28151_, new_n28152_, new_n28153_, new_n28154_,
    new_n28155_, new_n28156_, new_n28157_, new_n28158_, new_n28159_,
    new_n28160_, new_n28161_, new_n28162_, new_n28163_, new_n28164_,
    new_n28165_, new_n28166_, new_n28167_, new_n28168_, new_n28169_,
    new_n28170_, new_n28171_, new_n28172_, new_n28173_, new_n28174_,
    new_n28175_, new_n28176_, new_n28177_, new_n28178_, new_n28179_,
    new_n28180_, new_n28181_, new_n28182_, new_n28183_, new_n28184_,
    new_n28185_, new_n28186_, new_n28187_, new_n28188_, new_n28189_,
    new_n28190_, new_n28191_, new_n28192_, new_n28193_, new_n28194_,
    new_n28195_, new_n28196_, new_n28197_, new_n28198_, new_n28199_,
    new_n28200_, new_n28201_, new_n28202_, new_n28203_, new_n28204_,
    new_n28205_, new_n28206_, new_n28207_, new_n28208_, new_n28209_,
    new_n28210_, new_n28211_, new_n28212_, new_n28213_, new_n28214_,
    new_n28215_, new_n28216_, new_n28217_, new_n28218_, new_n28219_,
    new_n28220_, new_n28221_, new_n28222_, new_n28223_, new_n28224_,
    new_n28225_, new_n28226_, new_n28227_, new_n28228_, new_n28229_,
    new_n28230_, new_n28231_, new_n28232_, new_n28233_, new_n28234_,
    new_n28235_, new_n28236_, new_n28237_, new_n28238_, new_n28239_,
    new_n28240_, new_n28241_, new_n28242_, new_n28243_, new_n28244_,
    new_n28245_, new_n28246_, new_n28247_, new_n28248_, new_n28249_,
    new_n28250_, new_n28251_, new_n28252_, new_n28253_, new_n28254_,
    new_n28255_, new_n28256_, new_n28257_, new_n28258_, new_n28259_,
    new_n28260_, new_n28261_, new_n28262_, new_n28263_, new_n28264_,
    new_n28265_, new_n28266_, new_n28267_, new_n28268_, new_n28269_,
    new_n28270_, new_n28271_, new_n28272_, new_n28273_, new_n28274_,
    new_n28275_, new_n28276_, new_n28277_, new_n28278_, new_n28279_,
    new_n28280_, new_n28281_, new_n28282_, new_n28283_, new_n28284_,
    new_n28285_, new_n28286_, new_n28287_, new_n28288_, new_n28289_,
    new_n28290_, new_n28291_, new_n28292_, new_n28293_, new_n28294_,
    new_n28295_, new_n28296_, new_n28297_, new_n28298_, new_n28299_,
    new_n28300_, new_n28301_, new_n28302_, new_n28303_, new_n28304_,
    new_n28305_, new_n28306_, new_n28307_, new_n28308_, new_n28309_,
    new_n28310_, new_n28311_, new_n28312_, new_n28313_, new_n28314_,
    new_n28315_, new_n28316_, new_n28317_, new_n28318_, new_n28319_,
    new_n28320_, new_n28321_, new_n28322_, new_n28323_, new_n28324_,
    new_n28325_, new_n28326_, new_n28327_, new_n28328_, new_n28329_,
    new_n28330_, new_n28331_, new_n28332_, new_n28333_, new_n28334_,
    new_n28335_, new_n28336_, new_n28337_, new_n28338_, new_n28339_,
    new_n28340_, new_n28341_, new_n28342_, new_n28343_, new_n28344_,
    new_n28345_, new_n28346_, new_n28347_, new_n28348_, new_n28349_,
    new_n28350_, new_n28351_, new_n28352_, new_n28353_, new_n28354_,
    new_n28355_, new_n28356_, new_n28357_, new_n28358_, new_n28359_,
    new_n28360_, new_n28361_, new_n28362_, new_n28363_, new_n28364_,
    new_n28365_, new_n28366_, new_n28367_, new_n28368_, new_n28369_,
    new_n28370_, new_n28371_, new_n28372_, new_n28373_, new_n28374_,
    new_n28375_, new_n28376_, new_n28377_, new_n28378_, new_n28379_,
    new_n28380_, new_n28381_, new_n28382_, new_n28383_, new_n28384_,
    new_n28385_, new_n28386_, new_n28387_, new_n28388_, new_n28389_,
    new_n28390_, new_n28391_, new_n28392_, new_n28393_, new_n28394_,
    new_n28395_, new_n28396_, new_n28397_, new_n28398_, new_n28399_,
    new_n28400_, new_n28401_, new_n28402_, new_n28403_, new_n28404_,
    new_n28405_, new_n28406_, new_n28407_, new_n28408_, new_n28409_,
    new_n28410_, new_n28411_, new_n28412_, new_n28413_, new_n28414_,
    new_n28415_, new_n28416_, new_n28417_, new_n28418_, new_n28419_,
    new_n28420_, new_n28421_, new_n28422_, new_n28423_, new_n28424_,
    new_n28425_, new_n28426_, new_n28427_, new_n28428_, new_n28429_,
    new_n28430_, new_n28431_, new_n28432_, new_n28433_, new_n28434_,
    new_n28435_, new_n28436_, new_n28437_, new_n28438_, new_n28439_,
    new_n28440_, new_n28441_, new_n28442_, new_n28443_, new_n28444_,
    new_n28445_, new_n28446_, new_n28447_, new_n28448_, new_n28449_,
    new_n28450_, new_n28451_, new_n28452_, new_n28453_, new_n28454_,
    new_n28455_, new_n28456_, new_n28457_, new_n28458_, new_n28459_,
    new_n28460_, new_n28461_, new_n28462_, new_n28463_, new_n28464_,
    new_n28465_, new_n28466_, new_n28467_, new_n28468_, new_n28469_,
    new_n28470_, new_n28471_, new_n28472_, new_n28473_, new_n28474_,
    new_n28475_, new_n28476_, new_n28477_, new_n28478_, new_n28479_,
    new_n28480_, new_n28481_, new_n28482_, new_n28483_, new_n28484_,
    new_n28485_, new_n28486_, new_n28487_, new_n28488_, new_n28489_,
    new_n28490_, new_n28491_, new_n28492_, new_n28493_, new_n28494_,
    new_n28495_, new_n28496_, new_n28497_, new_n28498_, new_n28499_,
    new_n28500_, new_n28501_, new_n28502_, new_n28503_, new_n28504_,
    new_n28505_, new_n28506_, new_n28507_, new_n28508_, new_n28509_,
    new_n28510_, new_n28511_, new_n28512_, new_n28513_, new_n28514_,
    new_n28515_, new_n28516_, new_n28517_, new_n28518_, new_n28519_,
    new_n28520_, new_n28521_, new_n28522_, new_n28523_, new_n28524_,
    new_n28525_, new_n28526_, new_n28527_, new_n28528_, new_n28529_,
    new_n28530_, new_n28531_, new_n28532_, new_n28533_, new_n28534_,
    new_n28535_, new_n28536_, new_n28537_, new_n28538_, new_n28539_,
    new_n28540_, new_n28541_, new_n28542_, new_n28543_, new_n28544_,
    new_n28545_, new_n28546_, new_n28547_, new_n28548_, new_n28549_,
    new_n28550_, new_n28551_, new_n28552_, new_n28553_, new_n28554_,
    new_n28555_, new_n28556_, new_n28557_, new_n28558_, new_n28559_,
    new_n28560_, new_n28561_, new_n28562_, new_n28563_, new_n28564_,
    new_n28565_, new_n28566_, new_n28567_, new_n28568_, new_n28569_,
    new_n28570_, new_n28571_, new_n28572_, new_n28573_, new_n28574_,
    new_n28575_, new_n28576_, new_n28577_, new_n28578_, new_n28579_,
    new_n28580_, new_n28581_, new_n28582_, new_n28583_, new_n28584_,
    new_n28585_, new_n28586_, new_n28587_, new_n28588_, new_n28589_,
    new_n28590_, new_n28591_, new_n28592_, new_n28593_, new_n28594_,
    new_n28595_, new_n28596_, new_n28597_, new_n28598_, new_n28599_,
    new_n28600_, new_n28601_, new_n28602_, new_n28603_, new_n28604_,
    new_n28605_, new_n28606_, new_n28607_, new_n28608_, new_n28609_,
    new_n28610_, new_n28611_, new_n28612_, new_n28613_, new_n28614_,
    new_n28615_, new_n28616_, new_n28617_, new_n28618_, new_n28619_,
    new_n28620_, new_n28621_, new_n28622_, new_n28623_, new_n28624_,
    new_n28625_, new_n28626_, new_n28627_, new_n28628_, new_n28629_,
    new_n28630_, new_n28631_, new_n28632_, new_n28633_, new_n28634_,
    new_n28635_, new_n28636_, new_n28637_, new_n28638_, new_n28639_,
    new_n28640_, new_n28641_, new_n28642_, new_n28643_, new_n28644_,
    new_n28645_, new_n28646_, new_n28647_, new_n28648_, new_n28649_,
    new_n28650_, new_n28651_, new_n28652_, new_n28653_, new_n28654_,
    new_n28655_, new_n28656_, new_n28657_, new_n28658_, new_n28659_,
    new_n28660_, new_n28661_, new_n28662_, new_n28663_, new_n28664_,
    new_n28665_, new_n28666_, new_n28667_, new_n28668_, new_n28669_,
    new_n28670_, new_n28671_, new_n28672_, new_n28673_, new_n28674_,
    new_n28675_, new_n28676_, new_n28677_, new_n28678_, new_n28679_,
    new_n28680_, new_n28681_, new_n28682_, new_n28683_, new_n28684_,
    new_n28685_, new_n28686_, new_n28687_, new_n28688_, new_n28689_,
    new_n28690_, new_n28691_, new_n28692_, new_n28693_, new_n28694_,
    new_n28695_, new_n28696_, new_n28697_, new_n28698_, new_n28699_,
    new_n28700_, new_n28701_, new_n28702_, new_n28703_, new_n28704_,
    new_n28705_, new_n28706_, new_n28707_, new_n28708_, new_n28709_,
    new_n28710_, new_n28711_, new_n28712_, new_n28713_, new_n28714_,
    new_n28715_, new_n28716_, new_n28717_, new_n28718_, new_n28719_,
    new_n28720_, new_n28721_, new_n28722_, new_n28723_, new_n28724_,
    new_n28725_, new_n28726_, new_n28727_, new_n28728_, new_n28729_,
    new_n28730_, new_n28731_, new_n28732_, new_n28733_, new_n28734_,
    new_n28735_, new_n28736_, new_n28737_, new_n28738_, new_n28739_,
    new_n28740_, new_n28741_, new_n28742_, new_n28743_, new_n28744_,
    new_n28745_, new_n28746_, new_n28747_, new_n28748_, new_n28749_,
    new_n28750_, new_n28751_, new_n28752_, new_n28753_, new_n28754_,
    new_n28755_, new_n28756_, new_n28757_, new_n28758_, new_n28759_,
    new_n28760_, new_n28761_, new_n28762_, new_n28763_, new_n28764_,
    new_n28765_, new_n28766_, new_n28767_, new_n28768_, new_n28769_,
    new_n28770_, new_n28771_, new_n28772_, new_n28773_, new_n28774_,
    new_n28775_, new_n28776_, new_n28777_, new_n28778_, new_n28779_,
    new_n28780_, new_n28781_, new_n28782_, new_n28783_, new_n28784_,
    new_n28785_, new_n28786_, new_n28787_, new_n28788_, new_n28789_,
    new_n28790_, new_n28791_, new_n28792_, new_n28793_, new_n28794_,
    new_n28795_, new_n28796_, new_n28797_, new_n28798_, new_n28799_,
    new_n28800_, new_n28801_, new_n28802_, new_n28803_, new_n28804_,
    new_n28805_, new_n28806_, new_n28807_, new_n28808_, new_n28809_,
    new_n28810_, new_n28811_, new_n28812_, new_n28813_, new_n28814_,
    new_n28815_, new_n28816_, new_n28817_, new_n28818_, new_n28819_,
    new_n28820_, new_n28821_, new_n28822_, new_n28823_, new_n28824_,
    new_n28825_, new_n28826_, new_n28827_, new_n28828_, new_n28829_,
    new_n28830_, new_n28831_, new_n28832_, new_n28833_, new_n28834_,
    new_n28835_, new_n28836_, new_n28837_, new_n28838_, new_n28839_,
    new_n28840_, new_n28841_, new_n28842_, new_n28843_, new_n28844_,
    new_n28845_, new_n28846_, new_n28847_, new_n28848_, new_n28849_,
    new_n28850_, new_n28851_, new_n28852_, new_n28853_, new_n28854_,
    new_n28855_, new_n28856_, new_n28857_, new_n28858_, new_n28859_,
    new_n28860_, new_n28861_, new_n28862_, new_n28863_, new_n28864_,
    new_n28865_, new_n28866_, new_n28867_, new_n28868_, new_n28869_,
    new_n28870_, new_n28871_, new_n28872_, new_n28873_, new_n28874_,
    new_n28875_, new_n28876_, new_n28877_, new_n28878_, new_n28879_,
    new_n28880_, new_n28881_, new_n28882_, new_n28883_, new_n28884_,
    new_n28885_, new_n28886_, new_n28887_, new_n28888_, new_n28889_,
    new_n28890_, new_n28891_, new_n28892_, new_n28893_, new_n28894_,
    new_n28895_, new_n28896_, new_n28897_, new_n28898_, new_n28899_,
    new_n28900_, new_n28901_, new_n28902_, new_n28903_, new_n28904_,
    new_n28905_, new_n28906_, new_n28907_, new_n28908_, new_n28909_,
    new_n28910_, new_n28911_, new_n28912_, new_n28913_, new_n28914_,
    new_n28915_, new_n28916_, new_n28917_, new_n28918_, new_n28919_,
    new_n28920_, new_n28923_, new_n28924_, new_n28926_, new_n28927_,
    new_n28928_, new_n28929_, new_n28931_, new_n28932_, new_n28933_,
    new_n28934_, new_n28935_, new_n28936_, new_n28937_, new_n28938_,
    new_n28939_, new_n28940_, new_n28941_, new_n28942_, new_n28943_,
    new_n28944_, new_n28945_, new_n28946_, new_n28947_, new_n28948_,
    new_n28949_, new_n28950_, new_n28951_, new_n28952_, new_n28953_,
    new_n28954_, new_n28955_, new_n28956_, new_n28957_, new_n28958_,
    new_n28959_, new_n28960_, new_n28961_, new_n28962_, new_n28963_,
    new_n28964_, new_n28965_, new_n28966_, new_n28967_, new_n28968_,
    new_n28969_, new_n28970_, new_n28971_, new_n28972_, new_n28973_,
    new_n28974_, new_n28975_, new_n28976_, new_n28977_, new_n28978_,
    new_n28979_, new_n28980_, new_n28981_, new_n28982_, new_n28983_,
    new_n28984_, new_n28985_, new_n28986_, new_n28987_, new_n28988_,
    new_n28989_, new_n28990_, new_n28991_, new_n28992_, new_n28993_,
    new_n28994_, new_n28995_, new_n28996_, new_n28997_, new_n28998_,
    new_n28999_, new_n29000_, new_n29001_, new_n29002_, new_n29003_,
    new_n29004_, new_n29005_, new_n29006_, new_n29007_, new_n29008_,
    new_n29009_, new_n29010_, new_n29011_, new_n29012_, new_n29013_,
    new_n29014_, new_n29015_, new_n29016_, new_n29017_, new_n29018_,
    new_n29019_, new_n29020_, new_n29021_, new_n29022_, new_n29023_,
    new_n29024_, new_n29025_, new_n29026_, new_n29027_, new_n29028_,
    new_n29029_, new_n29030_, new_n29031_, new_n29032_, new_n29033_,
    new_n29034_, new_n29035_, new_n29036_, new_n29037_, new_n29038_,
    new_n29039_, new_n29040_, new_n29041_, new_n29042_, new_n29043_,
    new_n29044_, new_n29045_, new_n29046_, new_n29047_, new_n29048_,
    new_n29049_, new_n29050_, new_n29051_, new_n29052_, new_n29053_,
    new_n29054_, new_n29055_, new_n29056_, new_n29057_, new_n29058_,
    new_n29059_, new_n29060_, new_n29061_, new_n29062_, new_n29063_,
    new_n29064_, new_n29065_, new_n29066_, new_n29067_, new_n29068_,
    new_n29069_, new_n29070_, new_n29071_, new_n29072_, new_n29073_,
    new_n29074_, new_n29075_, new_n29076_, new_n29077_, new_n29078_,
    new_n29079_, new_n29080_, new_n29081_, new_n29082_, new_n29083_,
    new_n29084_, new_n29085_, new_n29086_, new_n29087_, new_n29088_,
    new_n29089_, new_n29090_, new_n29091_, new_n29092_, new_n29093_,
    new_n29094_, new_n29095_, new_n29096_, new_n29097_, new_n29098_,
    new_n29099_, new_n29100_, new_n29101_, new_n29102_, new_n29103_,
    new_n29104_, new_n29105_, new_n29106_, new_n29107_, new_n29108_,
    new_n29109_, new_n29110_, new_n29111_, new_n29112_, new_n29113_,
    new_n29114_, new_n29115_, new_n29116_, new_n29117_, new_n29118_,
    new_n29119_, new_n29120_, new_n29121_, new_n29122_, new_n29123_,
    new_n29124_, new_n29125_, new_n29126_, new_n29127_, new_n29128_,
    new_n29129_, new_n29130_, new_n29131_, new_n29132_, new_n29133_,
    new_n29134_, new_n29135_, new_n29136_, new_n29137_, new_n29138_,
    new_n29139_, new_n29140_, new_n29141_, new_n29142_, new_n29143_,
    new_n29144_, new_n29145_, new_n29146_, new_n29147_, new_n29148_,
    new_n29149_, new_n29150_, new_n29151_, new_n29152_, new_n29153_,
    new_n29154_, new_n29155_, new_n29156_, new_n29157_, new_n29158_,
    new_n29159_, new_n29160_, new_n29161_, new_n29162_, new_n29163_,
    new_n29164_, new_n29165_, new_n29166_, new_n29167_, new_n29168_,
    new_n29169_, new_n29170_, new_n29171_, new_n29172_, new_n29173_,
    new_n29174_, new_n29175_, new_n29176_, new_n29177_, new_n29178_,
    new_n29179_, new_n29180_, new_n29181_, new_n29182_, new_n29183_,
    new_n29184_, new_n29185_, new_n29186_, new_n29187_, new_n29188_,
    new_n29189_, new_n29190_, new_n29191_, new_n29192_, new_n29193_,
    new_n29194_, new_n29195_, new_n29196_, new_n29197_, new_n29198_,
    new_n29199_, new_n29200_, new_n29201_, new_n29202_, new_n29203_,
    new_n29204_, new_n29205_, new_n29206_, new_n29207_, new_n29208_,
    new_n29209_, new_n29210_, new_n29211_, new_n29212_, new_n29213_,
    new_n29214_, new_n29215_, new_n29216_, new_n29217_, new_n29218_,
    new_n29219_, new_n29220_, new_n29221_, new_n29222_, new_n29223_,
    new_n29224_, new_n29225_, new_n29226_, new_n29227_, new_n29228_,
    new_n29229_, new_n29230_, new_n29231_, new_n29232_, new_n29233_,
    new_n29234_, new_n29235_, new_n29236_, new_n29237_, new_n29238_,
    new_n29239_, new_n29240_, new_n29241_, new_n29242_, new_n29243_,
    new_n29244_, new_n29245_, new_n29246_, new_n29247_, new_n29248_,
    new_n29249_, new_n29250_, new_n29251_, new_n29252_, new_n29253_,
    new_n29254_, new_n29255_, new_n29256_, new_n29257_, new_n29258_,
    new_n29259_, new_n29260_, new_n29261_, new_n29262_, new_n29263_,
    new_n29264_, new_n29265_, new_n29266_, new_n29267_, new_n29268_,
    new_n29269_, new_n29270_, new_n29271_, new_n29272_, new_n29273_,
    new_n29274_, new_n29275_, new_n29276_, new_n29277_, new_n29278_,
    new_n29279_, new_n29280_, new_n29281_, new_n29282_, new_n29283_,
    new_n29284_, new_n29285_, new_n29286_, new_n29287_, new_n29288_,
    new_n29289_, new_n29290_, new_n29291_, new_n29292_, new_n29293_,
    new_n29294_, new_n29295_, new_n29296_, new_n29297_, new_n29298_,
    new_n29299_, new_n29300_, new_n29301_, new_n29302_, new_n29303_,
    new_n29304_, new_n29305_, new_n29306_, new_n29307_, new_n29308_,
    new_n29309_, new_n29310_, new_n29311_, new_n29312_, new_n29313_,
    new_n29314_, new_n29315_, new_n29316_, new_n29317_, new_n29318_,
    new_n29319_, new_n29320_, new_n29321_, new_n29322_, new_n29323_,
    new_n29324_, new_n29325_, new_n29326_, new_n29327_, new_n29328_,
    new_n29329_, new_n29330_, new_n29331_, new_n29332_, new_n29333_,
    new_n29334_, new_n29335_, new_n29336_, new_n29337_, new_n29338_,
    new_n29339_, new_n29340_, new_n29341_, new_n29342_, new_n29343_,
    new_n29344_, new_n29345_, new_n29346_, new_n29347_, new_n29348_,
    new_n29349_, new_n29350_, new_n29351_, new_n29352_, new_n29353_,
    new_n29354_, new_n29355_, new_n29356_, new_n29357_, new_n29358_,
    new_n29359_, new_n29360_, new_n29361_, new_n29362_, new_n29363_,
    new_n29364_, new_n29365_, new_n29366_, new_n29367_, new_n29368_,
    new_n29369_, new_n29370_, new_n29371_, new_n29372_, new_n29373_,
    new_n29374_, new_n29375_, new_n29376_, new_n29377_, new_n29378_,
    new_n29379_, new_n29380_, new_n29381_, new_n29382_, new_n29383_,
    new_n29384_, new_n29385_, new_n29386_, new_n29387_, new_n29388_,
    new_n29389_, new_n29390_, new_n29391_, new_n29392_, new_n29393_,
    new_n29394_, new_n29395_, new_n29396_, new_n29397_, new_n29398_,
    new_n29399_, new_n29400_, new_n29401_, new_n29402_, new_n29403_,
    new_n29404_, new_n29405_, new_n29406_, new_n29407_, new_n29408_,
    new_n29409_, new_n29410_, new_n29411_, new_n29412_, new_n29413_,
    new_n29414_, new_n29415_, new_n29416_, new_n29417_, new_n29418_,
    new_n29419_, new_n29420_, new_n29421_, new_n29422_, new_n29423_,
    new_n29424_, new_n29425_, new_n29426_, new_n29427_, new_n29428_,
    new_n29429_, new_n29430_, new_n29431_, new_n29432_, new_n29433_,
    new_n29434_, new_n29435_, new_n29436_, new_n29437_, new_n29438_,
    new_n29439_, new_n29440_, new_n29441_, new_n29442_, new_n29443_,
    new_n29444_, new_n29445_, new_n29446_, new_n29447_, new_n29448_,
    new_n29449_, new_n29450_, new_n29451_, new_n29452_, new_n29453_,
    new_n29454_, new_n29455_, new_n29456_, new_n29457_, new_n29458_,
    new_n29459_, new_n29460_, new_n29461_, new_n29462_, new_n29463_,
    new_n29464_, new_n29465_, new_n29466_, new_n29467_, new_n29468_,
    new_n29469_, new_n29470_, new_n29471_, new_n29472_, new_n29473_,
    new_n29474_, new_n29475_, new_n29476_, new_n29477_, new_n29478_,
    new_n29479_, new_n29480_, new_n29481_, new_n29482_, new_n29483_,
    new_n29484_, new_n29485_, new_n29486_, new_n29487_, new_n29488_,
    new_n29489_, new_n29490_, new_n29491_, new_n29492_, new_n29493_,
    new_n29494_, new_n29495_, new_n29496_, new_n29497_, new_n29498_,
    new_n29499_, new_n29500_, new_n29501_, new_n29502_, new_n29503_,
    new_n29504_, new_n29505_, new_n29506_, new_n29507_, new_n29508_,
    new_n29509_, new_n29510_, new_n29511_, new_n29512_, new_n29513_,
    new_n29514_, new_n29515_, new_n29516_, new_n29517_, new_n29518_,
    new_n29519_, new_n29520_, new_n29521_, new_n29522_, new_n29523_,
    new_n29524_, new_n29525_, new_n29526_, new_n29527_, new_n29528_,
    new_n29529_, new_n29530_, new_n29531_, new_n29532_, new_n29533_,
    new_n29534_, new_n29535_, new_n29536_, new_n29537_, new_n29538_,
    new_n29539_, new_n29540_, new_n29541_, new_n29542_, new_n29543_,
    new_n29544_, new_n29545_, new_n29546_, new_n29547_, new_n29548_,
    new_n29549_, new_n29550_, new_n29551_, new_n29552_, new_n29553_,
    new_n29554_, new_n29555_, new_n29556_, new_n29557_, new_n29558_,
    new_n29559_, new_n29560_, new_n29561_, new_n29562_, new_n29563_,
    new_n29564_, new_n29565_, new_n29566_, new_n29567_, new_n29568_,
    new_n29569_, new_n29570_, new_n29571_, new_n29572_, new_n29573_,
    new_n29574_, new_n29575_, new_n29576_, new_n29577_, new_n29578_,
    new_n29579_, new_n29580_, new_n29581_, new_n29582_, new_n29583_,
    new_n29584_, new_n29585_, new_n29586_, new_n29587_, new_n29588_,
    new_n29589_, new_n29590_, new_n29591_, new_n29592_, new_n29593_,
    new_n29594_, new_n29595_, new_n29596_, new_n29597_, new_n29598_,
    new_n29599_, new_n29600_, new_n29601_, new_n29602_, new_n29603_,
    new_n29604_, new_n29605_, new_n29606_, new_n29607_, new_n29608_,
    new_n29609_, new_n29610_, new_n29611_, new_n29612_, new_n29613_,
    new_n29614_, new_n29615_, new_n29616_, new_n29617_, new_n29618_,
    new_n29619_, new_n29620_, new_n29621_, new_n29622_, new_n29623_,
    new_n29624_, new_n29625_, new_n29626_, new_n29627_, new_n29628_,
    new_n29629_, new_n29630_, new_n29631_, new_n29632_, new_n29633_,
    new_n29634_, new_n29635_, new_n29636_, new_n29637_, new_n29638_,
    new_n29639_, new_n29640_, new_n29641_, new_n29642_, new_n29643_,
    new_n29644_, new_n29645_, new_n29646_, new_n29647_, new_n29648_,
    new_n29649_, new_n29650_, new_n29651_, new_n29652_, new_n29653_,
    new_n29654_, new_n29655_, new_n29656_, new_n29657_, new_n29658_,
    new_n29659_, new_n29660_, new_n29661_, new_n29662_, new_n29663_,
    new_n29664_, new_n29665_, new_n29666_, new_n29667_, new_n29668_,
    new_n29669_, new_n29670_, new_n29671_, new_n29672_, new_n29673_,
    new_n29674_, new_n29675_, new_n29676_, new_n29677_, new_n29678_,
    new_n29679_, new_n29680_, new_n29681_, new_n29682_, new_n29683_,
    new_n29684_, new_n29685_, new_n29686_, new_n29687_, new_n29688_,
    new_n29689_, new_n29690_, new_n29691_, new_n29692_, new_n29693_,
    new_n29694_, new_n29695_, new_n29696_, new_n29697_, new_n29698_,
    new_n29699_, new_n29700_, new_n29701_, new_n29702_, new_n29703_,
    new_n29704_, new_n29705_, new_n29706_, new_n29707_, new_n29708_,
    new_n29709_, new_n29710_, new_n29711_, new_n29712_, new_n29713_,
    new_n29714_, new_n29715_, new_n29716_, new_n29717_, new_n29718_,
    new_n29719_, new_n29720_, new_n29721_, new_n29722_, new_n29723_,
    new_n29724_, new_n29725_, new_n29726_, new_n29727_, new_n29728_,
    new_n29729_, new_n29730_, new_n29731_, new_n29732_, new_n29733_,
    new_n29734_, new_n29735_, new_n29736_, new_n29737_, new_n29738_,
    new_n29739_, new_n29740_, new_n29741_, new_n29742_, new_n29743_,
    new_n29744_, new_n29745_, new_n29746_, new_n29747_, new_n29748_,
    new_n29749_, new_n29750_, new_n29751_, new_n29752_, new_n29753_,
    new_n29754_, new_n29755_, new_n29756_, new_n29757_, new_n29758_,
    new_n29759_, new_n29760_, new_n29761_, new_n29762_, new_n29763_,
    new_n29764_, new_n29765_, new_n29766_, new_n29767_, new_n29768_,
    new_n29769_, new_n29770_, new_n29771_, new_n29772_, new_n29773_,
    new_n29774_, new_n29775_, new_n29776_, new_n29777_, new_n29778_,
    new_n29779_, new_n29780_, new_n29781_, new_n29782_, new_n29783_,
    new_n29784_, new_n29785_, new_n29786_, new_n29787_, new_n29788_,
    new_n29789_, new_n29790_, new_n29791_, new_n29792_, new_n29793_,
    new_n29794_, new_n29795_, new_n29796_, new_n29797_, new_n29798_,
    new_n29799_, new_n29800_, new_n29801_, new_n29802_, new_n29803_,
    new_n29804_, new_n29805_, new_n29806_, new_n29807_, new_n29808_,
    new_n29809_, new_n29810_, new_n29811_, new_n29812_, new_n29813_,
    new_n29814_, new_n29815_, new_n29816_, new_n29817_, new_n29818_,
    new_n29819_, new_n29820_, new_n29821_, new_n29822_, new_n29823_,
    new_n29824_, new_n29825_, new_n29826_, new_n29827_, new_n29828_,
    new_n29829_, new_n29830_, new_n29831_, new_n29832_, new_n29833_,
    new_n29834_, new_n29835_, new_n29836_, new_n29837_, new_n29838_,
    new_n29839_, new_n29840_, new_n29841_, new_n29842_, new_n29843_,
    new_n29844_, new_n29845_, new_n29846_, new_n29847_, new_n29848_,
    new_n29849_, new_n29850_, new_n29851_, new_n29852_, new_n29853_,
    new_n29854_, new_n29855_, new_n29856_, new_n29857_, new_n29858_,
    new_n29859_, new_n29860_, new_n29861_, new_n29862_, new_n29863_,
    new_n29864_, new_n29865_, new_n29866_, new_n29867_, new_n29868_,
    new_n29869_, new_n29870_, new_n29871_, new_n29872_, new_n29873_,
    new_n29874_, new_n29875_, new_n29876_, new_n29877_, new_n29878_,
    new_n29879_, new_n29880_, new_n29881_, new_n29882_, new_n29883_,
    new_n29884_, new_n29885_, new_n29886_, new_n29887_, new_n29888_,
    new_n29889_, new_n29890_, new_n29891_, new_n29892_, new_n29893_,
    new_n29894_, new_n29895_, new_n29896_, new_n29897_, new_n29898_,
    new_n29899_, new_n29900_, new_n29901_, new_n29902_, new_n29903_,
    new_n29904_, new_n29905_, new_n29906_, new_n29907_, new_n29908_,
    new_n29909_, new_n29910_, new_n29911_, new_n29912_, new_n29913_,
    new_n29914_, new_n29915_, new_n29916_, new_n29917_, new_n29918_,
    new_n29919_, new_n29920_, new_n29921_, new_n29922_, new_n29923_,
    new_n29924_, new_n29925_, new_n29926_, new_n29927_, new_n29928_,
    new_n29929_, new_n29930_, new_n29931_, new_n29932_, new_n29933_,
    new_n29934_, new_n29935_, new_n29936_, new_n29937_, new_n29938_,
    new_n29939_, new_n29940_, new_n29941_, new_n29942_, new_n29943_,
    new_n29944_, new_n29945_, new_n29946_, new_n29947_, new_n29948_,
    new_n29949_, new_n29950_, new_n29951_, new_n29952_, new_n29953_,
    new_n29954_, new_n29955_, new_n29956_, new_n29957_, new_n29958_,
    new_n29959_, new_n29960_, new_n29961_, new_n29962_, new_n29963_,
    new_n29964_, new_n29965_, new_n29966_, new_n29967_, new_n29968_,
    new_n29969_, new_n29970_, new_n29971_, new_n29972_, new_n29973_,
    new_n29974_, new_n29975_, new_n29976_, new_n29977_, new_n29978_,
    new_n29979_, new_n29980_, new_n29981_, new_n29982_, new_n29983_,
    new_n29984_, new_n29985_, new_n29986_, new_n29987_, new_n29988_,
    new_n29989_, new_n29990_, new_n29991_, new_n29992_, new_n29993_,
    new_n29994_, new_n29995_, new_n29996_, new_n29997_, new_n29998_,
    new_n29999_, new_n30000_, new_n30001_, new_n30002_, new_n30003_,
    new_n30004_, new_n30005_, new_n30006_, new_n30007_, new_n30008_,
    new_n30009_, new_n30010_, new_n30011_, new_n30012_, new_n30013_,
    new_n30014_, new_n30015_, new_n30016_, new_n30017_, new_n30018_,
    new_n30019_, new_n30020_, new_n30021_, new_n30022_, new_n30023_,
    new_n30024_, new_n30025_, new_n30026_, new_n30027_, new_n30028_,
    new_n30029_, new_n30030_, new_n30031_, new_n30032_, new_n30033_,
    new_n30034_, new_n30035_, new_n30036_, new_n30037_, new_n30038_,
    new_n30039_, new_n30040_, new_n30041_, new_n30042_, new_n30043_,
    new_n30044_, new_n30045_, new_n30046_, new_n30047_, new_n30048_,
    new_n30049_, new_n30050_, new_n30051_, new_n30052_, new_n30053_,
    new_n30054_, new_n30055_, new_n30056_, new_n30057_, new_n30058_,
    new_n30059_, new_n30060_, new_n30061_, new_n30062_, new_n30063_,
    new_n30064_, new_n30065_, new_n30066_, new_n30067_, new_n30068_,
    new_n30069_, new_n30070_, new_n30071_, new_n30072_, new_n30073_,
    new_n30074_, new_n30075_, new_n30076_, new_n30077_, new_n30078_,
    new_n30079_, new_n30080_, new_n30081_, new_n30082_, new_n30083_,
    new_n30084_, new_n30085_, new_n30086_, new_n30087_, new_n30088_,
    new_n30089_, new_n30090_, new_n30091_, new_n30092_, new_n30093_,
    new_n30094_, new_n30095_, new_n30096_, new_n30097_, new_n30098_,
    new_n30099_, new_n30100_, new_n30101_, new_n30102_, new_n30103_,
    new_n30104_, new_n30105_, new_n30106_, new_n30107_, new_n30108_,
    new_n30109_, new_n30110_, new_n30111_, new_n30112_, new_n30113_,
    new_n30114_, new_n30115_, new_n30116_, new_n30117_, new_n30118_,
    new_n30119_, new_n30120_, new_n30121_, new_n30122_, new_n30123_,
    new_n30124_, new_n30125_, new_n30126_, new_n30127_, new_n30128_,
    new_n30129_, new_n30130_, new_n30131_, new_n30132_, new_n30133_,
    new_n30134_, new_n30135_, new_n30136_, new_n30137_, new_n30138_,
    new_n30139_, new_n30140_, new_n30141_, new_n30142_, new_n30143_,
    new_n30144_, new_n30145_, new_n30146_, new_n30147_, new_n30148_,
    new_n30149_, new_n30150_, new_n30151_, new_n30152_, new_n30153_,
    new_n30154_, new_n30155_, new_n30156_, new_n30157_, new_n30158_,
    new_n30159_, new_n30160_, new_n30161_, new_n30162_, new_n30163_,
    new_n30164_, new_n30165_, new_n30166_, new_n30167_, new_n30168_,
    new_n30169_, new_n30170_, new_n30171_, new_n30172_, new_n30173_,
    new_n30174_, new_n30175_, new_n30176_, new_n30177_, new_n30178_,
    new_n30179_, new_n30180_, new_n30181_, new_n30182_, new_n30183_,
    new_n30184_, new_n30185_, new_n30186_, new_n30187_, new_n30188_,
    new_n30189_, new_n30190_, new_n30191_, new_n30192_, new_n30193_,
    new_n30194_, new_n30195_, new_n30196_, new_n30197_, new_n30198_,
    new_n30199_, new_n30200_, new_n30201_, new_n30202_, new_n30203_,
    new_n30204_, new_n30205_, new_n30206_, new_n30207_, new_n30208_,
    new_n30209_, new_n30210_, new_n30211_, new_n30212_, new_n30213_,
    new_n30214_, new_n30215_, new_n30216_, new_n30217_, new_n30218_,
    new_n30219_, new_n30220_, new_n30221_, new_n30222_, new_n30223_,
    new_n30224_, new_n30225_, new_n30226_, new_n30227_, new_n30228_,
    new_n30229_, new_n30230_, new_n30231_, new_n30232_, new_n30233_,
    new_n30234_, new_n30235_, new_n30236_, new_n30237_, new_n30238_,
    new_n30239_, new_n30240_, new_n30241_, new_n30242_, new_n30243_,
    new_n30244_, new_n30245_, new_n30246_, new_n30247_, new_n30248_,
    new_n30249_, new_n30250_, new_n30251_, new_n30252_, new_n30253_,
    new_n30254_, new_n30255_, new_n30256_, new_n30257_, new_n30258_,
    new_n30259_, new_n30260_, new_n30261_, new_n30262_, new_n30263_,
    new_n30264_, new_n30265_, new_n30266_, new_n30267_, new_n30268_,
    new_n30269_, new_n30270_, new_n30271_, new_n30272_, new_n30273_,
    new_n30274_, new_n30275_, new_n30276_, new_n30277_, new_n30278_,
    new_n30279_, new_n30280_, new_n30281_, new_n30282_, new_n30283_,
    new_n30284_, new_n30285_, new_n30286_, new_n30287_, new_n30288_,
    new_n30289_, new_n30290_, new_n30291_, new_n30292_, new_n30293_,
    new_n30294_, new_n30295_, new_n30296_, new_n30297_, new_n30298_,
    new_n30299_, new_n30300_, new_n30301_, new_n30302_, new_n30303_,
    new_n30304_, new_n30305_, new_n30306_, new_n30307_, new_n30308_,
    new_n30309_, new_n30310_, new_n30311_, new_n30312_, new_n30313_,
    new_n30314_, new_n30315_, new_n30316_, new_n30317_, new_n30318_,
    new_n30319_, new_n30320_, new_n30321_, new_n30322_, new_n30323_,
    new_n30324_, new_n30325_, new_n30326_, new_n30327_, new_n30328_,
    new_n30329_, new_n30330_, new_n30331_, new_n30332_, new_n30333_,
    new_n30334_, new_n30335_, new_n30336_, new_n30337_, new_n30338_,
    new_n30339_, new_n30340_, new_n30341_, new_n30342_, new_n30343_,
    new_n30344_, new_n30345_, new_n30346_, new_n30347_, new_n30348_,
    new_n30349_, new_n30350_, new_n30351_, new_n30352_, new_n30353_,
    new_n30354_, new_n30355_, new_n30356_, new_n30357_, new_n30358_,
    new_n30359_, new_n30360_, new_n30361_, new_n30362_, new_n30363_,
    new_n30364_, new_n30365_, new_n30366_, new_n30367_, new_n30368_,
    new_n30369_, new_n30370_, new_n30371_, new_n30372_, new_n30373_,
    new_n30374_, new_n30375_, new_n30376_, new_n30377_, new_n30378_,
    new_n30379_, new_n30380_, new_n30381_, new_n30382_, new_n30383_,
    new_n30384_, new_n30385_, new_n30386_, new_n30387_, new_n30388_,
    new_n30389_, new_n30390_, new_n30391_, new_n30392_, new_n30393_,
    new_n30394_, new_n30395_, new_n30396_, new_n30397_, new_n30398_,
    new_n30399_, new_n30400_, new_n30401_, new_n30402_, new_n30403_,
    new_n30404_, new_n30405_, new_n30406_, new_n30407_, new_n30408_,
    new_n30409_, new_n30410_, new_n30411_, new_n30412_, new_n30413_,
    new_n30414_, new_n30415_, new_n30416_, new_n30417_, new_n30418_,
    new_n30419_, new_n30420_, new_n30421_, new_n30422_, new_n30423_,
    new_n30424_, new_n30425_, new_n30426_, new_n30427_, new_n30428_,
    new_n30429_, new_n30430_, new_n30431_, new_n30432_, new_n30433_,
    new_n30434_, new_n30435_, new_n30436_, new_n30437_, new_n30438_,
    new_n30439_, new_n30440_, new_n30441_, new_n30442_, new_n30443_,
    new_n30444_, new_n30445_, new_n30446_, new_n30447_, new_n30448_,
    new_n30449_, new_n30450_, new_n30451_, new_n30452_, new_n30453_,
    new_n30454_, new_n30455_, new_n30456_, new_n30457_, new_n30458_,
    new_n30459_, new_n30460_, new_n30461_, new_n30462_, new_n30463_,
    new_n30464_, new_n30465_, new_n30466_, new_n30467_, new_n30468_,
    new_n30469_, new_n30470_, new_n30471_, new_n30472_, new_n30473_,
    new_n30474_, new_n30475_, new_n30476_, new_n30477_, new_n30478_,
    new_n30479_, new_n30480_, new_n30481_, new_n30482_, new_n30483_,
    new_n30484_, new_n30485_, new_n30486_, new_n30487_, new_n30488_,
    new_n30489_, new_n30490_, new_n30491_, new_n30492_, new_n30493_,
    new_n30494_, new_n30495_, new_n30496_, new_n30497_, new_n30498_,
    new_n30499_, new_n30500_, new_n30501_, new_n30502_, new_n30503_,
    new_n30504_, new_n30505_, new_n30506_, new_n30507_, new_n30508_,
    new_n30509_, new_n30510_, new_n30511_, new_n30512_, new_n30513_,
    new_n30514_, new_n30515_, new_n30516_, new_n30517_, new_n30518_,
    new_n30519_, new_n30520_, new_n30521_, new_n30522_, new_n30523_,
    new_n30524_, new_n30525_, new_n30526_, new_n30527_, new_n30528_,
    new_n30529_, new_n30530_, new_n30531_, new_n30532_, new_n30533_,
    new_n30534_, new_n30535_, new_n30536_, new_n30537_, new_n30538_,
    new_n30539_, new_n30540_, new_n30541_, new_n30542_, new_n30543_,
    new_n30544_, new_n30545_, new_n30546_, new_n30547_, new_n30548_,
    new_n30549_, new_n30550_, new_n30551_, new_n30552_, new_n30553_,
    new_n30554_, new_n30555_, new_n30556_, new_n30557_, new_n30558_,
    new_n30559_, new_n30560_, new_n30561_, new_n30562_, new_n30563_,
    new_n30564_, new_n30565_, new_n30566_, new_n30567_, new_n30568_,
    new_n30569_, new_n30570_, new_n30571_, new_n30572_, new_n30573_,
    new_n30574_, new_n30575_, new_n30576_, new_n30577_, new_n30578_,
    new_n30579_, new_n30580_, new_n30581_, new_n30582_, new_n30583_,
    new_n30584_, new_n30585_, new_n30586_, new_n30587_, new_n30588_,
    new_n30589_, new_n30590_, new_n30591_, new_n30592_, new_n30593_,
    new_n30594_, new_n30595_, new_n30596_, new_n30597_, new_n30598_,
    new_n30599_, new_n30600_, new_n30601_, new_n30602_, new_n30603_,
    new_n30604_, new_n30605_, new_n30606_, new_n30607_, new_n30608_,
    new_n30609_, new_n30610_, new_n30611_, new_n30612_, new_n30613_,
    new_n30614_, new_n30615_, new_n30616_, new_n30617_, new_n30618_,
    new_n30619_, new_n30620_, new_n30621_, new_n30622_, new_n30623_,
    new_n30624_, new_n30625_, new_n30626_, new_n30627_, new_n30628_,
    new_n30629_, new_n30630_, new_n30631_, new_n30632_, new_n30633_,
    new_n30634_, new_n30635_, new_n30636_, new_n30637_, new_n30638_,
    new_n30639_, new_n30640_, new_n30641_, new_n30642_, new_n30643_,
    new_n30644_, new_n30645_, new_n30646_, new_n30647_, new_n30648_,
    new_n30649_, new_n30650_, new_n30651_, new_n30652_, new_n30653_,
    new_n30654_, new_n30655_, new_n30656_, new_n30657_, new_n30658_,
    new_n30659_, new_n30660_, new_n30661_, new_n30662_, new_n30663_,
    new_n30664_, new_n30665_, new_n30666_, new_n30667_, new_n30668_,
    new_n30669_, new_n30670_, new_n30671_, new_n30672_, new_n30673_,
    new_n30674_, new_n30675_, new_n30676_, new_n30677_, new_n30678_,
    new_n30679_, new_n30680_, new_n30681_, new_n30682_, new_n30683_,
    new_n30684_, new_n30685_, new_n30686_, new_n30687_, new_n30688_,
    new_n30689_, new_n30690_, new_n30691_, new_n30692_, new_n30693_,
    new_n30694_, new_n30695_, new_n30696_, new_n30697_, new_n30698_,
    new_n30699_, new_n30700_, new_n30701_, new_n30702_, new_n30703_,
    new_n30704_, new_n30705_, new_n30706_, new_n30707_, new_n30708_,
    new_n30709_, new_n30710_, new_n30711_, new_n30712_, new_n30713_,
    new_n30714_, new_n30715_, new_n30716_, new_n30717_, new_n30718_,
    new_n30719_, new_n30720_, new_n30721_, new_n30722_, new_n30723_,
    new_n30724_, new_n30725_, new_n30726_, new_n30727_, new_n30728_,
    new_n30729_, new_n30730_, new_n30731_, new_n30732_, new_n30733_,
    new_n30734_, new_n30735_, new_n30736_, new_n30737_, new_n30738_,
    new_n30739_, new_n30740_, new_n30741_, new_n30742_, new_n30743_,
    new_n30744_, new_n30745_, new_n30746_, new_n30747_, new_n30748_,
    new_n30749_, new_n30750_, new_n30751_, new_n30752_, new_n30753_,
    new_n30754_, new_n30755_, new_n30756_, new_n30757_, new_n30758_,
    new_n30759_, new_n30760_, new_n30761_, new_n30762_, new_n30763_,
    new_n30764_, new_n30765_, new_n30766_, new_n30767_, new_n30768_,
    new_n30769_, new_n30770_, new_n30771_, new_n30772_, new_n30773_,
    new_n30774_, new_n30775_, new_n30776_, new_n30777_, new_n30778_,
    new_n30779_, new_n30780_, new_n30781_, new_n30782_, new_n30783_,
    new_n30784_, new_n30785_, new_n30786_, new_n30787_, new_n30788_,
    new_n30789_, new_n30790_, new_n30791_, new_n30792_, new_n30793_,
    new_n30794_, new_n30795_, new_n30796_, new_n30797_, new_n30798_,
    new_n30799_, new_n30800_, new_n30801_, new_n30802_, new_n30803_,
    new_n30804_, new_n30805_, new_n30806_, new_n30807_, new_n30808_,
    new_n30809_, new_n30810_, new_n30811_, new_n30812_, new_n30813_,
    new_n30814_, new_n30815_, new_n30816_, new_n30817_, new_n30818_,
    new_n30819_, new_n30820_, new_n30821_, new_n30822_, new_n30823_,
    new_n30824_, new_n30825_, new_n30826_, new_n30827_, new_n30828_,
    new_n30829_, new_n30830_, new_n30831_, new_n30832_, new_n30833_,
    new_n30834_, new_n30835_, new_n30836_, new_n30837_, new_n30838_,
    new_n30839_, new_n30840_, new_n30841_, new_n30842_, new_n30843_,
    new_n30844_, new_n30845_, new_n30846_, new_n30847_, new_n30848_,
    new_n30849_, new_n30850_, new_n30851_, new_n30852_, new_n30853_,
    new_n30854_, new_n30855_, new_n30856_, new_n30857_, new_n30858_,
    new_n30859_, new_n30860_, new_n30861_, new_n30862_, new_n30863_,
    new_n30864_, new_n30865_, new_n30866_, new_n30867_, new_n30868_,
    new_n30869_, new_n30870_, new_n30871_, new_n30872_, new_n30873_,
    new_n30874_, new_n30875_, new_n30876_, new_n30877_, new_n30878_,
    new_n30879_, new_n30880_, new_n30881_, new_n30882_, new_n30883_,
    new_n30884_, new_n30885_, new_n30886_, new_n30887_, new_n30888_,
    new_n30889_, new_n30890_, new_n30891_, new_n30892_, new_n30893_,
    new_n30894_, new_n30895_, new_n30896_, new_n30897_, new_n30898_,
    new_n30899_, new_n30900_, new_n30901_, new_n30902_, new_n30903_,
    new_n30904_, new_n30905_, new_n30906_, new_n30907_, new_n30908_,
    new_n30909_, new_n30910_, new_n30911_, new_n30912_, new_n30913_,
    new_n30914_, new_n30915_, new_n30916_, new_n30917_, new_n30918_,
    new_n30919_, new_n30920_, new_n30921_, new_n30922_, new_n30923_,
    new_n30924_, new_n30925_, new_n30926_, new_n30927_, new_n30928_,
    new_n30929_, new_n30930_, new_n30931_, new_n30932_, new_n30933_,
    new_n30934_, new_n30935_, new_n30936_, new_n30937_, new_n30938_,
    new_n30939_, new_n30940_, new_n30941_, new_n30942_, new_n30943_,
    new_n30944_, new_n30945_, new_n30946_, new_n30947_, new_n30948_,
    new_n30949_, new_n30950_, new_n30951_, new_n30952_, new_n30953_,
    new_n30954_, new_n30955_, new_n30956_, new_n30957_, new_n30958_,
    new_n30959_, new_n30960_, new_n30961_, new_n30962_, new_n30963_,
    new_n30964_, new_n30965_, new_n30966_, new_n30967_, new_n30968_,
    new_n30969_, new_n30970_, new_n30971_, new_n30972_, new_n30973_,
    new_n30974_, new_n30975_, new_n30976_, new_n30977_, new_n30978_,
    new_n30979_, new_n30980_, new_n30981_, new_n30982_, new_n30983_,
    new_n30984_, new_n30985_, new_n30986_, new_n30987_, new_n30988_,
    new_n30989_, new_n30990_, new_n30991_, new_n30992_, new_n30993_,
    new_n30994_, new_n30995_, new_n30996_, new_n30997_, new_n30998_,
    new_n30999_, new_n31000_, new_n31001_, new_n31002_, new_n31003_,
    new_n31004_, new_n31005_, new_n31006_, new_n31007_, new_n31008_,
    new_n31009_, new_n31010_, new_n31011_, new_n31012_, new_n31013_,
    new_n31014_, new_n31015_, new_n31016_, new_n31017_, new_n31018_,
    new_n31019_, new_n31020_, new_n31021_, new_n31022_, new_n31023_,
    new_n31024_, new_n31025_, new_n31026_, new_n31027_, new_n31028_,
    new_n31029_, new_n31030_, new_n31031_, new_n31032_, new_n31033_,
    new_n31034_, new_n31035_, new_n31036_, new_n31037_, new_n31038_,
    new_n31039_, new_n31040_, new_n31041_, new_n31042_, new_n31043_,
    new_n31044_, new_n31045_, new_n31046_, new_n31047_, new_n31048_,
    new_n31049_, new_n31050_, new_n31051_, new_n31052_, new_n31053_,
    new_n31054_, new_n31055_, new_n31056_, new_n31057_, new_n31058_,
    new_n31059_, new_n31060_, new_n31061_, new_n31062_, new_n31063_,
    new_n31064_, new_n31065_, new_n31066_, new_n31067_, new_n31068_,
    new_n31069_, new_n31070_, new_n31071_, new_n31072_, new_n31073_,
    new_n31074_, new_n31075_, new_n31076_, new_n31077_, new_n31078_,
    new_n31079_, new_n31080_, new_n31081_, new_n31082_, new_n31083_,
    new_n31084_, new_n31085_, new_n31086_, new_n31087_, new_n31088_,
    new_n31089_, new_n31090_, new_n31091_, new_n31092_, new_n31093_,
    new_n31094_, new_n31095_, new_n31096_, new_n31097_, new_n31098_,
    new_n31099_, new_n31100_, new_n31101_, new_n31102_, new_n31103_,
    new_n31104_, new_n31105_, new_n31106_, new_n31107_, new_n31108_,
    new_n31109_, new_n31110_, new_n31111_, new_n31112_, new_n31113_,
    new_n31114_, new_n31115_, new_n31116_, new_n31117_, new_n31118_,
    new_n31119_, new_n31120_, new_n31121_, new_n31122_, new_n31123_,
    new_n31124_, new_n31125_, new_n31126_, new_n31127_, new_n31128_,
    new_n31129_, new_n31130_, new_n31131_, new_n31132_, new_n31133_,
    new_n31134_, new_n31135_, new_n31136_, new_n31137_, new_n31138_,
    new_n31139_, new_n31140_, new_n31141_, new_n31142_, new_n31143_,
    new_n31144_, new_n31145_, new_n31146_, new_n31147_, new_n31148_,
    new_n31149_, new_n31150_, new_n31151_, new_n31152_, new_n31153_,
    new_n31154_, new_n31155_, new_n31156_, new_n31157_, new_n31158_,
    new_n31159_, new_n31160_, new_n31161_, new_n31162_, new_n31163_,
    new_n31164_, new_n31165_, new_n31166_, new_n31167_, new_n31168_,
    new_n31169_, new_n31170_, new_n31171_, new_n31172_, new_n31173_,
    new_n31174_, new_n31175_, new_n31176_, new_n31177_, new_n31178_,
    new_n31179_, new_n31180_, new_n31181_, new_n31182_, new_n31183_,
    new_n31184_, new_n31185_, new_n31186_, new_n31187_, new_n31188_,
    new_n31189_, new_n31190_, new_n31191_, new_n31192_, new_n31193_,
    new_n31194_, new_n31195_, new_n31196_, new_n31197_, new_n31198_,
    new_n31199_, new_n31200_, new_n31201_, new_n31202_, new_n31203_,
    new_n31204_, new_n31205_, new_n31206_, new_n31207_, new_n31208_,
    new_n31209_, new_n31210_, new_n31211_, new_n31212_, new_n31213_,
    new_n31214_, new_n31215_, new_n31216_, new_n31217_, new_n31218_,
    new_n31219_, new_n31220_, new_n31221_, new_n31222_, new_n31223_,
    new_n31224_, new_n31225_, new_n31226_, new_n31227_, new_n31228_,
    new_n31229_, new_n31230_, new_n31231_, new_n31232_, new_n31233_,
    new_n31234_, new_n31235_, new_n31236_, new_n31237_, new_n31238_,
    new_n31239_, new_n31240_, new_n31241_, new_n31242_, new_n31243_,
    new_n31244_, new_n31245_, new_n31246_, new_n31247_, new_n31248_,
    new_n31249_, new_n31250_, new_n31251_, new_n31252_, new_n31253_,
    new_n31254_, new_n31255_, new_n31256_, new_n31257_, new_n31258_,
    new_n31259_, new_n31260_, new_n31261_, new_n31262_, new_n31263_,
    new_n31264_, new_n31265_, new_n31266_, new_n31267_, new_n31268_,
    new_n31269_, new_n31270_, new_n31271_, new_n31272_, new_n31273_,
    new_n31274_, new_n31275_, new_n31276_, new_n31277_, new_n31278_,
    new_n31279_, new_n31280_, new_n31281_, new_n31282_, new_n31283_,
    new_n31284_, new_n31285_, new_n31286_, new_n31287_, new_n31288_,
    new_n31289_, new_n31290_, new_n31291_, new_n31292_, new_n31293_,
    new_n31294_, new_n31295_, new_n31296_, new_n31297_, new_n31298_,
    new_n31299_, new_n31300_, new_n31301_, new_n31302_, new_n31303_,
    new_n31304_, new_n31305_, new_n31306_, new_n31307_, new_n31308_,
    new_n31309_, new_n31310_, new_n31311_, new_n31312_, new_n31313_,
    new_n31314_, new_n31315_, new_n31316_, new_n31317_, new_n31318_,
    new_n31319_, new_n31320_, new_n31321_, new_n31322_, new_n31323_,
    new_n31324_, new_n31325_, new_n31326_, new_n31327_, new_n31328_,
    new_n31329_, new_n31330_, new_n31331_, new_n31332_, new_n31333_,
    new_n31334_, new_n31335_, new_n31336_, new_n31337_, new_n31338_,
    new_n31339_, new_n31340_, new_n31341_, new_n31342_, new_n31343_,
    new_n31344_, new_n31345_, new_n31346_, new_n31347_, new_n31348_,
    new_n31349_, new_n31350_, new_n31351_, new_n31352_, new_n31353_,
    new_n31354_, new_n31355_, new_n31356_, new_n31357_, new_n31358_,
    new_n31359_, new_n31360_, new_n31361_, new_n31362_, new_n31363_,
    new_n31364_, new_n31365_, new_n31366_, new_n31367_, new_n31368_,
    new_n31369_, new_n31370_, new_n31371_, new_n31372_, new_n31373_,
    new_n31374_, new_n31375_, new_n31376_, new_n31377_, new_n31378_,
    new_n31379_, new_n31380_, new_n31381_, new_n31382_, new_n31383_,
    new_n31384_, new_n31385_, new_n31386_, new_n31387_, new_n31388_,
    new_n31389_, new_n31390_, new_n31391_, new_n31392_, new_n31393_,
    new_n31394_, new_n31395_, new_n31396_, new_n31397_, new_n31398_,
    new_n31399_, new_n31400_, new_n31401_, new_n31402_, new_n31403_,
    new_n31404_, new_n31405_, new_n31406_, new_n31407_, new_n31408_,
    new_n31409_, new_n31410_, new_n31411_, new_n31412_, new_n31413_,
    new_n31414_, new_n31415_, new_n31416_, new_n31417_, new_n31418_,
    new_n31419_, new_n31420_, new_n31421_, new_n31422_, new_n31423_,
    new_n31424_, new_n31425_, new_n31426_, new_n31427_, new_n31428_,
    new_n31429_, new_n31430_, new_n31431_, new_n31432_, new_n31433_,
    new_n31434_, new_n31435_, new_n31436_, new_n31437_, new_n31438_,
    new_n31439_, new_n31440_, new_n31441_, new_n31442_, new_n31443_,
    new_n31444_, new_n31445_, new_n31446_, new_n31447_, new_n31448_,
    new_n31449_, new_n31450_, new_n31451_, new_n31452_, new_n31453_,
    new_n31454_, new_n31455_, new_n31456_, new_n31457_, new_n31458_,
    new_n31459_, new_n31460_, new_n31461_, new_n31462_, new_n31463_,
    new_n31464_, new_n31465_, new_n31466_, new_n31467_, new_n31468_,
    new_n31469_, new_n31470_, new_n31471_, new_n31472_, new_n31473_,
    new_n31474_, new_n31475_, new_n31476_, new_n31477_, new_n31478_,
    new_n31479_, new_n31480_, new_n31481_, new_n31482_, new_n31483_,
    new_n31484_, new_n31485_, new_n31486_, new_n31487_, new_n31488_,
    new_n31489_, new_n31490_, new_n31491_, new_n31492_, new_n31493_,
    new_n31494_, new_n31495_, new_n31496_, new_n31497_, new_n31498_,
    new_n31499_, new_n31500_, new_n31501_, new_n31502_, new_n31503_,
    new_n31504_, new_n31505_, new_n31506_, new_n31507_, new_n31508_,
    new_n31509_, new_n31510_, new_n31511_, new_n31512_, new_n31513_,
    new_n31514_, new_n31515_, new_n31516_, new_n31517_, new_n31518_,
    new_n31519_, new_n31520_, new_n31521_, new_n31522_, new_n31523_,
    new_n31524_, new_n31525_, new_n31526_, new_n31527_, new_n31528_,
    new_n31529_, new_n31530_, new_n31531_, new_n31532_, new_n31533_,
    new_n31534_, new_n31535_, new_n31536_, new_n31537_, new_n31538_,
    new_n31539_, new_n31540_, new_n31541_, new_n31542_, new_n31543_,
    new_n31544_, new_n31545_, new_n31546_, new_n31547_, new_n31548_,
    new_n31549_, new_n31550_, new_n31551_, new_n31552_, new_n31553_,
    new_n31554_, new_n31555_, new_n31556_, new_n31557_, new_n31558_,
    new_n31559_, new_n31560_, new_n31561_, new_n31562_, new_n31563_,
    new_n31564_, new_n31565_, new_n31566_, new_n31567_, new_n31568_,
    new_n31569_, new_n31570_, new_n31571_, new_n31572_, new_n31573_,
    new_n31574_, new_n31575_, new_n31576_, new_n31577_, new_n31578_,
    new_n31579_, new_n31580_, new_n31581_, new_n31582_, new_n31583_,
    new_n31584_, new_n31585_, new_n31586_, new_n31587_, new_n31588_,
    new_n31589_, new_n31590_, new_n31591_, new_n31592_, new_n31593_,
    new_n31594_, new_n31595_, new_n31596_, new_n31597_, new_n31598_,
    new_n31599_, new_n31600_, new_n31601_, new_n31602_, new_n31603_,
    new_n31604_, new_n31605_, new_n31606_, new_n31607_, new_n31608_,
    new_n31609_, new_n31610_, new_n31611_, new_n31612_, new_n31613_,
    new_n31614_, new_n31615_, new_n31616_, new_n31617_, new_n31618_,
    new_n31619_, new_n31620_, new_n31621_, new_n31622_, new_n31623_,
    new_n31624_, new_n31625_, new_n31626_, new_n31627_, new_n31628_,
    new_n31629_, new_n31630_, new_n31631_, new_n31632_, new_n31633_,
    new_n31634_, new_n31635_, new_n31636_, new_n31637_, new_n31638_,
    new_n31639_, new_n31640_, new_n31641_, new_n31642_, new_n31643_,
    new_n31644_, new_n31645_, new_n31646_, new_n31647_, new_n31648_,
    new_n31649_, new_n31650_, new_n31651_, new_n31652_, new_n31653_,
    new_n31654_, new_n31655_, new_n31656_, new_n31657_, new_n31658_,
    new_n31659_, new_n31660_, new_n31661_, new_n31662_, new_n31663_,
    new_n31664_, new_n31665_, new_n31666_, new_n31667_, new_n31668_,
    new_n31669_, new_n31670_, new_n31671_, new_n31672_, new_n31673_,
    new_n31674_, new_n31675_, new_n31676_, new_n31677_, new_n31678_,
    new_n31679_, new_n31680_, new_n31681_, new_n31682_, new_n31683_,
    new_n31684_, new_n31685_, new_n31686_, new_n31687_, new_n31688_,
    new_n31689_, new_n31690_, new_n31691_, new_n31692_, new_n31693_,
    new_n31694_, new_n31695_, new_n31696_, new_n31697_, new_n31698_,
    new_n31699_, new_n31700_, new_n31701_, new_n31702_, new_n31703_,
    new_n31704_, new_n31705_, new_n31706_, new_n31707_, new_n31708_,
    new_n31709_, new_n31710_, new_n31711_, new_n31712_, new_n31713_,
    new_n31714_, new_n31715_, new_n31716_, new_n31717_, new_n31718_,
    new_n31719_, new_n31720_, new_n31721_, new_n31722_, new_n31723_,
    new_n31724_, new_n31725_, new_n31726_, new_n31727_, new_n31728_,
    new_n31729_, new_n31730_, new_n31731_, new_n31732_, new_n31733_,
    new_n31734_, new_n31735_, new_n31736_, new_n31737_, new_n31738_,
    new_n31739_, new_n31740_, new_n31741_, new_n31742_, new_n31743_,
    new_n31744_, new_n31745_, new_n31746_, new_n31747_, new_n31748_,
    new_n31749_, new_n31750_, new_n31751_, new_n31752_, new_n31753_,
    new_n31754_, new_n31755_, new_n31756_, new_n31757_, new_n31758_,
    new_n31759_, new_n31760_, new_n31761_, new_n31762_, new_n31763_,
    new_n31764_, new_n31765_, new_n31766_, new_n31767_, new_n31768_,
    new_n31769_, new_n31770_, new_n31771_, new_n31772_, new_n31773_,
    new_n31774_, new_n31775_, new_n31776_, new_n31777_, new_n31778_,
    new_n31779_, new_n31780_, new_n31781_, new_n31782_, new_n31783_,
    new_n31784_, new_n31785_, new_n31786_, new_n31787_, new_n31788_,
    new_n31789_, new_n31790_, new_n31791_, new_n31792_, new_n31793_,
    new_n31794_, new_n31795_, new_n31796_, new_n31797_, new_n31798_,
    new_n31799_, new_n31800_, new_n31801_, new_n31802_, new_n31803_,
    new_n31804_, new_n31805_, new_n31806_, new_n31807_, new_n31808_,
    new_n31809_, new_n31810_, new_n31811_, new_n31812_, new_n31813_,
    new_n31814_, new_n31815_, new_n31816_, new_n31817_, new_n31818_,
    new_n31819_, new_n31820_, new_n31821_, new_n31822_, new_n31823_,
    new_n31824_, new_n31825_, new_n31826_, new_n31827_, new_n31828_,
    new_n31829_, new_n31830_, new_n31831_, new_n31832_, new_n31833_,
    new_n31834_, new_n31835_, new_n31836_, new_n31837_, new_n31838_,
    new_n31839_, new_n31840_, new_n31841_, new_n31842_, new_n31843_,
    new_n31844_, new_n31845_, new_n31846_, new_n31847_, new_n31848_,
    new_n31849_, new_n31850_, new_n31851_, new_n31852_, new_n31853_,
    new_n31854_, new_n31855_, new_n31856_, new_n31857_, new_n31858_,
    new_n31859_, new_n31860_, new_n31861_, new_n31862_, new_n31863_,
    new_n31864_, new_n31865_, new_n31866_, new_n31867_, new_n31868_,
    new_n31869_, new_n31870_, new_n31871_, new_n31872_, new_n31873_,
    new_n31874_, new_n31875_, new_n31876_, new_n31877_, new_n31878_,
    new_n31879_, new_n31880_, new_n31881_, new_n31882_, new_n31883_,
    new_n31884_, new_n31885_, new_n31886_, new_n31887_, new_n31888_,
    new_n31889_, new_n31890_, new_n31891_, new_n31892_, new_n31893_,
    new_n31894_, new_n31895_, new_n31896_, new_n31897_, new_n31898_,
    new_n31899_, new_n31900_, new_n31901_, new_n31902_, new_n31903_,
    new_n31904_, new_n31905_, new_n31906_, new_n31907_, new_n31908_,
    new_n31909_, new_n31910_, new_n31911_, new_n31912_, new_n31913_,
    new_n31914_, new_n31915_, new_n31916_, new_n31917_, new_n31918_,
    new_n31919_, new_n31920_, new_n31921_, new_n31922_, new_n31923_,
    new_n31924_, new_n31925_, new_n31926_, new_n31927_, new_n31928_,
    new_n31929_, new_n31930_, new_n31931_, new_n31932_, new_n31933_,
    new_n31934_, new_n31935_, new_n31936_, new_n31937_, new_n31938_,
    new_n31939_, new_n31940_, new_n31941_, new_n31942_, new_n31943_,
    new_n31944_, new_n31945_, new_n31946_, new_n31947_, new_n31948_,
    new_n31949_, new_n31950_, new_n31951_, new_n31952_, new_n31953_,
    new_n31954_, new_n31955_, new_n31956_, new_n31957_, new_n31958_,
    new_n31959_, new_n31960_, new_n31961_, new_n31962_, new_n31963_,
    new_n31964_, new_n31965_, new_n31966_, new_n31967_, new_n31968_,
    new_n31969_, new_n31970_, new_n31971_, new_n31972_, new_n31973_,
    new_n31974_, new_n31975_, new_n31976_, new_n31977_, new_n31978_,
    new_n31979_, new_n31980_, new_n31981_, new_n31982_, new_n31983_,
    new_n31984_, new_n31985_, new_n31986_, new_n31987_, new_n31988_,
    new_n31989_, new_n31990_, new_n31991_, new_n31992_, new_n31993_,
    new_n31994_, new_n31995_, new_n31996_, new_n31997_, new_n31998_,
    new_n31999_, new_n32000_, new_n32001_, new_n32002_, new_n32003_,
    new_n32004_, new_n32005_, new_n32006_, new_n32007_, new_n32008_,
    new_n32009_, new_n32010_, new_n32011_, new_n32012_, new_n32013_,
    new_n32014_, new_n32015_, new_n32016_, new_n32017_, new_n32018_,
    new_n32019_, new_n32020_, new_n32021_, new_n32022_, new_n32023_,
    new_n32024_, new_n32025_, new_n32026_, new_n32027_, new_n32028_,
    new_n32029_, new_n32030_, new_n32031_, new_n32032_, new_n32033_,
    new_n32034_, new_n32035_, new_n32036_, new_n32037_, new_n32038_,
    new_n32039_, new_n32040_, new_n32041_, new_n32042_, new_n32043_,
    new_n32044_, new_n32045_, new_n32046_, new_n32047_, new_n32048_,
    new_n32049_, new_n32050_, new_n32051_, new_n32052_, new_n32053_,
    new_n32054_, new_n32055_, new_n32056_, new_n32057_, new_n32058_,
    new_n32059_, new_n32060_, new_n32061_, new_n32062_, new_n32063_,
    new_n32064_, new_n32065_, new_n32066_, new_n32067_, new_n32068_,
    new_n32069_, new_n32070_, new_n32071_, new_n32072_, new_n32073_,
    new_n32074_, new_n32075_, new_n32076_, new_n32077_, new_n32078_,
    new_n32079_, new_n32080_, new_n32081_, new_n32082_, new_n32083_,
    new_n32084_, new_n32085_, new_n32086_, new_n32087_, new_n32088_,
    new_n32089_, new_n32090_, new_n32091_, new_n32092_, new_n32093_,
    new_n32094_, new_n32095_, new_n32096_, new_n32097_, new_n32098_,
    new_n32099_, new_n32100_, new_n32101_, new_n32102_, new_n32103_,
    new_n32104_, new_n32105_, new_n32106_, new_n32107_, new_n32108_,
    new_n32109_, new_n32110_, new_n32111_, new_n32112_, new_n32113_,
    new_n32114_, new_n32115_, new_n32116_, new_n32117_, new_n32118_,
    new_n32119_, new_n32120_, new_n32121_, new_n32122_, new_n32123_,
    new_n32124_, new_n32125_, new_n32126_, new_n32127_, new_n32128_,
    new_n32129_, new_n32130_, new_n32131_, new_n32132_, new_n32133_,
    new_n32134_, new_n32135_, new_n32136_, new_n32137_, new_n32138_,
    new_n32139_, new_n32140_, new_n32141_, new_n32142_, new_n32143_,
    new_n32144_, new_n32145_, new_n32146_, new_n32147_, new_n32148_,
    new_n32149_, new_n32150_, new_n32151_, new_n32152_, new_n32153_,
    new_n32154_, new_n32155_, new_n32156_, new_n32157_, new_n32158_,
    new_n32159_, new_n32160_, new_n32161_, new_n32162_, new_n32163_,
    new_n32164_, new_n32165_, new_n32166_, new_n32167_, new_n32168_,
    new_n32169_, new_n32170_, new_n32171_, new_n32172_, new_n32173_,
    new_n32174_, new_n32175_, new_n32176_, new_n32177_, new_n32178_,
    new_n32179_, new_n32180_, new_n32181_, new_n32182_, new_n32183_,
    new_n32184_, new_n32185_, new_n32186_, new_n32187_, new_n32188_,
    new_n32189_, new_n32190_, new_n32191_, new_n32192_, new_n32193_,
    new_n32194_, new_n32195_, new_n32196_, new_n32197_, new_n32198_,
    new_n32199_, new_n32200_, new_n32201_, new_n32202_, new_n32203_,
    new_n32204_, new_n32205_, new_n32206_, new_n32207_, new_n32208_,
    new_n32209_, new_n32210_, new_n32211_, new_n32212_, new_n32213_,
    new_n32214_, new_n32215_, new_n32216_, new_n32217_, new_n32218_,
    new_n32219_, new_n32220_, new_n32221_, new_n32222_, new_n32223_,
    new_n32224_, new_n32225_, new_n32226_, new_n32227_, new_n32228_,
    new_n32229_, new_n32230_, new_n32231_, new_n32232_, new_n32233_,
    new_n32234_, new_n32235_, new_n32236_, new_n32237_, new_n32238_,
    new_n32239_, new_n32240_, new_n32241_, new_n32242_, new_n32243_,
    new_n32244_, new_n32245_, new_n32246_, new_n32247_, new_n32248_,
    new_n32249_, new_n32250_, new_n32251_, new_n32252_, new_n32253_,
    new_n32254_, new_n32255_, new_n32256_, new_n32257_, new_n32258_,
    new_n32259_, new_n32260_, new_n32261_, new_n32262_, new_n32263_,
    new_n32264_, new_n32265_, new_n32266_, new_n32267_, new_n32268_,
    new_n32269_, new_n32270_, new_n32271_, new_n32272_, new_n32273_,
    new_n32274_, new_n32275_, new_n32276_, new_n32277_, new_n32278_,
    new_n32279_, new_n32280_, new_n32281_, new_n32282_, new_n32283_,
    new_n32284_, new_n32285_, new_n32286_, new_n32287_, new_n32288_,
    new_n32289_, new_n32290_, new_n32291_, new_n32292_, new_n32293_,
    new_n32294_, new_n32295_, new_n32296_, new_n32297_, new_n32298_,
    new_n32299_, new_n32300_, new_n32301_, new_n32302_, new_n32303_,
    new_n32304_, new_n32305_, new_n32306_, new_n32307_, new_n32308_,
    new_n32309_, new_n32310_, new_n32311_, new_n32312_, new_n32313_,
    new_n32314_, new_n32315_, new_n32316_, new_n32317_, new_n32318_,
    new_n32319_, new_n32320_, new_n32321_, new_n32322_, new_n32323_,
    new_n32324_, new_n32325_, new_n32326_, new_n32327_, new_n32328_,
    new_n32329_, new_n32330_, new_n32331_, new_n32332_, new_n32333_,
    new_n32334_, new_n32335_, new_n32336_, new_n32337_, new_n32338_,
    new_n32339_, new_n32340_, new_n32341_, new_n32342_, new_n32343_,
    new_n32344_, new_n32345_, new_n32346_, new_n32347_, new_n32348_,
    new_n32349_, new_n32350_, new_n32351_, new_n32352_, new_n32353_,
    new_n32354_, new_n32355_, new_n32356_, new_n32357_, new_n32358_,
    new_n32359_, new_n32360_, new_n32361_, new_n32362_, new_n32363_,
    new_n32364_, new_n32365_, new_n32366_, new_n32367_, new_n32368_,
    new_n32369_, new_n32370_, new_n32371_, new_n32372_, new_n32373_,
    new_n32374_, new_n32375_, new_n32376_, new_n32377_, new_n32378_,
    new_n32379_, new_n32380_, new_n32381_, new_n32382_, new_n32383_,
    new_n32384_, new_n32385_, new_n32386_, new_n32387_, new_n32388_,
    new_n32389_, new_n32390_, new_n32391_, new_n32392_, new_n32393_,
    new_n32394_, new_n32395_, new_n32396_, new_n32397_, new_n32398_,
    new_n32399_, new_n32400_, new_n32401_, new_n32402_, new_n32403_,
    new_n32404_, new_n32405_, new_n32406_, new_n32407_, new_n32408_,
    new_n32409_, new_n32410_, new_n32411_, new_n32412_, new_n32413_,
    new_n32414_, new_n32415_, new_n32416_, new_n32417_, new_n32418_,
    new_n32419_, new_n32420_, new_n32421_, new_n32422_, new_n32423_,
    new_n32424_, new_n32425_, new_n32426_, new_n32427_, new_n32428_,
    new_n32429_, new_n32430_, new_n32431_, new_n32432_, new_n32433_,
    new_n32434_, new_n32435_, new_n32436_, new_n32437_, new_n32438_,
    new_n32439_, new_n32440_, new_n32441_, new_n32442_, new_n32443_,
    new_n32444_, new_n32445_, new_n32446_, new_n32447_, new_n32448_,
    new_n32449_, new_n32450_, new_n32451_, new_n32452_, new_n32453_,
    new_n32454_, new_n32455_, new_n32456_, new_n32457_, new_n32458_,
    new_n32459_, new_n32460_, new_n32461_, new_n32462_, new_n32463_,
    new_n32464_, new_n32465_, new_n32466_, new_n32467_, new_n32468_,
    new_n32469_, new_n32470_, new_n32471_, new_n32472_, new_n32473_,
    new_n32474_, new_n32475_, new_n32476_, new_n32477_, new_n32478_,
    new_n32479_, new_n32480_, new_n32481_, new_n32482_, new_n32483_,
    new_n32484_, new_n32485_, new_n32486_, new_n32487_, new_n32488_,
    new_n32489_, new_n32490_, new_n32491_, new_n32492_, new_n32493_,
    new_n32494_, new_n32495_, new_n32496_, new_n32497_, new_n32498_,
    new_n32499_, new_n32500_, new_n32501_, new_n32502_, new_n32503_,
    new_n32504_, new_n32505_, new_n32506_, new_n32507_, new_n32508_,
    new_n32509_, new_n32510_, new_n32511_, new_n32512_, new_n32513_,
    new_n32514_, new_n32515_, new_n32516_, new_n32517_, new_n32518_,
    new_n32519_, new_n32520_, new_n32521_, new_n32522_, new_n32523_,
    new_n32524_, new_n32525_, new_n32526_, new_n32527_, new_n32528_,
    new_n32529_, new_n32530_, new_n32531_, new_n32532_, new_n32533_,
    new_n32534_, new_n32535_, new_n32536_, new_n32537_, new_n32538_,
    new_n32539_, new_n32540_, new_n32541_, new_n32542_, new_n32543_,
    new_n32544_, new_n32545_, new_n32546_, new_n32547_, new_n32548_,
    new_n32549_, new_n32550_, new_n32551_, new_n32552_, new_n32553_,
    new_n32554_, new_n32555_, new_n32556_, new_n32557_, new_n32558_,
    new_n32559_, new_n32560_, new_n32561_, new_n32562_, new_n32563_,
    new_n32564_, new_n32565_, new_n32566_, new_n32567_, new_n32568_,
    new_n32569_, new_n32570_, new_n32571_, new_n32572_, new_n32573_,
    new_n32574_, new_n32575_, new_n32576_, new_n32577_, new_n32578_,
    new_n32579_, new_n32580_, new_n32581_, new_n32582_, new_n32583_,
    new_n32584_, new_n32585_, new_n32586_, new_n32587_, new_n32588_,
    new_n32589_, new_n32590_, new_n32591_, new_n32592_, new_n32593_,
    new_n32594_, new_n32595_, new_n32596_, new_n32597_, new_n32598_,
    new_n32599_, new_n32600_, new_n32601_, new_n32602_, new_n32603_,
    new_n32604_, new_n32605_, new_n32606_, new_n32607_, new_n32608_,
    new_n32609_, new_n32610_, new_n32611_, new_n32612_, new_n32613_,
    new_n32614_, new_n32615_, new_n32616_, new_n32617_, new_n32618_,
    new_n32619_, new_n32620_, new_n32621_, new_n32622_, new_n32623_,
    new_n32624_, new_n32625_, new_n32626_, new_n32627_, new_n32628_,
    new_n32629_, new_n32630_, new_n32631_, new_n32632_, new_n32633_,
    new_n32634_, new_n32635_, new_n32636_, new_n32637_, new_n32638_,
    new_n32639_, new_n32640_, new_n32641_, new_n32642_, new_n32643_,
    new_n32644_, new_n32645_, new_n32646_, new_n32647_, new_n32648_,
    new_n32649_, new_n32650_, new_n32651_, new_n32652_, new_n32653_,
    new_n32654_, new_n32655_, new_n32656_, new_n32657_, new_n32658_,
    new_n32659_, new_n32660_, new_n32661_, new_n32662_, new_n32663_,
    new_n32664_, new_n32665_, new_n32666_, new_n32667_, new_n32668_,
    new_n32669_, new_n32670_, new_n32671_, new_n32672_, new_n32673_,
    new_n32674_, new_n32675_, new_n32676_, new_n32677_, new_n32678_,
    new_n32679_, new_n32680_, new_n32681_, new_n32682_, new_n32683_,
    new_n32684_, new_n32685_, new_n32686_, new_n32687_, new_n32688_,
    new_n32689_, new_n32690_, new_n32691_, new_n32692_, new_n32693_,
    new_n32694_, new_n32695_, new_n32696_, new_n32697_, new_n32698_,
    new_n32699_, new_n32700_, new_n32701_, new_n32702_, new_n32703_,
    new_n32704_, new_n32705_, new_n32706_, new_n32707_, new_n32708_,
    new_n32709_, new_n32710_, new_n32711_, new_n32712_, new_n32713_,
    new_n32714_, new_n32715_, new_n32716_, new_n32717_, new_n32718_,
    new_n32719_, new_n32720_, new_n32721_, new_n32722_, new_n32723_,
    new_n32724_, new_n32725_, new_n32726_, new_n32727_, new_n32728_,
    new_n32729_, new_n32730_, new_n32731_, new_n32732_, new_n32733_,
    new_n32734_, new_n32735_, new_n32736_, new_n32737_, new_n32738_,
    new_n32739_, new_n32740_, new_n32741_, new_n32742_, new_n32743_,
    new_n32744_, new_n32745_, new_n32746_, new_n32747_, new_n32748_,
    new_n32749_, new_n32750_, new_n32751_, new_n32752_, new_n32753_,
    new_n32754_, new_n32755_, new_n32756_, new_n32757_, new_n32758_,
    new_n32759_, new_n32760_, new_n32761_, new_n32762_, new_n32763_,
    new_n32764_, new_n32765_, new_n32766_, new_n32767_, new_n32768_,
    new_n32769_, new_n32770_, new_n32771_, new_n32772_, new_n32773_,
    new_n32774_, new_n32775_, new_n32776_, new_n32777_, new_n32778_,
    new_n32779_, new_n32780_, new_n32781_, new_n32782_, new_n32783_,
    new_n32784_, new_n32785_, new_n32786_, new_n32787_, new_n32788_,
    new_n32789_, new_n32790_, new_n32791_, new_n32792_, new_n32793_,
    new_n32794_, new_n32795_, new_n32796_, new_n32797_, new_n32798_,
    new_n32799_, new_n32800_, new_n32801_, new_n32802_, new_n32803_,
    new_n32804_, new_n32805_, new_n32806_, new_n32807_, new_n32808_,
    new_n32809_, new_n32810_, new_n32811_, new_n32812_, new_n32813_,
    new_n32814_, new_n32815_, new_n32816_, new_n32817_, new_n32818_,
    new_n32819_, new_n32820_, new_n32821_, new_n32822_, new_n32823_,
    new_n32824_, new_n32825_, new_n32826_, new_n32827_, new_n32828_,
    new_n32829_, new_n32830_, new_n32831_, new_n32832_, new_n32833_,
    new_n32834_, new_n32835_, new_n32836_, new_n32837_, new_n32838_,
    new_n32839_, new_n32840_, new_n32841_, new_n32842_, new_n32843_,
    new_n32844_, new_n32845_, new_n32846_, new_n32847_, new_n32848_,
    new_n32849_, new_n32850_, new_n32851_, new_n32852_, new_n32853_,
    new_n32854_, new_n32855_, new_n32856_, new_n32857_, new_n32858_,
    new_n32859_, new_n32860_, new_n32861_, new_n32862_, new_n32863_,
    new_n32864_, new_n32865_, new_n32866_, new_n32867_, new_n32868_,
    new_n32869_, new_n32870_, new_n32871_, new_n32872_, new_n32873_,
    new_n32874_, new_n32875_, new_n32876_, new_n32877_, new_n32878_,
    new_n32879_, new_n32880_, new_n32881_, new_n32882_, new_n32883_,
    new_n32884_, new_n32885_, new_n32886_, new_n32887_, new_n32888_,
    new_n32889_, new_n32890_, new_n32891_, new_n32892_, new_n32893_,
    new_n32894_, new_n32895_, new_n32896_, new_n32897_, new_n32898_,
    new_n32899_, new_n32900_, new_n32901_, new_n32902_, new_n32903_,
    new_n32904_, new_n32905_, new_n32906_, new_n32907_, new_n32908_,
    new_n32909_, new_n32910_, new_n32911_, new_n32912_, new_n32913_,
    new_n32914_, new_n32915_, new_n32916_, new_n32917_, new_n32918_,
    new_n32919_, new_n32920_, new_n32921_, new_n32922_, new_n32923_,
    new_n32924_, new_n32925_, new_n32926_, new_n32927_, new_n32928_,
    new_n32929_, new_n32930_, new_n32931_, new_n32932_, new_n32933_,
    new_n32934_, new_n32935_, new_n32936_, new_n32937_, new_n32938_,
    new_n32939_, new_n32940_, new_n32941_, new_n32942_, new_n32943_,
    new_n32944_, new_n32945_, new_n32946_, new_n32947_, new_n32948_,
    new_n32949_, new_n32950_, new_n32951_, new_n32952_, new_n32953_,
    new_n32954_, new_n32955_, new_n32956_, new_n32957_, new_n32958_,
    new_n32959_, new_n32960_, new_n32961_, new_n32962_, new_n32963_,
    new_n32964_, new_n32965_, new_n32966_, new_n32967_, new_n32968_,
    new_n32969_, new_n32970_, new_n32971_, new_n32972_, new_n32973_,
    new_n32974_, new_n32975_, new_n32976_, new_n32977_, new_n32978_,
    new_n32979_, new_n32980_, new_n32981_, new_n32982_, new_n32983_,
    new_n32984_, new_n32985_, new_n32986_, new_n32987_, new_n32988_,
    new_n32989_, new_n32990_, new_n32991_, new_n32992_, new_n32993_,
    new_n32994_, new_n32995_, new_n32996_, new_n32997_, new_n32998_,
    new_n32999_, new_n33000_, new_n33001_, new_n33002_, new_n33003_,
    new_n33004_, new_n33005_, new_n33006_, new_n33007_, new_n33008_,
    new_n33009_, new_n33010_, new_n33011_, new_n33012_, new_n33013_,
    new_n33014_, new_n33015_, new_n33016_, new_n33017_, new_n33018_,
    new_n33019_, new_n33020_, new_n33021_, new_n33022_, new_n33023_,
    new_n33024_, new_n33025_, new_n33026_, new_n33027_, new_n33028_,
    new_n33029_, new_n33030_, new_n33031_, new_n33032_, new_n33033_,
    new_n33034_, new_n33035_, new_n33036_, new_n33037_, new_n33038_,
    new_n33039_, new_n33040_, new_n33041_, new_n33042_, new_n33043_,
    new_n33044_, new_n33045_, new_n33046_, new_n33047_, new_n33048_,
    new_n33049_, new_n33050_, new_n33051_, new_n33052_, new_n33053_,
    new_n33054_, new_n33055_, new_n33056_, new_n33057_, new_n33058_,
    new_n33059_, new_n33060_, new_n33061_, new_n33062_, new_n33063_,
    new_n33064_, new_n33065_, new_n33066_, new_n33067_, new_n33068_,
    new_n33069_, new_n33070_, new_n33071_, new_n33072_, new_n33073_,
    new_n33074_, new_n33075_, new_n33076_, new_n33077_, new_n33078_,
    new_n33079_, new_n33080_, new_n33081_, new_n33082_, new_n33083_,
    new_n33084_, new_n33085_, new_n33086_, new_n33087_, new_n33088_,
    new_n33089_, new_n33090_, new_n33091_, new_n33092_, new_n33093_,
    new_n33094_, new_n33095_, new_n33096_, new_n33097_, new_n33098_,
    new_n33099_, new_n33100_, new_n33101_, new_n33102_, new_n33103_,
    new_n33104_, new_n33105_, new_n33106_, new_n33107_, new_n33108_,
    new_n33109_, new_n33110_, new_n33111_, new_n33112_, new_n33113_,
    new_n33114_, new_n33115_, new_n33116_, new_n33117_, new_n33118_,
    new_n33119_, new_n33120_, new_n33121_, new_n33122_, new_n33123_,
    new_n33124_, new_n33125_, new_n33126_, new_n33127_, new_n33128_,
    new_n33129_, new_n33130_, new_n33131_, new_n33132_, new_n33133_,
    new_n33134_, new_n33135_, new_n33136_, new_n33137_, new_n33138_,
    new_n33139_, new_n33140_, new_n33141_, new_n33142_, new_n33143_,
    new_n33144_, new_n33145_, new_n33146_, new_n33147_, new_n33148_,
    new_n33149_, new_n33150_, new_n33151_, new_n33152_, new_n33153_,
    new_n33154_, new_n33155_, new_n33156_, new_n33157_, new_n33158_,
    new_n33159_, new_n33160_, new_n33161_, new_n33162_, new_n33163_,
    new_n33164_, new_n33165_, new_n33166_, new_n33167_, new_n33168_,
    new_n33169_, new_n33170_, new_n33171_, new_n33172_, new_n33173_,
    new_n33174_, new_n33175_, new_n33176_, new_n33177_, new_n33178_,
    new_n33179_, new_n33180_, new_n33181_, new_n33182_, new_n33183_,
    new_n33184_, new_n33185_, new_n33186_, new_n33187_, new_n33188_,
    new_n33189_, new_n33190_, new_n33191_, new_n33192_, new_n33193_,
    new_n33194_, new_n33195_, new_n33196_, new_n33197_, new_n33198_,
    new_n33199_, new_n33200_, new_n33201_, new_n33202_, new_n33203_,
    new_n33204_, new_n33205_, new_n33206_, new_n33207_, new_n33208_,
    new_n33209_, new_n33210_, new_n33211_, new_n33212_, new_n33213_,
    new_n33214_, new_n33215_, new_n33216_, new_n33217_, new_n33218_,
    new_n33219_, new_n33220_, new_n33221_, new_n33222_, new_n33223_,
    new_n33224_, new_n33225_, new_n33226_, new_n33227_, new_n33228_,
    new_n33229_, new_n33230_, new_n33231_, new_n33232_, new_n33233_,
    new_n33234_, new_n33235_, new_n33236_, new_n33237_, new_n33238_,
    new_n33239_, new_n33240_, new_n33241_, new_n33242_, new_n33243_,
    new_n33244_, new_n33245_, new_n33246_, new_n33247_, new_n33248_,
    new_n33249_, new_n33250_, new_n33251_, new_n33252_, new_n33253_,
    new_n33254_, new_n33255_, new_n33256_, new_n33257_, new_n33258_,
    new_n33259_, new_n33260_, new_n33261_, new_n33262_, new_n33263_,
    new_n33264_, new_n33265_, new_n33266_, new_n33267_, new_n33268_,
    new_n33269_, new_n33270_, new_n33271_, new_n33272_, new_n33273_,
    new_n33274_, new_n33275_, new_n33276_, new_n33277_, new_n33278_,
    new_n33279_, new_n33280_, new_n33281_, new_n33282_, new_n33283_,
    new_n33284_, new_n33285_, new_n33286_, new_n33287_, new_n33288_,
    new_n33289_, new_n33290_, new_n33291_, new_n33292_, new_n33293_,
    new_n33294_, new_n33295_, new_n33296_, new_n33297_, new_n33298_,
    new_n33299_, new_n33300_, new_n33301_, new_n33302_, new_n33303_,
    new_n33304_, new_n33305_, new_n33306_, new_n33307_, new_n33308_,
    new_n33309_, new_n33310_, new_n33311_, new_n33312_, new_n33313_,
    new_n33314_, new_n33315_, new_n33316_, new_n33317_, new_n33318_,
    new_n33319_, new_n33320_, new_n33321_, new_n33322_, new_n33323_,
    new_n33324_, new_n33325_, new_n33326_, new_n33327_, new_n33328_,
    new_n33329_, new_n33330_, new_n33331_, new_n33332_, new_n33333_,
    new_n33334_, new_n33335_, new_n33336_, new_n33337_, new_n33338_,
    new_n33339_, new_n33340_, new_n33341_, new_n33342_, new_n33343_,
    new_n33344_, new_n33345_, new_n33346_, new_n33347_, new_n33348_,
    new_n33349_, new_n33350_, new_n33351_, new_n33352_, new_n33353_,
    new_n33354_, new_n33355_, new_n33356_, new_n33357_, new_n33358_,
    new_n33359_, new_n33360_, new_n33361_, new_n33362_, new_n33363_,
    new_n33364_, new_n33365_, new_n33366_, new_n33367_, new_n33368_,
    new_n33369_, new_n33370_, new_n33371_, new_n33372_, new_n33373_,
    new_n33374_, new_n33375_, new_n33376_, new_n33377_, new_n33378_,
    new_n33379_, new_n33380_, new_n33381_, new_n33382_, new_n33383_,
    new_n33384_, new_n33385_, new_n33386_, new_n33387_, new_n33388_,
    new_n33389_, new_n33390_, new_n33391_, new_n33392_, new_n33393_,
    new_n33394_, new_n33395_, new_n33396_, new_n33397_, new_n33398_,
    new_n33399_, new_n33400_, new_n33401_, new_n33402_, new_n33403_,
    new_n33404_, new_n33405_, new_n33406_, new_n33407_, new_n33408_,
    new_n33409_, new_n33410_, new_n33411_, new_n33412_, new_n33413_,
    new_n33414_, new_n33415_, new_n33416_, new_n33417_, new_n33418_,
    new_n33419_, new_n33420_, new_n33421_, new_n33422_, new_n33423_,
    new_n33424_, new_n33425_, new_n33426_, new_n33427_, new_n33428_,
    new_n33429_, new_n33430_, new_n33431_, new_n33432_, new_n33433_,
    new_n33434_, new_n33435_, new_n33436_, new_n33437_, new_n33438_,
    new_n33439_, new_n33440_, new_n33441_, new_n33442_, new_n33443_,
    new_n33444_, new_n33445_, new_n33446_, new_n33447_, new_n33448_,
    new_n33449_, new_n33450_, new_n33451_, new_n33452_, new_n33453_,
    new_n33454_, new_n33455_, new_n33456_, new_n33457_, new_n33458_,
    new_n33459_, new_n33460_, new_n33461_, new_n33462_, new_n33463_,
    new_n33464_, new_n33465_, new_n33466_, new_n33467_, new_n33468_,
    new_n33469_, new_n33470_, new_n33471_, new_n33472_, new_n33473_,
    new_n33474_, new_n33475_, new_n33476_, new_n33477_, new_n33478_,
    new_n33479_, new_n33480_, new_n33481_, new_n33482_, new_n33483_,
    new_n33484_, new_n33485_, new_n33486_, new_n33487_, new_n33488_,
    new_n33489_, new_n33490_, new_n33491_, new_n33492_, new_n33493_,
    new_n33494_, new_n33495_, new_n33496_, new_n33497_, new_n33498_,
    new_n33499_, new_n33500_, new_n33501_, new_n33502_, new_n33503_,
    new_n33504_, new_n33505_, new_n33506_, new_n33507_, new_n33508_,
    new_n33509_, new_n33510_, new_n33511_, new_n33512_, new_n33513_,
    new_n33514_, new_n33515_, new_n33516_, new_n33517_, new_n33518_,
    new_n33519_, new_n33520_, new_n33521_, new_n33522_, new_n33523_,
    new_n33524_, new_n33525_, new_n33526_, new_n33527_, new_n33528_,
    new_n33529_, new_n33530_, new_n33531_, new_n33532_, new_n33533_,
    new_n33534_, new_n33535_, new_n33536_, new_n33537_, new_n33538_,
    new_n33539_, new_n33540_, new_n33541_, new_n33542_, new_n33543_,
    new_n33544_, new_n33545_, new_n33546_, new_n33547_, new_n33548_,
    new_n33549_, new_n33550_, new_n33551_, new_n33552_, new_n33553_,
    new_n33554_, new_n33555_, new_n33556_, new_n33557_, new_n33558_,
    new_n33559_, new_n33560_, new_n33561_, new_n33562_, new_n33563_,
    new_n33564_, new_n33565_, new_n33566_, new_n33567_, new_n33568_,
    new_n33569_, new_n33570_, new_n33571_, new_n33572_, new_n33573_,
    new_n33574_, new_n33575_, new_n33576_, new_n33577_, new_n33578_,
    new_n33579_, new_n33580_, new_n33581_, new_n33582_, new_n33583_,
    new_n33584_, new_n33585_, new_n33586_, new_n33587_, new_n33588_,
    new_n33589_, new_n33590_, new_n33591_, new_n33592_, new_n33593_,
    new_n33594_, new_n33595_, new_n33596_, new_n33597_, new_n33598_,
    new_n33599_, new_n33600_, new_n33601_, new_n33602_, new_n33603_,
    new_n33604_, new_n33605_, new_n33606_, new_n33607_, new_n33608_,
    new_n33609_, new_n33610_, new_n33611_, new_n33612_, new_n33613_,
    new_n33614_, new_n33615_, new_n33616_, new_n33617_, new_n33618_,
    new_n33619_, new_n33620_, new_n33621_, new_n33622_, new_n33623_,
    new_n33624_, new_n33625_, new_n33626_, new_n33627_, new_n33628_,
    new_n33629_, new_n33630_, new_n33631_, new_n33632_, new_n33633_,
    new_n33634_, new_n33635_, new_n33636_, new_n33637_, new_n33638_,
    new_n33639_, new_n33640_, new_n33641_, new_n33642_, new_n33643_,
    new_n33644_, new_n33645_, new_n33646_, new_n33647_, new_n33648_,
    new_n33649_, new_n33650_, new_n33651_, new_n33652_, new_n33653_,
    new_n33654_, new_n33655_, new_n33656_, new_n33657_, new_n33658_,
    new_n33659_, new_n33660_, new_n33661_, new_n33662_, new_n33663_,
    new_n33664_, new_n33665_, new_n33666_, new_n33667_, new_n33668_,
    new_n33669_, new_n33670_, new_n33671_, new_n33672_, new_n33673_,
    new_n33674_, new_n33675_, new_n33676_, new_n33677_, new_n33678_,
    new_n33679_, new_n33680_, new_n33681_, new_n33682_, new_n33683_,
    new_n33684_, new_n33685_, new_n33686_, new_n33687_, new_n33688_,
    new_n33689_, new_n33690_, new_n33691_, new_n33692_, new_n33693_,
    new_n33694_, new_n33695_, new_n33696_, new_n33697_, new_n33698_,
    new_n33699_, new_n33700_, new_n33701_, new_n33702_, new_n33703_,
    new_n33704_, new_n33705_, new_n33706_, new_n33707_, new_n33708_,
    new_n33709_, new_n33710_, new_n33711_, new_n33712_, new_n33713_,
    new_n33714_, new_n33715_, new_n33716_, new_n33717_, new_n33718_,
    new_n33719_, new_n33720_, new_n33721_, new_n33722_, new_n33723_,
    new_n33724_, new_n33725_, new_n33726_, new_n33727_, new_n33728_,
    new_n33729_, new_n33730_, new_n33731_, new_n33732_, new_n33733_,
    new_n33734_, new_n33735_, new_n33736_, new_n33737_, new_n33738_,
    new_n33739_, new_n33740_, new_n33741_, new_n33742_, new_n33743_,
    new_n33744_, new_n33745_, new_n33746_, new_n33747_, new_n33748_,
    new_n33749_, new_n33750_, new_n33751_, new_n33752_, new_n33753_,
    new_n33754_, new_n33755_, new_n33756_, new_n33757_, new_n33758_,
    new_n33759_, new_n33760_, new_n33761_, new_n33762_, new_n33763_,
    new_n33764_, new_n33765_, new_n33766_, new_n33767_, new_n33768_,
    new_n33769_, new_n33770_, new_n33771_, new_n33772_, new_n33773_,
    new_n33774_, new_n33775_, new_n33776_, new_n33777_, new_n33778_,
    new_n33779_, new_n33780_, new_n33781_, new_n33782_, new_n33783_,
    new_n33784_, new_n33785_, new_n33786_, new_n33787_, new_n33788_,
    new_n33789_, new_n33790_, new_n33791_, new_n33792_, new_n33793_,
    new_n33794_, new_n33795_, new_n33796_, new_n33797_, new_n33798_,
    new_n33799_, new_n33800_, new_n33801_, new_n33802_, new_n33803_,
    new_n33804_, new_n33805_, new_n33806_, new_n33807_, new_n33808_,
    new_n33809_, new_n33810_, new_n33811_, new_n33812_, new_n33813_,
    new_n33814_, new_n33815_, new_n33816_, new_n33817_, new_n33818_,
    new_n33819_, new_n33820_, new_n33821_, new_n33822_, new_n33823_,
    new_n33824_, new_n33825_, new_n33826_, new_n33827_, new_n33828_,
    new_n33829_, new_n33830_, new_n33831_, new_n33832_, new_n33833_,
    new_n33834_, new_n33835_, new_n33836_, new_n33837_, new_n33838_,
    new_n33839_, new_n33840_, new_n33841_, new_n33842_, new_n33843_,
    new_n33844_, new_n33845_, new_n33846_, new_n33847_, new_n33848_,
    new_n33849_, new_n33850_, new_n33851_, new_n33852_, new_n33853_,
    new_n33854_, new_n33855_, new_n33856_, new_n33857_, new_n33858_,
    new_n33859_, new_n33860_, new_n33861_, new_n33862_, new_n33863_,
    new_n33864_, new_n33865_, new_n33866_, new_n33867_, new_n33868_,
    new_n33869_, new_n33870_, new_n33871_, new_n33872_, new_n33873_,
    new_n33874_, new_n33875_, new_n33876_, new_n33877_, new_n33878_,
    new_n33879_, new_n33880_, new_n33881_, new_n33882_, new_n33883_,
    new_n33884_, new_n33885_, new_n33886_, new_n33887_, new_n33888_,
    new_n33889_, new_n33890_, new_n33891_, new_n33892_, new_n33893_,
    new_n33894_, new_n33895_, new_n33896_, new_n33897_, new_n33898_,
    new_n33899_, new_n33900_, new_n33901_, new_n33902_, new_n33903_,
    new_n33904_, new_n33905_, new_n33906_, new_n33907_, new_n33908_,
    new_n33909_, new_n33910_, new_n33911_, new_n33912_, new_n33913_,
    new_n33914_, new_n33915_, new_n33916_, new_n33917_, new_n33918_,
    new_n33919_, new_n33920_, new_n33921_, new_n33922_, new_n33923_,
    new_n33924_, new_n33925_, new_n33926_, new_n33927_, new_n33928_,
    new_n33929_, new_n33930_, new_n33931_, new_n33932_, new_n33933_,
    new_n33934_, new_n33935_, new_n33936_, new_n33937_, new_n33938_,
    new_n33939_, new_n33940_, new_n33941_, new_n33942_, new_n33943_,
    new_n33944_, new_n33945_, new_n33946_, new_n33947_, new_n33948_,
    new_n33949_, new_n33950_, new_n33951_, new_n33952_, new_n33953_,
    new_n33954_, new_n33955_, new_n33956_, new_n33957_, new_n33958_,
    new_n33959_, new_n33960_, new_n33961_, new_n33962_, new_n33963_,
    new_n33964_, new_n33965_, new_n33966_, new_n33967_, new_n33968_,
    new_n33969_, new_n33970_, new_n33971_, new_n33972_, new_n33973_,
    new_n33974_, new_n33975_, new_n33976_, new_n33977_, new_n33978_,
    new_n33979_, new_n33980_, new_n33981_, new_n33982_, new_n33983_,
    new_n33984_, new_n33985_, new_n33986_, new_n33987_, new_n33988_,
    new_n33989_, new_n33990_, new_n33991_, new_n33992_, new_n33993_,
    new_n33994_, new_n33995_, new_n33996_, new_n33997_, new_n33998_,
    new_n33999_, new_n34000_, new_n34001_, new_n34002_, new_n34003_,
    new_n34004_, new_n34005_, new_n34006_, new_n34007_, new_n34008_,
    new_n34009_, new_n34010_, new_n34011_, new_n34012_, new_n34013_,
    new_n34014_, new_n34015_, new_n34016_, new_n34017_, new_n34018_,
    new_n34019_, new_n34020_, new_n34021_, new_n34022_, new_n34023_,
    new_n34024_, new_n34025_, new_n34026_, new_n34027_, new_n34028_,
    new_n34029_, new_n34030_, new_n34031_, new_n34032_, new_n34033_,
    new_n34034_, new_n34035_, new_n34036_, new_n34037_, new_n34038_,
    new_n34039_, new_n34040_, new_n34041_, new_n34042_, new_n34043_,
    new_n34044_, new_n34045_, new_n34046_, new_n34047_, new_n34048_,
    new_n34049_, new_n34050_, new_n34051_, new_n34052_, new_n34053_,
    new_n34054_, new_n34055_, new_n34056_, new_n34057_, new_n34058_,
    new_n34059_, new_n34060_, new_n34061_, new_n34062_, new_n34063_,
    new_n34064_, new_n34065_, new_n34066_, new_n34067_, new_n34068_,
    new_n34069_, new_n34070_, new_n34071_, new_n34072_, new_n34073_,
    new_n34074_, new_n34075_, new_n34076_, new_n34077_, new_n34078_,
    new_n34079_, new_n34080_, new_n34081_, new_n34082_, new_n34083_,
    new_n34084_, new_n34085_, new_n34086_, new_n34087_, new_n34088_,
    new_n34089_, new_n34090_, new_n34091_, new_n34092_, new_n34093_,
    new_n34094_, new_n34095_, new_n34096_, new_n34097_, new_n34098_,
    new_n34099_, new_n34100_, new_n34101_, new_n34102_, new_n34103_,
    new_n34104_, new_n34105_, new_n34106_, new_n34107_, new_n34108_,
    new_n34109_, new_n34110_, new_n34111_, new_n34112_, new_n34113_,
    new_n34114_, new_n34115_, new_n34116_, new_n34117_, new_n34118_,
    new_n34119_, new_n34120_, new_n34121_, new_n34122_, new_n34123_,
    new_n34124_, new_n34125_, new_n34126_, new_n34127_, new_n34128_,
    new_n34129_, new_n34130_, new_n34131_, new_n34132_, new_n34133_,
    new_n34134_, new_n34135_, new_n34136_, new_n34137_, new_n34138_,
    new_n34139_, new_n34140_, new_n34141_, new_n34142_, new_n34143_,
    new_n34144_, new_n34145_, new_n34146_, new_n34147_, new_n34148_,
    new_n34149_, new_n34150_, new_n34151_, new_n34152_, new_n34153_,
    new_n34154_, new_n34155_, new_n34156_, new_n34157_, new_n34158_,
    new_n34159_, new_n34160_, new_n34161_, new_n34162_, new_n34163_,
    new_n34164_, new_n34165_, new_n34166_, new_n34167_, new_n34168_,
    new_n34169_, new_n34170_, new_n34171_, new_n34172_, new_n34173_,
    new_n34174_, new_n34175_, new_n34176_, new_n34177_, new_n34178_,
    new_n34179_, new_n34180_, new_n34181_, new_n34182_, new_n34183_,
    new_n34184_, new_n34185_, new_n34186_, new_n34187_, new_n34188_,
    new_n34189_, new_n34190_, new_n34191_, new_n34192_, new_n34193_,
    new_n34194_, new_n34195_, new_n34196_, new_n34197_, new_n34198_,
    new_n34199_, new_n34200_, new_n34201_, new_n34202_, new_n34203_,
    new_n34204_, new_n34205_, new_n34206_, new_n34207_, new_n34208_,
    new_n34209_, new_n34210_, new_n34211_, new_n34212_, new_n34213_,
    new_n34214_, new_n34215_, new_n34216_, new_n34217_, new_n34218_,
    new_n34219_, new_n34220_, new_n34221_, new_n34222_, new_n34223_,
    new_n34224_, new_n34225_, new_n34226_, new_n34227_, new_n34228_,
    new_n34229_, new_n34230_, new_n34231_, new_n34232_, new_n34233_,
    new_n34234_, new_n34235_, new_n34236_, new_n34237_, new_n34238_,
    new_n34239_, new_n34240_, new_n34241_, new_n34242_, new_n34243_,
    new_n34244_, new_n34245_, new_n34246_, new_n34247_, new_n34248_,
    new_n34249_, new_n34250_, new_n34251_, new_n34252_, new_n34253_,
    new_n34254_, new_n34255_, new_n34256_, new_n34257_, new_n34258_,
    new_n34259_, new_n34260_, new_n34261_, new_n34262_, new_n34263_,
    new_n34264_, new_n34265_, new_n34266_, new_n34267_, new_n34268_,
    new_n34269_, new_n34270_, new_n34271_, new_n34272_, new_n34273_,
    new_n34274_, new_n34275_, new_n34276_, new_n34277_, new_n34278_,
    new_n34279_, new_n34280_, new_n34281_, new_n34282_, new_n34283_,
    new_n34284_, new_n34285_, new_n34286_, new_n34287_, new_n34288_,
    new_n34289_, new_n34290_, new_n34291_, new_n34292_, new_n34293_,
    new_n34294_, new_n34295_, new_n34296_, new_n34297_, new_n34298_,
    new_n34299_, new_n34300_, new_n34301_, new_n34302_, new_n34303_,
    new_n34304_, new_n34305_, new_n34306_, new_n34307_, new_n34308_,
    new_n34309_, new_n34310_, new_n34311_, new_n34312_, new_n34313_,
    new_n34314_, new_n34315_, new_n34316_, new_n34317_, new_n34318_,
    new_n34319_, new_n34320_, new_n34321_, new_n34322_, new_n34323_,
    new_n34324_, new_n34325_, new_n34326_, new_n34327_, new_n34328_,
    new_n34329_, new_n34330_, new_n34331_, new_n34332_, new_n34333_,
    new_n34334_, new_n34335_, new_n34336_, new_n34337_, new_n34338_,
    new_n34339_, new_n34340_, new_n34341_, new_n34342_, new_n34343_,
    new_n34344_, new_n34345_, new_n34346_, new_n34347_, new_n34348_,
    new_n34349_, new_n34350_, new_n34351_, new_n34352_, new_n34353_,
    new_n34354_, new_n34355_, new_n34356_, new_n34357_, new_n34358_,
    new_n34359_, new_n34360_, new_n34361_, new_n34362_, new_n34363_,
    new_n34364_, new_n34365_, new_n34366_, new_n34367_, new_n34368_,
    new_n34369_, new_n34370_, new_n34371_, new_n34372_, new_n34373_,
    new_n34374_, new_n34375_, new_n34376_, new_n34377_, new_n34378_,
    new_n34379_, new_n34380_, new_n34381_, new_n34382_, new_n34383_,
    new_n34384_, new_n34385_, new_n34386_, new_n34387_, new_n34388_,
    new_n34389_, new_n34390_, new_n34391_, new_n34392_, new_n34393_,
    new_n34394_, new_n34395_, new_n34396_, new_n34397_, new_n34398_,
    new_n34399_, new_n34400_, new_n34401_, new_n34402_, new_n34403_,
    new_n34404_, new_n34405_, new_n34406_, new_n34407_, new_n34408_,
    new_n34409_, new_n34410_, new_n34411_, new_n34412_, new_n34413_,
    new_n34414_, new_n34415_, new_n34416_, new_n34417_, new_n34418_,
    new_n34419_, new_n34420_, new_n34421_, new_n34422_, new_n34423_,
    new_n34424_, new_n34425_, new_n34426_, new_n34427_, new_n34428_,
    new_n34429_, new_n34430_, new_n34431_, new_n34432_, new_n34433_,
    new_n34434_, new_n34435_, new_n34436_, new_n34437_, new_n34438_,
    new_n34439_, new_n34440_, new_n34441_, new_n34442_, new_n34443_,
    new_n34444_, new_n34445_, new_n34446_, new_n34447_, new_n34448_,
    new_n34449_, new_n34450_, new_n34451_, new_n34452_, new_n34453_,
    new_n34454_, new_n34455_, new_n34456_, new_n34457_, new_n34458_,
    new_n34459_, new_n34460_, new_n34461_, new_n34462_, new_n34463_,
    new_n34464_, new_n34465_, new_n34466_, new_n34467_, new_n34468_,
    new_n34469_, new_n34470_, new_n34471_, new_n34472_, new_n34473_,
    new_n34474_, new_n34475_, new_n34476_, new_n34477_, new_n34478_,
    new_n34479_, new_n34480_, new_n34481_, new_n34482_, new_n34483_,
    new_n34484_, new_n34485_, new_n34486_, new_n34487_, new_n34488_,
    new_n34489_, new_n34490_, new_n34491_, new_n34492_, new_n34493_,
    new_n34494_, new_n34495_, new_n34496_, new_n34497_, new_n34498_,
    new_n34499_, new_n34500_, new_n34501_, new_n34502_, new_n34503_,
    new_n34504_, new_n34505_, new_n34506_, new_n34507_, new_n34508_,
    new_n34509_, new_n34510_, new_n34511_, new_n34512_, new_n34513_,
    new_n34514_, new_n34515_, new_n34516_, new_n34517_, new_n34518_,
    new_n34519_, new_n34520_, new_n34521_, new_n34522_, new_n34523_,
    new_n34524_, new_n34525_, new_n34526_, new_n34527_, new_n34528_,
    new_n34529_, new_n34530_, new_n34531_, new_n34532_, new_n34533_,
    new_n34534_, new_n34535_, new_n34536_, new_n34537_, new_n34538_,
    new_n34539_, new_n34540_, new_n34541_, new_n34542_, new_n34543_,
    new_n34544_, new_n34545_, new_n34546_, new_n34547_, new_n34548_,
    new_n34549_, new_n34550_, new_n34551_, new_n34552_, new_n34553_,
    new_n34554_, new_n34555_, new_n34556_, new_n34557_, new_n34558_,
    new_n34559_, new_n34560_, new_n34561_, new_n34562_, new_n34563_,
    new_n34564_, new_n34565_, new_n34566_, new_n34567_, new_n34568_,
    new_n34569_, new_n34570_, new_n34571_, new_n34572_, new_n34573_,
    new_n34574_, new_n34575_, new_n34576_, new_n34577_, new_n34578_,
    new_n34579_, new_n34580_, new_n34581_, new_n34582_, new_n34583_,
    new_n34584_, new_n34585_, new_n34586_, new_n34587_, new_n34588_,
    new_n34589_, new_n34590_, new_n34591_, new_n34592_, new_n34593_,
    new_n34594_, new_n34595_, new_n34596_, new_n34597_, new_n34598_,
    new_n34599_, new_n34600_, new_n34601_, new_n34602_, new_n34603_,
    new_n34604_, new_n34605_, new_n34606_, new_n34607_, new_n34608_,
    new_n34609_, new_n34610_, new_n34611_, new_n34612_, new_n34613_,
    new_n34614_, new_n34615_, new_n34616_, new_n34617_, new_n34618_,
    new_n34619_, new_n34620_, new_n34621_, new_n34622_, new_n34623_,
    new_n34624_, new_n34625_, new_n34626_, new_n34627_, new_n34628_,
    new_n34629_, new_n34630_, new_n34631_, new_n34632_, new_n34633_,
    new_n34634_, new_n34635_, new_n34636_, new_n34637_, new_n34638_,
    new_n34639_, new_n34640_, new_n34641_, new_n34642_, new_n34643_,
    new_n34644_, new_n34645_, new_n34646_, new_n34647_, new_n34648_,
    new_n34649_, new_n34650_, new_n34651_, new_n34652_, new_n34653_,
    new_n34654_, new_n34655_, new_n34656_, new_n34657_, new_n34658_,
    new_n34659_, new_n34660_, new_n34661_, new_n34662_, new_n34663_,
    new_n34664_, new_n34665_, new_n34666_, new_n34667_, new_n34668_,
    new_n34669_, new_n34670_, new_n34671_, new_n34672_, new_n34673_,
    new_n34674_, new_n34675_, new_n34676_, new_n34677_, new_n34678_,
    new_n34679_, new_n34680_, new_n34681_, new_n34682_, new_n34683_,
    new_n34684_, new_n34685_, new_n34686_, new_n34687_, new_n34688_,
    new_n34689_, new_n34690_, new_n34691_, new_n34692_, new_n34693_,
    new_n34694_, new_n34695_, new_n34696_, new_n34697_, new_n34698_,
    new_n34699_, new_n34700_, new_n34701_, new_n34702_, new_n34703_,
    new_n34704_, new_n34705_, new_n34706_, new_n34707_, new_n34708_,
    new_n34709_, new_n34710_, new_n34711_, new_n34712_, new_n34713_,
    new_n34714_, new_n34715_, new_n34716_, new_n34717_, new_n34718_,
    new_n34719_, new_n34720_, new_n34721_, new_n34722_, new_n34723_,
    new_n34724_, new_n34725_, new_n34726_, new_n34727_, new_n34728_,
    new_n34729_, new_n34730_, new_n34731_, new_n34732_, new_n34733_,
    new_n34734_, new_n34735_, new_n34736_, new_n34737_, new_n34738_,
    new_n34739_, new_n34740_, new_n34741_, new_n34742_, new_n34743_,
    new_n34744_, new_n34745_, new_n34746_, new_n34747_, new_n34748_,
    new_n34749_, new_n34750_, new_n34751_, new_n34752_, new_n34753_,
    new_n34754_, new_n34755_, new_n34756_, new_n34757_, new_n34758_,
    new_n34759_, new_n34760_, new_n34761_, new_n34762_, new_n34763_,
    new_n34764_, new_n34765_, new_n34766_, new_n34767_, new_n34768_,
    new_n34769_, new_n34770_, new_n34771_, new_n34772_, new_n34773_,
    new_n34774_, new_n34775_, new_n34776_, new_n34777_, new_n34778_,
    new_n34779_, new_n34780_, new_n34781_, new_n34782_, new_n34783_,
    new_n34784_, new_n34785_, new_n34786_, new_n34787_, new_n34788_,
    new_n34789_, new_n34790_, new_n34791_, new_n34792_, new_n34793_,
    new_n34794_, new_n34795_, new_n34796_, new_n34797_, new_n34798_,
    new_n34799_, new_n34800_, new_n34801_, new_n34802_, new_n34803_,
    new_n34804_, new_n34805_, new_n34806_, new_n34807_, new_n34808_,
    new_n34809_, new_n34810_, new_n34811_, new_n34812_, new_n34813_,
    new_n34814_, new_n34815_, new_n34816_, new_n34817_, new_n34818_,
    new_n34819_, new_n34820_, new_n34821_, new_n34822_, new_n34823_,
    new_n34824_, new_n34825_, new_n34826_, new_n34827_, new_n34828_,
    new_n34829_, new_n34830_, new_n34831_, new_n34832_, new_n34833_,
    new_n34834_, new_n34835_, new_n34836_, new_n34837_, new_n34838_,
    new_n34839_, new_n34840_, new_n34841_, new_n34842_, new_n34843_,
    new_n34844_, new_n34845_, new_n34846_, new_n34847_, new_n34848_,
    new_n34849_, new_n34850_, new_n34851_, new_n34852_, new_n34853_,
    new_n34854_, new_n34855_, new_n34856_, new_n34857_, new_n34858_,
    new_n34859_, new_n34860_, new_n34861_, new_n34862_, new_n34863_,
    new_n34864_, new_n34865_, new_n34866_, new_n34867_, new_n34868_,
    new_n34869_, new_n34870_, new_n34871_, new_n34872_, new_n34873_,
    new_n34874_, new_n34875_, new_n34876_, new_n34877_, new_n34878_,
    new_n34879_, new_n34880_, new_n34881_, new_n34882_, new_n34883_,
    new_n34884_, new_n34885_, new_n34886_, new_n34887_, new_n34888_,
    new_n34889_, new_n34890_, new_n34891_, new_n34892_, new_n34893_,
    new_n34894_, new_n34895_, new_n34896_, new_n34897_, new_n34898_,
    new_n34899_, new_n34900_, new_n34901_, new_n34902_, new_n34903_,
    new_n34904_, new_n34905_, new_n34906_, new_n34907_, new_n34908_,
    new_n34909_, new_n34910_, new_n34911_, new_n34912_, new_n34913_,
    new_n34914_, new_n34915_, new_n34916_, new_n34917_, new_n34918_,
    new_n34919_, new_n34920_, new_n34921_, new_n34922_, new_n34923_,
    new_n34924_, new_n34925_, new_n34926_, new_n34927_, new_n34928_,
    new_n34929_, new_n34930_, new_n34931_, new_n34932_, new_n34933_,
    new_n34934_, new_n34935_, new_n34936_, new_n34937_, new_n34938_,
    new_n34939_, new_n34940_, new_n34941_, new_n34942_, new_n34943_,
    new_n34944_, new_n34945_, new_n34946_, new_n34947_, new_n34948_,
    new_n34949_, new_n34950_, new_n34951_, new_n34952_, new_n34953_,
    new_n34954_, new_n34955_, new_n34956_, new_n34957_, new_n34958_,
    new_n34959_, new_n34960_, new_n34961_, new_n34962_, new_n34963_,
    new_n34964_, new_n34965_, new_n34966_, new_n34967_, new_n34968_,
    new_n34969_, new_n34970_, new_n34971_, new_n34972_, new_n34973_,
    new_n34974_, new_n34975_, new_n34976_, new_n34977_, new_n34978_,
    new_n34979_, new_n34980_, new_n34981_, new_n34982_, new_n34983_,
    new_n34984_, new_n34985_, new_n34986_, new_n34987_, new_n34988_,
    new_n34989_, new_n34990_, new_n34991_, new_n34992_, new_n34993_,
    new_n34994_, new_n34995_, new_n34996_, new_n34997_, new_n34998_,
    new_n34999_, new_n35000_, new_n35001_, new_n35002_, new_n35003_,
    new_n35004_, new_n35005_, new_n35006_, new_n35007_, new_n35008_,
    new_n35009_, new_n35010_, new_n35011_, new_n35012_, new_n35013_,
    new_n35014_, new_n35015_, new_n35016_, new_n35017_, new_n35018_,
    new_n35019_, new_n35020_, new_n35021_, new_n35022_, new_n35023_,
    new_n35024_, new_n35025_, new_n35026_, new_n35027_, new_n35028_,
    new_n35029_, new_n35030_, new_n35031_, new_n35032_, new_n35033_,
    new_n35034_, new_n35035_, new_n35036_, new_n35037_, new_n35038_,
    new_n35039_, new_n35040_, new_n35041_, new_n35042_, new_n35043_,
    new_n35044_, new_n35045_, new_n35046_, new_n35047_, new_n35048_,
    new_n35049_, new_n35050_, new_n35051_, new_n35052_, new_n35053_,
    new_n35054_, new_n35055_, new_n35056_, new_n35057_, new_n35058_,
    new_n35059_, new_n35060_, new_n35061_, new_n35062_, new_n35063_,
    new_n35064_, new_n35065_, new_n35066_, new_n35067_, new_n35068_,
    new_n35069_, new_n35070_, new_n35071_, new_n35072_, new_n35073_,
    new_n35074_, new_n35075_, new_n35076_, new_n35077_, new_n35078_,
    new_n35079_, new_n35080_, new_n35081_, new_n35082_, new_n35083_,
    new_n35084_, new_n35085_, new_n35086_, new_n35087_, new_n35088_,
    new_n35089_, new_n35090_, new_n35091_, new_n35092_, new_n35093_,
    new_n35094_, new_n35095_, new_n35096_, new_n35097_, new_n35098_,
    new_n35099_, new_n35100_, new_n35101_, new_n35102_, new_n35103_,
    new_n35104_, new_n35105_, new_n35106_, new_n35107_, new_n35108_,
    new_n35109_, new_n35110_, new_n35111_, new_n35112_, new_n35113_,
    new_n35114_, new_n35115_, new_n35116_, new_n35117_, new_n35118_,
    new_n35119_, new_n35120_, new_n35121_, new_n35122_, new_n35123_,
    new_n35124_, new_n35125_, new_n35126_, new_n35127_, new_n35128_,
    new_n35129_, new_n35130_, new_n35131_, new_n35132_, new_n35133_,
    new_n35134_, new_n35135_, new_n35136_, new_n35137_, new_n35138_,
    new_n35139_, new_n35140_, new_n35141_, new_n35142_, new_n35143_,
    new_n35144_, new_n35145_, new_n35146_, new_n35147_, new_n35148_,
    new_n35149_, new_n35150_, new_n35151_, new_n35152_, new_n35153_,
    new_n35154_, new_n35155_, new_n35156_, new_n35157_, new_n35158_,
    new_n35159_, new_n35160_, new_n35161_, new_n35162_, new_n35163_,
    new_n35164_, new_n35165_, new_n35166_, new_n35167_, new_n35168_,
    new_n35169_, new_n35170_, new_n35171_, new_n35172_, new_n35173_,
    new_n35174_, new_n35175_, new_n35176_, new_n35177_, new_n35178_,
    new_n35179_, new_n35180_, new_n35181_, new_n35182_, new_n35183_,
    new_n35184_, new_n35185_, new_n35186_, new_n35187_, new_n35188_,
    new_n35189_, new_n35190_, new_n35191_, new_n35192_, new_n35193_,
    new_n35194_, new_n35195_, new_n35196_, new_n35197_, new_n35198_,
    new_n35199_, new_n35200_, new_n35201_, new_n35202_, new_n35203_,
    new_n35204_, new_n35205_, new_n35206_, new_n35207_, new_n35208_,
    new_n35209_, new_n35210_, new_n35211_, new_n35212_, new_n35213_,
    new_n35214_, new_n35215_, new_n35216_, new_n35217_, new_n35218_,
    new_n35219_, new_n35220_, new_n35221_, new_n35222_, new_n35223_,
    new_n35224_, new_n35225_, new_n35226_, new_n35227_, new_n35228_,
    new_n35229_, new_n35230_, new_n35231_, new_n35232_, new_n35233_,
    new_n35234_, new_n35235_, new_n35236_, new_n35237_, new_n35238_,
    new_n35239_, new_n35240_, new_n35241_, new_n35242_, new_n35243_,
    new_n35244_, new_n35245_, new_n35246_, new_n35247_, new_n35248_,
    new_n35249_, new_n35250_, new_n35251_, new_n35252_, new_n35253_,
    new_n35254_, new_n35255_, new_n35256_, new_n35257_, new_n35258_,
    new_n35259_, new_n35260_, new_n35261_, new_n35262_, new_n35263_,
    new_n35264_, new_n35265_, new_n35266_, new_n35267_, new_n35268_,
    new_n35269_, new_n35270_, new_n35271_, new_n35272_, new_n35273_,
    new_n35274_, new_n35275_, new_n35276_, new_n35277_, new_n35278_,
    new_n35279_, new_n35280_, new_n35281_, new_n35282_, new_n35283_,
    new_n35284_, new_n35285_, new_n35286_, new_n35287_, new_n35288_,
    new_n35289_, new_n35290_, new_n35291_, new_n35292_, new_n35293_,
    new_n35294_, new_n35295_, new_n35296_, new_n35297_, new_n35298_,
    new_n35299_, new_n35300_, new_n35301_, new_n35302_, new_n35303_,
    new_n35304_, new_n35305_, new_n35306_, new_n35307_, new_n35308_,
    new_n35309_, new_n35310_, new_n35311_, new_n35312_, new_n35313_,
    new_n35314_, new_n35315_, new_n35316_, new_n35317_, new_n35318_,
    new_n35319_, new_n35320_, new_n35321_, new_n35322_, new_n35323_,
    new_n35324_, new_n35325_, new_n35326_, new_n35327_, new_n35328_,
    new_n35329_, new_n35330_, new_n35331_, new_n35332_, new_n35333_,
    new_n35334_, new_n35335_, new_n35336_, new_n35337_, new_n35338_,
    new_n35339_, new_n35340_, new_n35341_, new_n35342_, new_n35343_,
    new_n35344_, new_n35345_, new_n35346_, new_n35347_, new_n35348_,
    new_n35349_, new_n35350_, new_n35351_, new_n35352_, new_n35353_,
    new_n35354_, new_n35355_, new_n35356_, new_n35357_, new_n35358_,
    new_n35359_, new_n35360_, new_n35361_, new_n35362_, new_n35363_,
    new_n35364_, new_n35365_, new_n35366_, new_n35367_, new_n35368_,
    new_n35369_, new_n35370_, new_n35371_, new_n35372_, new_n35373_,
    new_n35374_, new_n35375_, new_n35376_, new_n35377_, new_n35378_,
    new_n35379_, new_n35380_, new_n35381_, new_n35382_, new_n35383_,
    new_n35384_, new_n35385_, new_n35386_, new_n35387_, new_n35388_,
    new_n35389_, new_n35390_, new_n35391_, new_n35392_, new_n35393_,
    new_n35394_, new_n35395_, new_n35396_, new_n35397_, new_n35398_,
    new_n35399_, new_n35400_, new_n35401_, new_n35402_, new_n35403_,
    new_n35404_, new_n35405_, new_n35406_, new_n35407_, new_n35408_,
    new_n35409_, new_n35410_, new_n35411_, new_n35412_, new_n35413_,
    new_n35414_, new_n35415_, new_n35416_, new_n35417_, new_n35418_,
    new_n35419_, new_n35420_, new_n35421_, new_n35422_, new_n35423_,
    new_n35424_, new_n35425_, new_n35426_, new_n35427_, new_n35428_,
    new_n35429_, new_n35430_, new_n35431_, new_n35432_, new_n35433_,
    new_n35434_, new_n35435_, new_n35436_, new_n35437_, new_n35438_,
    new_n35439_, new_n35440_, new_n35441_, new_n35442_, new_n35443_,
    new_n35444_, new_n35445_, new_n35446_, new_n35447_, new_n35448_,
    new_n35449_, new_n35450_, new_n35451_, new_n35452_, new_n35453_,
    new_n35454_, new_n35455_, new_n35456_, new_n35457_, new_n35458_,
    new_n35459_, new_n35460_, new_n35461_, new_n35462_, new_n35463_,
    new_n35464_, new_n35465_, new_n35466_, new_n35467_, new_n35468_,
    new_n35469_, new_n35470_, new_n35471_, new_n35472_, new_n35473_,
    new_n35474_, new_n35475_, new_n35476_, new_n35477_, new_n35478_,
    new_n35479_, new_n35480_, new_n35481_, new_n35482_, new_n35483_,
    new_n35484_, new_n35485_, new_n35486_, new_n35487_, new_n35488_,
    new_n35489_, new_n35490_, new_n35491_, new_n35492_, new_n35493_,
    new_n35494_, new_n35495_, new_n35496_, new_n35497_, new_n35498_,
    new_n35499_, new_n35500_, new_n35501_, new_n35502_, new_n35503_,
    new_n35504_, new_n35505_, new_n35506_, new_n35507_, new_n35508_,
    new_n35509_, new_n35510_, new_n35511_, new_n35512_, new_n35513_,
    new_n35514_, new_n35515_, new_n35516_, new_n35517_, new_n35518_,
    new_n35519_, new_n35520_, new_n35521_, new_n35522_, new_n35523_,
    new_n35524_, new_n35525_, new_n35526_, new_n35527_, new_n35528_,
    new_n35529_, new_n35530_, new_n35531_, new_n35532_, new_n35533_,
    new_n35534_, new_n35535_, new_n35536_, new_n35537_, new_n35538_,
    new_n35539_, new_n35540_, new_n35541_, new_n35542_, new_n35543_,
    new_n35544_, new_n35545_, new_n35546_, new_n35547_, new_n35548_,
    new_n35549_, new_n35550_, new_n35551_, new_n35552_, new_n35553_,
    new_n35554_, new_n35555_, new_n35556_, new_n35557_, new_n35558_,
    new_n35559_, new_n35560_, new_n35561_, new_n35562_, new_n35563_,
    new_n35564_, new_n35565_, new_n35566_, new_n35567_, new_n35568_,
    new_n35569_, new_n35570_, new_n35571_, new_n35572_, new_n35573_,
    new_n35574_, new_n35575_, new_n35576_, new_n35577_, new_n35578_,
    new_n35579_, new_n35580_, new_n35581_, new_n35582_, new_n35583_,
    new_n35584_, new_n35585_, new_n35586_, new_n35587_, new_n35588_,
    new_n35589_, new_n35590_, new_n35591_, new_n35592_, new_n35593_,
    new_n35594_, new_n35595_, new_n35596_, new_n35597_, new_n35598_,
    new_n35599_, new_n35600_, new_n35601_, new_n35602_, new_n35603_,
    new_n35604_, new_n35605_, new_n35606_, new_n35607_, new_n35608_,
    new_n35609_, new_n35610_, new_n35611_, new_n35612_, new_n35613_,
    new_n35614_, new_n35615_, new_n35616_, new_n35617_, new_n35618_,
    new_n35619_, new_n35620_, new_n35621_, new_n35622_, new_n35623_,
    new_n35624_, new_n35625_, new_n35626_, new_n35627_, new_n35628_,
    new_n35629_, new_n35630_, new_n35631_, new_n35632_, new_n35633_,
    new_n35634_, new_n35635_, new_n35636_, new_n35637_, new_n35638_,
    new_n35639_, new_n35640_, new_n35641_, new_n35642_, new_n35643_,
    new_n35644_, new_n35645_, new_n35646_, new_n35647_, new_n35648_,
    new_n35649_, new_n35650_, new_n35651_, new_n35652_, new_n35653_,
    new_n35654_, new_n35655_, new_n35656_, new_n35657_, new_n35658_,
    new_n35659_, new_n35660_, new_n35661_, new_n35662_, new_n35663_,
    new_n35664_, new_n35665_, new_n35666_, new_n35667_, new_n35668_,
    new_n35669_, new_n35670_, new_n35671_, new_n35672_, new_n35673_,
    new_n35674_, new_n35675_, new_n35676_, new_n35677_, new_n35678_,
    new_n35679_, new_n35680_, new_n35681_, new_n35682_, new_n35683_,
    new_n35684_, new_n35685_, new_n35686_, new_n35687_, new_n35688_,
    new_n35689_, new_n35690_, new_n35691_, new_n35692_, new_n35693_,
    new_n35694_, new_n35695_, new_n35696_, new_n35697_, new_n35698_,
    new_n35699_, new_n35700_, new_n35701_, new_n35702_, new_n35703_,
    new_n35704_, new_n35705_, new_n35706_, new_n35707_, new_n35708_,
    new_n35709_, new_n35710_, new_n35711_, new_n35712_, new_n35713_,
    new_n35714_, new_n35715_, new_n35716_, new_n35717_, new_n35718_,
    new_n35719_, new_n35720_, new_n35721_, new_n35722_, new_n35723_,
    new_n35724_, new_n35725_, new_n35726_, new_n35727_, new_n35728_,
    new_n35729_, new_n35730_, new_n35731_, new_n35732_, new_n35733_,
    new_n35734_, new_n35735_, new_n35736_, new_n35737_, new_n35738_,
    new_n35739_, new_n35740_, new_n35741_, new_n35742_, new_n35743_,
    new_n35744_, new_n35745_, new_n35746_, new_n35747_, new_n35748_,
    new_n35749_, new_n35750_, new_n35751_, new_n35752_, new_n35753_,
    new_n35754_, new_n35755_, new_n35756_, new_n35757_, new_n35758_,
    new_n35759_, new_n35760_, new_n35761_, new_n35762_, new_n35763_,
    new_n35764_, new_n35765_, new_n35766_, new_n35767_, new_n35768_,
    new_n35769_, new_n35770_, new_n35771_, new_n35772_, new_n35773_,
    new_n35774_, new_n35775_, new_n35776_, new_n35777_, new_n35778_,
    new_n35779_, new_n35780_, new_n35781_, new_n35782_, new_n35783_,
    new_n35784_, new_n35785_, new_n35786_, new_n35787_, new_n35788_,
    new_n35789_, new_n35790_, new_n35791_, new_n35792_, new_n35793_,
    new_n35794_, new_n35795_, new_n35796_, new_n35797_, new_n35798_,
    new_n35799_, new_n35800_, new_n35801_, new_n35802_, new_n35803_,
    new_n35804_, new_n35805_, new_n35806_, new_n35807_, new_n35808_,
    new_n35809_, new_n35810_, new_n35811_, new_n35812_, new_n35813_,
    new_n35814_, new_n35815_, new_n35816_, new_n35817_, new_n35818_,
    new_n35819_, new_n35820_, new_n35821_, new_n35822_, new_n35823_,
    new_n35824_, new_n35825_, new_n35826_, new_n35827_, new_n35828_,
    new_n35829_, new_n35830_, new_n35831_, new_n35832_, new_n35833_,
    new_n35834_, new_n35835_, new_n35836_, new_n35837_, new_n35838_,
    new_n35839_, new_n35840_, new_n35841_, new_n35842_, new_n35843_,
    new_n35844_, new_n35845_, new_n35846_, new_n35847_, new_n35848_,
    new_n35849_, new_n35850_, new_n35851_, new_n35852_, new_n35853_,
    new_n35854_, new_n35855_, new_n35856_, new_n35857_, new_n35858_,
    new_n35859_, new_n35860_, new_n35861_, new_n35862_, new_n35863_,
    new_n35864_, new_n35865_, new_n35866_, new_n35867_, new_n35868_,
    new_n35869_, new_n35870_, new_n35871_, new_n35872_, new_n35873_,
    new_n35874_, new_n35875_, new_n35876_, new_n35877_, new_n35878_,
    new_n35879_, new_n35880_, new_n35881_, new_n35882_, new_n35883_,
    new_n35884_, new_n35885_, new_n35886_, new_n35887_, new_n35888_,
    new_n35889_, new_n35890_, new_n35891_, new_n35892_, new_n35893_,
    new_n35894_, new_n35895_, new_n35896_, new_n35897_, new_n35898_,
    new_n35899_, new_n35900_, new_n35901_, new_n35902_, new_n35903_,
    new_n35904_, new_n35905_, new_n35906_, new_n35907_, new_n35908_,
    new_n35909_, new_n35910_, new_n35911_, new_n35912_, new_n35913_,
    new_n35914_, new_n35915_, new_n35916_, new_n35917_, new_n35918_,
    new_n35919_, new_n35920_, new_n35921_, new_n35922_, new_n35923_,
    new_n35924_, new_n35925_, new_n35926_, new_n35927_, new_n35928_,
    new_n35929_, new_n35930_, new_n35931_, new_n35932_, new_n35933_,
    new_n35934_, new_n35935_, new_n35936_, new_n35937_, new_n35938_,
    new_n35939_, new_n35940_, new_n35941_, new_n35942_, new_n35943_,
    new_n35944_, new_n35945_, new_n35946_, new_n35947_, new_n35948_,
    new_n35949_, new_n35950_, new_n35951_, new_n35952_, new_n35953_,
    new_n35954_, new_n35955_, new_n35956_, new_n35957_, new_n35958_,
    new_n35959_, new_n35960_, new_n35961_, new_n35962_, new_n35963_,
    new_n35964_, new_n35965_, new_n35966_, new_n35967_, new_n35968_,
    new_n35969_, new_n35970_, new_n35971_, new_n35972_, new_n35973_,
    new_n35974_, new_n35975_, new_n35976_, new_n35977_, new_n35978_,
    new_n35979_, new_n35980_, new_n35981_, new_n35982_, new_n35983_,
    new_n35984_, new_n35985_, new_n35986_, new_n35987_, new_n35988_,
    new_n35989_, new_n35990_, new_n35991_, new_n35992_, new_n35993_,
    new_n35994_, new_n35995_, new_n35996_, new_n35997_, new_n35998_,
    new_n35999_, new_n36000_, new_n36001_, new_n36002_, new_n36003_,
    new_n36004_, new_n36005_, new_n36006_, new_n36007_, new_n36008_,
    new_n36009_, new_n36010_, new_n36011_, new_n36012_, new_n36013_,
    new_n36014_, new_n36015_, new_n36016_, new_n36017_, new_n36018_,
    new_n36019_, new_n36020_, new_n36021_, new_n36022_, new_n36023_,
    new_n36024_, new_n36025_, new_n36026_, new_n36027_, new_n36028_,
    new_n36029_, new_n36030_, new_n36031_, new_n36032_, new_n36033_,
    new_n36034_, new_n36035_, new_n36036_, new_n36037_, new_n36038_,
    new_n36039_, new_n36040_, new_n36041_, new_n36042_, new_n36043_,
    new_n36044_, new_n36045_, new_n36046_, new_n36047_, new_n36048_,
    new_n36049_, new_n36050_, new_n36051_, new_n36052_, new_n36053_,
    new_n36054_, new_n36055_, new_n36056_, new_n36057_, new_n36058_,
    new_n36059_, new_n36060_, new_n36061_, new_n36062_, new_n36063_,
    new_n36064_, new_n36065_, new_n36066_, new_n36067_, new_n36068_,
    new_n36069_, new_n36070_, new_n36071_, new_n36072_, new_n36073_,
    new_n36074_, new_n36075_, new_n36076_, new_n36077_, new_n36078_,
    new_n36079_, new_n36080_, new_n36081_, new_n36082_, new_n36083_,
    new_n36084_, new_n36085_, new_n36086_, new_n36087_, new_n36088_,
    new_n36089_, new_n36090_, new_n36091_, new_n36092_, new_n36093_,
    new_n36094_, new_n36095_, new_n36096_, new_n36097_, new_n36098_,
    new_n36099_, new_n36100_, new_n36101_, new_n36102_, new_n36103_,
    new_n36104_, new_n36105_, new_n36106_, new_n36107_, new_n36108_,
    new_n36109_, new_n36110_, new_n36111_, new_n36112_, new_n36113_,
    new_n36114_, new_n36115_, new_n36116_, new_n36117_, new_n36118_,
    new_n36119_, new_n36120_, new_n36121_, new_n36122_, new_n36123_,
    new_n36124_, new_n36125_, new_n36126_, new_n36127_, new_n36128_,
    new_n36129_, new_n36130_, new_n36131_, new_n36132_, new_n36133_,
    new_n36134_, new_n36135_, new_n36136_, new_n36137_, new_n36138_,
    new_n36139_, new_n36140_, new_n36141_, new_n36142_, new_n36143_,
    new_n36144_, new_n36145_, new_n36146_, new_n36147_, new_n36148_,
    new_n36149_, new_n36150_, new_n36151_, new_n36152_, new_n36153_,
    new_n36154_, new_n36155_, new_n36156_, new_n36157_, new_n36158_,
    new_n36159_, new_n36160_, new_n36161_, new_n36162_, new_n36163_,
    new_n36164_, new_n36165_, new_n36166_, new_n36167_, new_n36168_,
    new_n36169_, new_n36170_, new_n36171_, new_n36172_, new_n36173_,
    new_n36174_, new_n36175_, new_n36176_, new_n36177_, new_n36178_,
    new_n36179_, new_n36180_, new_n36181_, new_n36182_, new_n36183_,
    new_n36184_, new_n36185_, new_n36186_, new_n36187_, new_n36188_,
    new_n36189_, new_n36190_, new_n36191_, new_n36192_, new_n36193_,
    new_n36194_, new_n36195_, new_n36196_, new_n36197_, new_n36198_,
    new_n36199_, new_n36200_, new_n36201_, new_n36202_, new_n36203_,
    new_n36204_, new_n36205_, new_n36206_, new_n36207_, new_n36208_,
    new_n36209_, new_n36210_, new_n36211_, new_n36212_, new_n36213_,
    new_n36214_, new_n36215_, new_n36216_, new_n36217_, new_n36218_,
    new_n36219_, new_n36220_, new_n36221_, new_n36222_, new_n36223_,
    new_n36224_, new_n36225_, new_n36226_, new_n36227_, new_n36228_,
    new_n36229_, new_n36230_, new_n36231_, new_n36232_, new_n36233_,
    new_n36234_, new_n36235_, new_n36236_, new_n36237_, new_n36238_,
    new_n36239_, new_n36240_, new_n36241_, new_n36242_, new_n36243_,
    new_n36244_, new_n36245_, new_n36246_, new_n36247_, new_n36248_,
    new_n36249_, new_n36250_, new_n36251_, new_n36252_, new_n36253_,
    new_n36254_, new_n36255_, new_n36256_, new_n36257_, new_n36258_,
    new_n36259_, new_n36260_, new_n36261_, new_n36262_, new_n36263_,
    new_n36264_, new_n36265_, new_n36266_, new_n36267_, new_n36268_,
    new_n36269_, new_n36270_, new_n36271_, new_n36272_, new_n36273_,
    new_n36274_, new_n36275_, new_n36276_, new_n36277_, new_n36278_,
    new_n36279_, new_n36280_, new_n36281_, new_n36282_, new_n36283_,
    new_n36284_, new_n36285_, new_n36286_, new_n36287_, new_n36288_,
    new_n36289_, new_n36290_, new_n36291_, new_n36292_, new_n36293_,
    new_n36294_, new_n36295_, new_n36296_, new_n36297_, new_n36298_,
    new_n36299_, new_n36300_, new_n36301_, new_n36302_, new_n36303_,
    new_n36304_, new_n36305_, new_n36306_, new_n36307_, new_n36308_,
    new_n36309_, new_n36310_, new_n36311_, new_n36312_, new_n36313_,
    new_n36314_, new_n36315_, new_n36316_, new_n36317_, new_n36318_,
    new_n36319_, new_n36320_, new_n36321_, new_n36322_, new_n36323_,
    new_n36324_, new_n36325_, new_n36326_, new_n36327_, new_n36328_,
    new_n36329_, new_n36330_, new_n36331_, new_n36332_, new_n36333_,
    new_n36334_, new_n36335_, new_n36336_, new_n36337_, new_n36338_,
    new_n36339_, new_n36340_, new_n36341_, new_n36342_, new_n36343_,
    new_n36344_, new_n36345_, new_n36346_, new_n36347_, new_n36348_,
    new_n36349_, new_n36350_, new_n36351_, new_n36352_, new_n36353_,
    new_n36354_, new_n36355_, new_n36356_, new_n36357_, new_n36358_,
    new_n36359_, new_n36360_, new_n36361_, new_n36362_, new_n36363_,
    new_n36364_, new_n36365_, new_n36366_, new_n36367_, new_n36368_,
    new_n36369_, new_n36370_, new_n36371_, new_n36372_, new_n36373_,
    new_n36374_, new_n36375_, new_n36376_, new_n36377_, new_n36378_,
    new_n36379_, new_n36380_, new_n36381_, new_n36382_, new_n36383_,
    new_n36384_, new_n36385_, new_n36386_, new_n36387_, new_n36388_,
    new_n36389_, new_n36390_, new_n36391_, new_n36392_, new_n36393_,
    new_n36394_, new_n36395_, new_n36396_, new_n36397_, new_n36398_,
    new_n36399_, new_n36400_, new_n36401_, new_n36402_, new_n36403_,
    new_n36404_, new_n36405_, new_n36406_, new_n36407_, new_n36408_,
    new_n36409_, new_n36410_, new_n36411_, new_n36412_, new_n36413_,
    new_n36414_, new_n36415_, new_n36416_, new_n36417_, new_n36418_,
    new_n36419_, new_n36420_, new_n36421_, new_n36422_, new_n36423_,
    new_n36424_, new_n36425_, new_n36426_, new_n36427_, new_n36428_,
    new_n36429_, new_n36430_, new_n36431_, new_n36432_, new_n36433_,
    new_n36434_, new_n36435_, new_n36436_, new_n36437_, new_n36438_,
    new_n36439_, new_n36440_, new_n36441_, new_n36442_, new_n36443_,
    new_n36444_, new_n36445_, new_n36446_, new_n36447_, new_n36448_,
    new_n36449_, new_n36450_, new_n36451_, new_n36452_, new_n36453_,
    new_n36454_, new_n36455_, new_n36456_, new_n36457_, new_n36458_,
    new_n36459_, new_n36460_, new_n36461_, new_n36462_, new_n36463_,
    new_n36464_, new_n36465_, new_n36466_, new_n36467_, new_n36468_,
    new_n36469_, new_n36470_, new_n36471_, new_n36472_, new_n36473_,
    new_n36474_, new_n36475_, new_n36476_, new_n36477_, new_n36478_,
    new_n36479_, new_n36480_, new_n36481_, new_n36482_, new_n36483_,
    new_n36484_, new_n36485_, new_n36486_, new_n36487_, new_n36488_,
    new_n36489_, new_n36490_, new_n36491_, new_n36492_, new_n36493_,
    new_n36494_, new_n36495_, new_n36496_, new_n36497_, new_n36498_,
    new_n36499_, new_n36500_, new_n36501_, new_n36502_, new_n36503_,
    new_n36504_, new_n36505_, new_n36506_, new_n36507_, new_n36508_,
    new_n36509_, new_n36510_, new_n36511_, new_n36512_, new_n36513_,
    new_n36514_, new_n36515_, new_n36516_, new_n36517_, new_n36518_,
    new_n36519_, new_n36520_, new_n36521_, new_n36522_, new_n36523_,
    new_n36524_, new_n36525_, new_n36526_, new_n36527_, new_n36528_,
    new_n36529_, new_n36530_, new_n36531_, new_n36532_, new_n36533_,
    new_n36534_, new_n36535_, new_n36536_, new_n36537_, new_n36538_,
    new_n36539_, new_n36540_, new_n36541_, new_n36542_, new_n36543_,
    new_n36544_, new_n36545_, new_n36546_, new_n36547_, new_n36548_,
    new_n36549_, new_n36550_, new_n36551_, new_n36552_, new_n36553_,
    new_n36554_, new_n36555_, new_n36556_, new_n36557_, new_n36558_,
    new_n36559_, new_n36560_, new_n36561_, new_n36562_, new_n36563_,
    new_n36564_, new_n36565_, new_n36566_, new_n36567_, new_n36568_,
    new_n36569_, new_n36570_, new_n36571_, new_n36572_, new_n36573_,
    new_n36574_, new_n36575_, new_n36576_, new_n36577_, new_n36578_,
    new_n36579_, new_n36580_, new_n36581_, new_n36582_, new_n36583_,
    new_n36584_, new_n36585_, new_n36586_, new_n36587_, new_n36588_,
    new_n36589_, new_n36590_, new_n36591_, new_n36592_, new_n36593_,
    new_n36594_, new_n36595_, new_n36596_, new_n36597_, new_n36598_,
    new_n36599_, new_n36600_, new_n36601_, new_n36602_, new_n36603_,
    new_n36604_, new_n36605_, new_n36606_, new_n36607_, new_n36608_,
    new_n36609_, new_n36610_, new_n36611_, new_n36612_, new_n36613_,
    new_n36614_, new_n36615_, new_n36616_, new_n36617_, new_n36618_,
    new_n36619_, new_n36620_, new_n36621_, new_n36622_, new_n36623_,
    new_n36624_, new_n36625_, new_n36626_, new_n36627_, new_n36628_,
    new_n36629_, new_n36630_, new_n36631_, new_n36632_, new_n36633_,
    new_n36634_, new_n36635_, new_n36636_, new_n36637_, new_n36638_,
    new_n36639_, new_n36640_, new_n36641_, new_n36642_, new_n36643_,
    new_n36644_, new_n36645_, new_n36646_, new_n36647_, new_n36648_,
    new_n36649_, new_n36650_, new_n36651_, new_n36652_, new_n36653_,
    new_n36654_, new_n36655_, new_n36656_, new_n36657_, new_n36658_,
    new_n36659_, new_n36660_, new_n36661_, new_n36662_, new_n36663_,
    new_n36664_, new_n36665_, new_n36666_, new_n36667_, new_n36668_,
    new_n36669_, new_n36670_, new_n36671_, new_n36672_, new_n36673_,
    new_n36674_, new_n36675_, new_n36676_, new_n36677_, new_n36678_,
    new_n36679_, new_n36680_, new_n36681_, new_n36682_, new_n36683_,
    new_n36684_, new_n36685_, new_n36686_, new_n36687_, new_n36688_,
    new_n36689_, new_n36690_, new_n36691_, new_n36692_, new_n36693_,
    new_n36694_, new_n36695_, new_n36696_, new_n36697_, new_n36698_,
    new_n36699_, new_n36700_, new_n36701_, new_n36702_, new_n36703_,
    new_n36704_, new_n36705_, new_n36706_, new_n36707_, new_n36708_,
    new_n36709_, new_n36710_, new_n36711_, new_n36712_, new_n36713_,
    new_n36714_, new_n36715_, new_n36716_, new_n36717_, new_n36718_,
    new_n36719_, new_n36720_, new_n36721_, new_n36722_, new_n36723_,
    new_n36724_, new_n36725_, new_n36726_, new_n36727_, new_n36728_,
    new_n36729_, new_n36730_, new_n36731_, new_n36732_, new_n36733_,
    new_n36734_, new_n36735_, new_n36736_, new_n36737_, new_n36738_,
    new_n36739_, new_n36740_, new_n36741_, new_n36742_, new_n36743_,
    new_n36744_, new_n36745_, new_n36746_, new_n36747_, new_n36748_,
    new_n36749_, new_n36750_, new_n36751_, new_n36752_, new_n36753_,
    new_n36754_, new_n36755_, new_n36756_, new_n36757_, new_n36758_,
    new_n36759_, new_n36760_, new_n36761_, new_n36762_, new_n36763_,
    new_n36764_, new_n36765_, new_n36766_, new_n36767_, new_n36768_,
    new_n36769_, new_n36770_, new_n36771_, new_n36772_, new_n36773_,
    new_n36774_, new_n36775_, new_n36776_, new_n36777_, new_n36778_,
    new_n36779_, new_n36780_, new_n36781_, new_n36782_, new_n36783_,
    new_n36784_, new_n36785_, new_n36786_, new_n36787_, new_n36788_,
    new_n36789_, new_n36790_, new_n36791_, new_n36792_, new_n36793_,
    new_n36794_, new_n36795_, new_n36796_, new_n36797_, new_n36798_,
    new_n36799_, new_n36800_, new_n36801_, new_n36802_, new_n36803_,
    new_n36804_, new_n36805_, new_n36806_, new_n36807_, new_n36808_,
    new_n36809_, new_n36810_, new_n36811_, new_n36812_, new_n36813_,
    new_n36814_, new_n36815_, new_n36816_, new_n36817_, new_n36818_,
    new_n36819_, new_n36820_, new_n36821_, new_n36822_, new_n36823_,
    new_n36824_, new_n36825_, new_n36826_, new_n36827_, new_n36828_,
    new_n36829_, new_n36830_, new_n36831_, new_n36832_, new_n36833_,
    new_n36834_, new_n36835_, new_n36836_, new_n36837_, new_n36838_,
    new_n36839_, new_n36840_, new_n36841_, new_n36842_, new_n36843_,
    new_n36844_, new_n36845_, new_n36846_, new_n36847_, new_n36848_,
    new_n36849_, new_n36850_, new_n36851_, new_n36852_, new_n36853_,
    new_n36854_, new_n36855_, new_n36856_, new_n36857_, new_n36858_,
    new_n36859_, new_n36860_, new_n36861_, new_n36862_, new_n36863_,
    new_n36864_, new_n36865_, new_n36866_, new_n36867_, new_n36868_,
    new_n36869_, new_n36870_, new_n36871_, new_n36872_, new_n36873_,
    new_n36874_, new_n36875_, new_n36876_, new_n36877_, new_n36878_,
    new_n36879_, new_n36880_, new_n36881_, new_n36882_, new_n36883_,
    new_n36884_, new_n36885_, new_n36886_, new_n36887_, new_n36888_,
    new_n36889_, new_n36890_, new_n36891_, new_n36892_, new_n36893_,
    new_n36894_, new_n36895_, new_n36896_, new_n36897_, new_n36898_,
    new_n36899_, new_n36900_, new_n36901_, new_n36902_, new_n36903_,
    new_n36904_, new_n36905_, new_n36906_, new_n36907_, new_n36908_,
    new_n36909_, new_n36910_, new_n36911_, new_n36912_, new_n36913_,
    new_n36914_, new_n36915_, new_n36916_, new_n36917_, new_n36918_,
    new_n36919_, new_n36920_, new_n36921_, new_n36922_, new_n36923_,
    new_n36924_, new_n36925_, new_n36926_, new_n36927_, new_n36928_,
    new_n36929_, new_n36930_, new_n36931_, new_n36932_, new_n36933_,
    new_n36934_, new_n36935_, new_n36936_, new_n36937_, new_n36938_,
    new_n36939_, new_n36940_, new_n36941_, new_n36942_, new_n36943_,
    new_n36944_, new_n36945_, new_n36946_, new_n36947_, new_n36948_,
    new_n36949_, new_n36950_, new_n36951_, new_n36952_, new_n36953_,
    new_n36954_, new_n36955_, new_n36956_, new_n36957_, new_n36958_,
    new_n36959_, new_n36960_, new_n36961_, new_n36962_, new_n36963_,
    new_n36964_, new_n36965_, new_n36966_, new_n36967_, new_n36968_,
    new_n36969_, new_n36970_, new_n36971_, new_n36972_, new_n36973_,
    new_n36974_, new_n36975_, new_n36976_, new_n36977_, new_n36978_,
    new_n36979_, new_n36980_, new_n36981_, new_n36982_, new_n36983_,
    new_n36984_, new_n36985_, new_n36986_, new_n36987_, new_n36988_,
    new_n36989_, new_n36990_, new_n36991_, new_n36992_, new_n36993_,
    new_n36994_, new_n36995_, new_n36996_, new_n36997_, new_n36998_,
    new_n36999_, new_n37000_, new_n37001_, new_n37002_, new_n37003_,
    new_n37004_, new_n37005_, new_n37006_, new_n37007_, new_n37008_,
    new_n37009_, new_n37010_, new_n37011_, new_n37012_, new_n37013_,
    new_n37014_, new_n37015_, new_n37016_, new_n37017_, new_n37018_,
    new_n37019_, new_n37020_, new_n37021_, new_n37022_, new_n37023_,
    new_n37024_, new_n37025_, new_n37026_, new_n37027_, new_n37028_,
    new_n37029_, new_n37030_, new_n37031_, new_n37032_, new_n37033_,
    new_n37034_, new_n37035_, new_n37036_, new_n37037_, new_n37038_,
    new_n37039_, new_n37040_, new_n37041_, new_n37042_, new_n37043_,
    new_n37044_, new_n37045_, new_n37046_, new_n37047_, new_n37048_,
    new_n37049_, new_n37050_, new_n37051_, new_n37052_, new_n37053_,
    new_n37054_, new_n37055_, new_n37056_, new_n37057_, new_n37058_,
    new_n37059_, new_n37060_, new_n37061_, new_n37062_, new_n37063_,
    new_n37064_, new_n37065_, new_n37066_, new_n37067_, new_n37068_,
    new_n37069_, new_n37070_, new_n37071_, new_n37072_, new_n37073_,
    new_n37074_, new_n37075_, new_n37076_, new_n37077_, new_n37078_,
    new_n37079_, new_n37080_, new_n37081_, new_n37082_, new_n37083_,
    new_n37084_, new_n37085_, new_n37086_, new_n37087_, new_n37088_,
    new_n37089_, new_n37090_, new_n37091_, new_n37092_, new_n37093_,
    new_n37094_, new_n37095_, new_n37096_, new_n37097_, new_n37098_,
    new_n37099_, new_n37100_, new_n37101_, new_n37102_, new_n37103_,
    new_n37104_, new_n37105_, new_n37106_, new_n37107_, new_n37108_,
    new_n37109_, new_n37110_, new_n37111_, new_n37112_, new_n37113_,
    new_n37114_, new_n37115_, new_n37116_, new_n37117_, new_n37118_,
    new_n37119_, new_n37120_, new_n37121_, new_n37122_, new_n37123_,
    new_n37124_, new_n37125_, new_n37126_, new_n37127_, new_n37128_,
    new_n37129_, new_n37130_, new_n37131_, new_n37132_, new_n37133_,
    new_n37134_, new_n37135_, new_n37136_, new_n37137_, new_n37138_,
    new_n37139_, new_n37140_, new_n37141_, new_n37142_, new_n37143_,
    new_n37144_, new_n37145_, new_n37146_, new_n37147_, new_n37148_,
    new_n37149_, new_n37150_, new_n37151_, new_n37152_, new_n37153_,
    new_n37154_, new_n37155_, new_n37156_, new_n37157_, new_n37158_,
    new_n37159_, new_n37160_, new_n37161_, new_n37162_, new_n37163_,
    new_n37164_, new_n37165_, new_n37166_, new_n37167_, new_n37168_,
    new_n37169_, new_n37170_, new_n37171_, new_n37172_, new_n37173_,
    new_n37174_, new_n37175_, new_n37176_, new_n37177_, new_n37178_,
    new_n37179_, new_n37180_, new_n37181_, new_n37182_, new_n37183_,
    new_n37184_, new_n37185_, new_n37186_, new_n37187_, new_n37188_,
    new_n37189_, new_n37190_, new_n37191_, new_n37192_, new_n37193_,
    new_n37194_, new_n37195_, new_n37196_, new_n37197_, new_n37198_,
    new_n37199_, new_n37200_, new_n37201_, new_n37202_, new_n37203_,
    new_n37204_, new_n37205_, new_n37206_, new_n37207_, new_n37208_,
    new_n37209_, new_n37210_, new_n37211_, new_n37212_, new_n37213_,
    new_n37214_, new_n37215_, new_n37216_, new_n37217_, new_n37218_,
    new_n37219_, new_n37220_, new_n37221_, new_n37222_, new_n37223_,
    new_n37224_, new_n37225_, new_n37226_, new_n37227_, new_n37228_,
    new_n37229_, new_n37230_, new_n37231_, new_n37232_, new_n37233_,
    new_n37234_, new_n37235_, new_n37236_, new_n37237_, new_n37238_,
    new_n37239_, new_n37240_, new_n37241_, new_n37242_, new_n37243_,
    new_n37244_, new_n37245_, new_n37246_, new_n37247_, new_n37248_,
    new_n37249_, new_n37250_, new_n37251_, new_n37252_, new_n37253_,
    new_n37254_, new_n37255_, new_n37256_, new_n37257_, new_n37258_,
    new_n37259_, new_n37260_, new_n37261_, new_n37262_, new_n37263_,
    new_n37264_, new_n37265_, new_n37266_, new_n37267_, new_n37268_,
    new_n37269_, new_n37270_, new_n37271_, new_n37272_, new_n37273_,
    new_n37274_, new_n37275_, new_n37276_, new_n37277_, new_n37278_,
    new_n37279_, new_n37280_, new_n37281_, new_n37282_, new_n37283_,
    new_n37284_, new_n37285_, new_n37286_, new_n37287_, new_n37288_,
    new_n37289_, new_n37290_, new_n37291_, new_n37292_, new_n37293_,
    new_n37294_, new_n37295_, new_n37296_, new_n37297_, new_n37298_,
    new_n37299_, new_n37300_, new_n37301_, new_n37302_, new_n37303_,
    new_n37304_, new_n37305_, new_n37306_, new_n37307_, new_n37308_,
    new_n37309_, new_n37310_, new_n37311_, new_n37312_, new_n37313_,
    new_n37314_, new_n37315_, new_n37316_, new_n37317_, new_n37318_,
    new_n37319_, new_n37320_, new_n37321_, new_n37322_, new_n37323_,
    new_n37324_, new_n37325_, new_n37326_, new_n37327_, new_n37328_,
    new_n37329_, new_n37330_, new_n37331_, new_n37332_, new_n37333_,
    new_n37334_, new_n37335_, new_n37336_, new_n37337_, new_n37338_,
    new_n37339_, new_n37340_, new_n37341_, new_n37342_, new_n37343_,
    new_n37344_, new_n37345_, new_n37346_, new_n37347_, new_n37348_,
    new_n37349_, new_n37350_, new_n37351_, new_n37352_, new_n37353_,
    new_n37354_, new_n37355_, new_n37356_, new_n37357_, new_n37358_,
    new_n37359_, new_n37360_, new_n37361_, new_n37362_, new_n37363_,
    new_n37364_, new_n37365_, new_n37366_, new_n37367_, new_n37368_,
    new_n37369_, new_n37370_, new_n37371_, new_n37372_, new_n37373_,
    new_n37374_, new_n37375_, new_n37376_, new_n37377_, new_n37378_,
    new_n37379_, new_n37380_, new_n37381_, new_n37382_, new_n37383_,
    new_n37384_, new_n37385_, new_n37386_, new_n37387_, new_n37388_,
    new_n37389_, new_n37390_, new_n37391_, new_n37392_, new_n37393_,
    new_n37394_, new_n37395_, new_n37396_, new_n37397_, new_n37398_,
    new_n37399_, new_n37400_, new_n37401_, new_n37402_, new_n37403_,
    new_n37404_, new_n37405_, new_n37406_, new_n37407_, new_n37408_,
    new_n37409_, new_n37410_, new_n37411_, new_n37412_, new_n37413_,
    new_n37414_, new_n37415_, new_n37416_, new_n37417_, new_n37418_,
    new_n37419_, new_n37420_, new_n37421_, new_n37422_, new_n37423_,
    new_n37424_, new_n37425_, new_n37426_, new_n37427_, new_n37428_,
    new_n37429_, new_n37430_, new_n37431_, new_n37432_, new_n37433_,
    new_n37434_, new_n37435_, new_n37436_, new_n37437_, new_n37438_,
    new_n37439_, new_n37440_, new_n37441_, new_n37442_, new_n37443_,
    new_n37444_, new_n37445_, new_n37446_, new_n37447_, new_n37448_,
    new_n37449_, new_n37450_, new_n37451_, new_n37452_, new_n37453_,
    new_n37454_, new_n37455_, new_n37456_, new_n37457_, new_n37458_,
    new_n37459_, new_n37460_, new_n37461_, new_n37462_, new_n37463_,
    new_n37464_, new_n37465_, new_n37466_, new_n37467_, new_n37468_,
    new_n37469_, new_n37470_, new_n37471_, new_n37472_, new_n37473_,
    new_n37474_, new_n37475_, new_n37476_, new_n37477_, new_n37478_,
    new_n37479_, new_n37480_, new_n37481_, new_n37482_, new_n37483_,
    new_n37484_, new_n37485_, new_n37486_, new_n37487_, new_n37488_,
    new_n37489_, new_n37490_, new_n37491_, new_n37492_, new_n37493_,
    new_n37494_, new_n37495_, new_n37496_, new_n37497_, new_n37498_,
    new_n37499_, new_n37500_, new_n37501_, new_n37502_, new_n37503_,
    new_n37504_, new_n37505_, new_n37506_, new_n37507_, new_n37508_,
    new_n37509_, new_n37510_, new_n37511_, new_n37512_, new_n37513_,
    new_n37514_, new_n37515_, new_n37516_, new_n37517_, new_n37518_,
    new_n37519_, new_n37520_, new_n37521_, new_n37522_, new_n37523_,
    new_n37524_, new_n37525_, new_n37526_, new_n37527_, new_n37528_,
    new_n37529_, new_n37530_, new_n37531_, new_n37532_, new_n37533_,
    new_n37534_, new_n37535_, new_n37536_, new_n37537_, new_n37538_,
    new_n37539_, new_n37540_, new_n37541_, new_n37542_, new_n37543_,
    new_n37544_, new_n37545_, new_n37546_, new_n37547_, new_n37548_,
    new_n37549_, new_n37550_, new_n37551_, new_n37552_, new_n37553_,
    new_n37554_, new_n37555_, new_n37556_, new_n37557_, new_n37558_,
    new_n37559_, new_n37560_, new_n37561_, new_n37562_, new_n37563_,
    new_n37564_, new_n37565_, new_n37566_, new_n37567_, new_n37568_,
    new_n37569_, new_n37570_, new_n37571_, new_n37572_, new_n37573_,
    new_n37574_, new_n37575_, new_n37576_, new_n37577_, new_n37578_,
    new_n37579_, new_n37580_, new_n37581_, new_n37582_, new_n37583_,
    new_n37584_, new_n37585_, new_n37586_, new_n37587_, new_n37588_,
    new_n37589_, new_n37590_, new_n37591_, new_n37592_, new_n37593_,
    new_n37594_, new_n37595_, new_n37596_, new_n37597_, new_n37598_,
    new_n37599_, new_n37600_, new_n37601_, new_n37602_, new_n37603_,
    new_n37604_, new_n37605_, new_n37606_, new_n37607_, new_n37608_,
    new_n37609_, new_n37610_, new_n37611_, new_n37612_, new_n37613_,
    new_n37614_, new_n37615_, new_n37616_, new_n37617_, new_n37618_,
    new_n37619_, new_n37620_, new_n37621_, new_n37622_, new_n37623_,
    new_n37624_, new_n37625_, new_n37626_, new_n37627_, new_n37628_,
    new_n37629_, new_n37630_, new_n37631_, new_n37632_, new_n37633_,
    new_n37634_, new_n37635_, new_n37636_, new_n37637_, new_n37638_,
    new_n37639_, new_n37640_, new_n37641_, new_n37642_, new_n37643_,
    new_n37644_, new_n37645_, new_n37646_, new_n37647_, new_n37648_,
    new_n37649_, new_n37650_, new_n37651_, new_n37652_, new_n37653_,
    new_n37654_, new_n37655_, new_n37656_, new_n37657_, new_n37658_,
    new_n37659_, new_n37660_, new_n37661_, new_n37662_, new_n37663_,
    new_n37664_, new_n37665_, new_n37666_, new_n37667_, new_n37668_,
    new_n37669_, new_n37670_, new_n37671_, new_n37672_, new_n37673_,
    new_n37674_, new_n37675_, new_n37676_, new_n37677_, new_n37678_,
    new_n37679_, new_n37680_, new_n37681_, new_n37682_, new_n37683_,
    new_n37684_, new_n37685_, new_n37686_, new_n37687_, new_n37688_,
    new_n37689_, new_n37690_, new_n37691_, new_n37692_, new_n37693_,
    new_n37694_, new_n37695_, new_n37696_, new_n37697_, new_n37698_,
    new_n37699_, new_n37700_, new_n37701_, new_n37702_, new_n37703_,
    new_n37704_, new_n37705_, new_n37706_, new_n37707_, new_n37708_,
    new_n37709_, new_n37710_, new_n37711_, new_n37712_, new_n37713_,
    new_n37714_, new_n37715_, new_n37716_, new_n37717_, new_n37718_,
    new_n37719_, new_n37720_, new_n37721_, new_n37722_, new_n37723_,
    new_n37724_, new_n37725_, new_n37726_, new_n37727_, new_n37728_,
    new_n37729_, new_n37730_, new_n37731_, new_n37732_, new_n37733_,
    new_n37734_, new_n37735_, new_n37736_, new_n37737_, new_n37738_,
    new_n37739_, new_n37740_, new_n37741_, new_n37742_, new_n37743_,
    new_n37744_, new_n37745_, new_n37746_, new_n37747_, new_n37748_,
    new_n37749_, new_n37750_, new_n37751_, new_n37752_, new_n37753_,
    new_n37754_, new_n37755_, new_n37756_, new_n37757_, new_n37758_,
    new_n37759_, new_n37760_, new_n37761_, new_n37762_, new_n37763_,
    new_n37764_, new_n37765_, new_n37766_, new_n37767_, new_n37768_,
    new_n37769_, new_n37770_, new_n37771_, new_n37772_, new_n37773_,
    new_n37774_, new_n37775_, new_n37776_, new_n37777_, new_n37778_,
    new_n37779_, new_n37780_, new_n37781_, new_n37782_, new_n37783_,
    new_n37784_, new_n37785_, new_n37786_, new_n37787_, new_n37788_,
    new_n37789_, new_n37790_, new_n37791_, new_n37792_, new_n37793_,
    new_n37794_, new_n37795_, new_n37796_, new_n37797_, new_n37798_,
    new_n37799_, new_n37800_, new_n37801_, new_n37802_, new_n37803_,
    new_n37804_, new_n37805_, new_n37806_, new_n37807_, new_n37808_,
    new_n37809_, new_n37810_, new_n37811_, new_n37812_, new_n37813_,
    new_n37814_, new_n37815_, new_n37816_, new_n37817_, new_n37818_,
    new_n37819_, new_n37820_, new_n37821_, new_n37822_, new_n37823_,
    new_n37824_, new_n37825_, new_n37826_, new_n37827_, new_n37828_,
    new_n37829_, new_n37830_, new_n37831_, new_n37832_, new_n37833_,
    new_n37834_, new_n37835_, new_n37836_, new_n37837_, new_n37838_,
    new_n37839_, new_n37840_, new_n37841_, new_n37842_, new_n37843_,
    new_n37844_, new_n37845_, new_n37846_, new_n37847_, new_n37848_,
    new_n37849_, new_n37850_, new_n37851_, new_n37852_, new_n37853_,
    new_n37854_, new_n37855_, new_n37856_, new_n37857_, new_n37858_,
    new_n37859_, new_n37860_, new_n37861_, new_n37862_, new_n37863_,
    new_n37864_, new_n37865_, new_n37866_, new_n37867_, new_n37868_,
    new_n37869_, new_n37870_, new_n37871_, new_n37872_, new_n37873_,
    new_n37874_, new_n37875_, new_n37876_, new_n37877_, new_n37878_,
    new_n37879_, new_n37880_, new_n37881_, new_n37882_, new_n37883_,
    new_n37884_, new_n37885_, new_n37886_, new_n37887_, new_n37888_,
    new_n37889_, new_n37890_, new_n37891_, new_n37892_, new_n37893_,
    new_n37894_, new_n37895_, new_n37896_, new_n37897_, new_n37898_,
    new_n37899_, new_n37900_, new_n37901_, new_n37902_, new_n37903_,
    new_n37904_, new_n37905_, new_n37906_, new_n37907_, new_n37908_,
    new_n37909_, new_n37910_, new_n37911_, new_n37912_, new_n37913_,
    new_n37914_, new_n37915_, new_n37916_, new_n37917_, new_n37918_,
    new_n37919_, new_n37920_, new_n37921_, new_n37922_, new_n37923_,
    new_n37924_, new_n37925_, new_n37926_, new_n37927_, new_n37928_,
    new_n37929_, new_n37930_, new_n37931_, new_n37932_, new_n37933_,
    new_n37934_, new_n37935_, new_n37936_, new_n37937_, new_n37938_,
    new_n37939_, new_n37940_, new_n37941_, new_n37942_, new_n37943_,
    new_n37944_, new_n37945_, new_n37946_, new_n37947_, new_n37948_,
    new_n37949_, new_n37950_, new_n37951_, new_n37952_, new_n37953_,
    new_n37954_, new_n37955_, new_n37956_, new_n37957_, new_n37958_,
    new_n37959_, new_n37960_, new_n37961_, new_n37962_, new_n37963_,
    new_n37964_, new_n37965_, new_n37966_, new_n37967_, new_n37968_,
    new_n37969_, new_n37970_, new_n37971_, new_n37972_, new_n37973_,
    new_n37974_, new_n37975_, new_n37976_, new_n37977_, new_n37978_,
    new_n37979_, new_n37980_, new_n37981_, new_n37982_, new_n37983_,
    new_n37984_, new_n37985_, new_n37986_, new_n37987_, new_n37988_,
    new_n37989_, new_n37990_, new_n37991_, new_n37992_, new_n37993_,
    new_n37994_, new_n37995_, new_n37996_, new_n37997_, new_n37998_,
    new_n37999_, new_n38000_, new_n38001_, new_n38002_, new_n38003_,
    new_n38004_, new_n38005_, new_n38006_, new_n38007_, new_n38008_,
    new_n38009_, new_n38010_, new_n38011_, new_n38012_, new_n38013_,
    new_n38014_, new_n38015_, new_n38016_, new_n38017_, new_n38018_,
    new_n38019_, new_n38020_, new_n38021_, new_n38022_, new_n38023_,
    new_n38024_, new_n38025_, new_n38026_, new_n38027_, new_n38028_,
    new_n38029_, new_n38030_, new_n38031_, new_n38032_, new_n38033_,
    new_n38034_, new_n38035_, new_n38036_, new_n38037_, new_n38038_,
    new_n38039_, new_n38040_, new_n38041_, new_n38042_, new_n38043_,
    new_n38044_, new_n38045_, new_n38046_, new_n38047_, new_n38048_,
    new_n38049_, new_n38050_, new_n38051_, new_n38052_, new_n38053_,
    new_n38054_, new_n38055_, new_n38056_, new_n38057_, new_n38058_,
    new_n38059_, new_n38060_, new_n38061_, new_n38062_, new_n38063_,
    new_n38064_, new_n38065_, new_n38066_, new_n38067_, new_n38068_,
    new_n38069_, new_n38070_, new_n38071_, new_n38072_, new_n38073_,
    new_n38074_, new_n38075_, new_n38076_, new_n38077_, new_n38078_,
    new_n38079_, new_n38080_, new_n38081_, new_n38082_, new_n38083_,
    new_n38084_, new_n38085_, new_n38086_, new_n38087_, new_n38088_,
    new_n38089_, new_n38090_, new_n38091_, new_n38092_, new_n38093_,
    new_n38094_, new_n38095_, new_n38096_, new_n38097_, new_n38098_,
    new_n38099_, new_n38100_, new_n38101_, new_n38102_, new_n38103_,
    new_n38104_, new_n38105_, new_n38106_, new_n38107_, new_n38108_,
    new_n38109_, new_n38110_, new_n38111_, new_n38112_, new_n38113_,
    new_n38114_, new_n38115_, new_n38116_, new_n38117_, new_n38118_,
    new_n38119_, new_n38120_, new_n38121_, new_n38122_, new_n38123_,
    new_n38124_, new_n38125_, new_n38126_, new_n38127_, new_n38128_,
    new_n38129_, new_n38130_, new_n38131_, new_n38132_, new_n38133_,
    new_n38134_, new_n38135_, new_n38136_, new_n38137_, new_n38138_,
    new_n38139_, new_n38140_, new_n38141_, new_n38142_, new_n38143_,
    new_n38144_, new_n38145_, new_n38146_, new_n38147_, new_n38148_,
    new_n38149_, new_n38150_, new_n38151_, new_n38152_, new_n38153_,
    new_n38154_, new_n38155_, new_n38156_, new_n38157_, new_n38158_,
    new_n38159_, new_n38160_, new_n38161_, new_n38162_, new_n38163_,
    new_n38164_, new_n38165_, new_n38166_, new_n38167_, new_n38168_,
    new_n38169_, new_n38170_, new_n38171_, new_n38172_, new_n38173_,
    new_n38174_, new_n38175_, new_n38176_, new_n38177_, new_n38178_,
    new_n38179_, new_n38180_, new_n38181_, new_n38182_, new_n38183_,
    new_n38184_, new_n38185_, new_n38186_, new_n38187_, new_n38188_,
    new_n38189_, new_n38190_, new_n38191_, new_n38192_, new_n38193_,
    new_n38194_, new_n38195_, new_n38196_, new_n38197_, new_n38198_,
    new_n38199_, new_n38200_, new_n38201_, new_n38202_, new_n38203_,
    new_n38204_, new_n38205_, new_n38206_, new_n38207_, new_n38208_,
    new_n38209_, new_n38210_, new_n38211_, new_n38212_, new_n38213_,
    new_n38214_, new_n38215_, new_n38216_, new_n38217_, new_n38218_,
    new_n38219_, new_n38220_, new_n38221_, new_n38222_, new_n38223_,
    new_n38224_, new_n38225_, new_n38226_, new_n38227_, new_n38228_,
    new_n38229_, new_n38230_, new_n38231_, new_n38232_, new_n38233_,
    new_n38234_, new_n38235_, new_n38236_, new_n38237_, new_n38238_,
    new_n38239_, new_n38240_, new_n38241_, new_n38242_, new_n38243_,
    new_n38244_, new_n38245_, new_n38246_, new_n38247_, new_n38248_,
    new_n38249_, new_n38250_, new_n38251_, new_n38252_, new_n38253_,
    new_n38254_, new_n38255_, new_n38256_, new_n38257_, new_n38258_,
    new_n38259_, new_n38260_, new_n38261_, new_n38262_, new_n38263_,
    new_n38264_, new_n38265_, new_n38266_, new_n38267_, new_n38268_,
    new_n38269_, new_n38270_, new_n38271_, new_n38272_, new_n38273_,
    new_n38274_, new_n38275_, new_n38276_, new_n38277_, new_n38278_,
    new_n38279_, new_n38280_, new_n38281_, new_n38282_, new_n38283_,
    new_n38284_, new_n38285_, new_n38286_, new_n38287_, new_n38288_,
    new_n38289_, new_n38290_, new_n38291_, new_n38292_, new_n38293_,
    new_n38294_, new_n38295_, new_n38296_, new_n38297_, new_n38298_,
    new_n38299_, new_n38300_, new_n38301_, new_n38302_, new_n38303_,
    new_n38304_, new_n38305_, new_n38306_, new_n38307_, new_n38308_,
    new_n38309_, new_n38310_, new_n38311_, new_n38312_, new_n38313_,
    new_n38314_, new_n38315_, new_n38316_, new_n38317_, new_n38318_,
    new_n38319_, new_n38320_, new_n38321_, new_n38322_, new_n38323_,
    new_n38324_, new_n38325_, new_n38326_, new_n38327_, new_n38328_,
    new_n38329_, new_n38330_, new_n38331_, new_n38332_, new_n38333_,
    new_n38334_, new_n38335_, new_n38336_, new_n38337_, new_n38338_,
    new_n38339_, new_n38340_, new_n38341_, new_n38342_, new_n38343_,
    new_n38344_, new_n38345_, new_n38346_, new_n38347_, new_n38348_,
    new_n38349_, new_n38350_, new_n38351_, new_n38352_, new_n38353_,
    new_n38354_, new_n38355_, new_n38356_, new_n38357_, new_n38358_,
    new_n38359_, new_n38360_, new_n38361_, new_n38362_, new_n38363_,
    new_n38364_, new_n38365_, new_n38366_, new_n38367_, new_n38368_,
    new_n38369_, new_n38370_, new_n38371_, new_n38372_, new_n38373_,
    new_n38374_, new_n38375_, new_n38376_, new_n38377_, new_n38378_,
    new_n38379_, new_n38380_, new_n38381_, new_n38382_, new_n38383_,
    new_n38384_, new_n38385_, new_n38386_, new_n38387_, new_n38388_,
    new_n38389_, new_n38390_, new_n38391_, new_n38392_, new_n38393_,
    new_n38394_, new_n38395_, new_n38396_, new_n38397_, new_n38398_,
    new_n38399_, new_n38400_, new_n38401_, new_n38402_, new_n38403_,
    new_n38404_, new_n38405_, new_n38406_, new_n38407_, new_n38408_,
    new_n38409_, new_n38410_, new_n38411_, new_n38412_, new_n38413_,
    new_n38414_, new_n38415_, new_n38416_, new_n38417_, new_n38418_,
    new_n38419_, new_n38420_, new_n38421_, new_n38422_, new_n38423_,
    new_n38424_, new_n38425_, new_n38426_, new_n38427_, new_n38428_,
    new_n38429_, new_n38430_, new_n38431_, new_n38432_, new_n38433_,
    new_n38434_, new_n38435_, new_n38436_, new_n38437_, new_n38438_,
    new_n38439_, new_n38440_, new_n38441_, new_n38442_, new_n38443_,
    new_n38444_, new_n38445_, new_n38446_, new_n38447_, new_n38448_,
    new_n38449_, new_n38450_, new_n38451_, new_n38452_, new_n38453_,
    new_n38454_, new_n38455_, new_n38456_, new_n38457_, new_n38458_,
    new_n38459_, new_n38460_, new_n38461_, new_n38462_, new_n38463_,
    new_n38464_, new_n38465_, new_n38466_, new_n38467_, new_n38468_,
    new_n38469_, new_n38470_, new_n38471_, new_n38472_, new_n38473_,
    new_n38474_, new_n38475_, new_n38476_, new_n38477_, new_n38478_,
    new_n38479_, new_n38480_, new_n38481_, new_n38482_, new_n38483_,
    new_n38484_, new_n38485_, new_n38486_, new_n38487_, new_n38488_,
    new_n38489_, new_n38490_, new_n38491_, new_n38492_, new_n38493_,
    new_n38494_, new_n38495_, new_n38496_, new_n38497_, new_n38498_,
    new_n38499_, new_n38500_, new_n38501_, new_n38502_, new_n38503_,
    new_n38504_, new_n38505_, new_n38506_, new_n38507_, new_n38508_,
    new_n38509_, new_n38510_, new_n38511_, new_n38512_, new_n38513_,
    new_n38514_, new_n38515_, new_n38516_, new_n38517_, new_n38518_,
    new_n38519_, new_n38520_, new_n38521_, new_n38522_, new_n38523_,
    new_n38524_, new_n38525_, new_n38526_, new_n38527_, new_n38528_,
    new_n38529_, new_n38530_, new_n38531_, new_n38532_, new_n38533_,
    new_n38534_, new_n38535_, new_n38536_, new_n38537_, new_n38538_,
    new_n38539_, new_n38540_, new_n38541_, new_n38542_, new_n38543_,
    new_n38544_, new_n38545_, new_n38546_, new_n38547_, new_n38548_,
    new_n38549_, new_n38550_, new_n38551_, new_n38552_, new_n38553_,
    new_n38554_, new_n38555_, new_n38556_, new_n38557_, new_n38558_,
    new_n38559_, new_n38560_, new_n38561_, new_n38562_, new_n38563_,
    new_n38564_, new_n38565_, new_n38566_, new_n38567_, new_n38568_,
    new_n38569_, new_n38570_, new_n38571_, new_n38572_, new_n38573_,
    new_n38574_, new_n38575_, new_n38576_, new_n38577_, new_n38578_,
    new_n38579_, new_n38580_, new_n38581_, new_n38582_, new_n38583_,
    new_n38584_, new_n38585_, new_n38586_, new_n38587_, new_n38588_,
    new_n38589_, new_n38590_, new_n38591_, new_n38592_, new_n38593_,
    new_n38594_, new_n38595_, new_n38596_, new_n38597_, new_n38598_,
    new_n38599_, new_n38600_, new_n38601_, new_n38602_, new_n38603_,
    new_n38604_, new_n38605_, new_n38606_, new_n38607_, new_n38608_,
    new_n38609_, new_n38610_, new_n38611_, new_n38612_, new_n38613_,
    new_n38614_, new_n38615_, new_n38616_, new_n38617_, new_n38618_,
    new_n38619_, new_n38620_, new_n38621_, new_n38622_, new_n38623_,
    new_n38624_, new_n38625_, new_n38626_, new_n38627_, new_n38628_,
    new_n38629_, new_n38630_, new_n38631_, new_n38632_, new_n38633_,
    new_n38634_, new_n38635_, new_n38636_, new_n38637_, new_n38638_,
    new_n38639_, new_n38640_, new_n38641_, new_n38642_, new_n38643_,
    new_n38644_, new_n38645_, new_n38646_, new_n38647_, new_n38648_,
    new_n38649_, new_n38650_, new_n38651_, new_n38652_, new_n38653_,
    new_n38654_, new_n38655_, new_n38656_, new_n38657_, new_n38658_,
    new_n38659_, new_n38660_, new_n38661_, new_n38662_, new_n38663_,
    new_n38664_, new_n38665_, new_n38666_, new_n38667_, new_n38668_,
    new_n38669_, new_n38670_, new_n38671_, new_n38672_, new_n38673_,
    new_n38674_, new_n38675_, new_n38676_, new_n38677_, new_n38678_,
    new_n38679_, new_n38680_, new_n38681_, new_n38682_, new_n38683_,
    new_n38684_, new_n38685_, new_n38686_, new_n38687_, new_n38688_,
    new_n38689_, new_n38690_, new_n38691_, new_n38692_, new_n38693_,
    new_n38694_, new_n38695_, new_n38696_, new_n38697_, new_n38698_,
    new_n38699_, new_n38700_, new_n38701_, new_n38702_, new_n38703_,
    new_n38704_, new_n38705_, new_n38706_, new_n38707_, new_n38708_,
    new_n38709_, new_n38710_, new_n38711_, new_n38712_, new_n38713_,
    new_n38714_, new_n38715_, new_n38716_, new_n38717_, new_n38718_,
    new_n38719_, new_n38720_, new_n38721_, new_n38722_, new_n38723_,
    new_n38724_, new_n38725_, new_n38726_, new_n38727_, new_n38728_,
    new_n38729_, new_n38730_, new_n38731_, new_n38732_, new_n38733_,
    new_n38734_, new_n38735_, new_n38736_, new_n38737_, new_n38738_,
    new_n38739_, new_n38740_, new_n38741_, new_n38742_, new_n38743_,
    new_n38744_, new_n38745_, new_n38746_, new_n38747_, new_n38748_,
    new_n38749_, new_n38750_, new_n38751_, new_n38752_, new_n38753_,
    new_n38754_, new_n38755_, new_n38756_, new_n38757_, new_n38758_,
    new_n38759_, new_n38760_, new_n38761_, new_n38762_, new_n38763_,
    new_n38764_, new_n38765_, new_n38766_, new_n38767_, new_n38768_,
    new_n38769_, new_n38770_, new_n38771_, new_n38772_, new_n38773_,
    new_n38774_, new_n38775_, new_n38776_, new_n38777_, new_n38778_,
    new_n38779_, new_n38780_, new_n38781_, new_n38782_, new_n38783_,
    new_n38784_, new_n38785_, new_n38786_, new_n38787_, new_n38788_,
    new_n38789_, new_n38790_, new_n38791_, new_n38792_, new_n38793_,
    new_n38794_, new_n38795_, new_n38796_, new_n38797_, new_n38798_,
    new_n38799_, new_n38800_, new_n38801_, new_n38802_, new_n38803_,
    new_n38804_, new_n38805_, new_n38806_, new_n38807_, new_n38808_,
    new_n38809_, new_n38810_, new_n38811_, new_n38812_, new_n38813_,
    new_n38814_, new_n38815_, new_n38816_, new_n38817_, new_n38818_,
    new_n38819_, new_n38820_, new_n38821_, new_n38822_, new_n38823_,
    new_n38824_, new_n38825_, new_n38826_, new_n38827_, new_n38828_,
    new_n38829_, new_n38830_, new_n38831_, new_n38832_, new_n38833_,
    new_n38834_, new_n38835_, new_n38836_, new_n38837_, new_n38838_,
    new_n38839_, new_n38840_, new_n38841_, new_n38842_, new_n38843_,
    new_n38844_, new_n38845_, new_n38846_, new_n38847_, new_n38848_,
    new_n38849_, new_n38850_, new_n38851_, new_n38852_, new_n38853_,
    new_n38854_, new_n38855_, new_n38856_, new_n38857_, new_n38858_,
    new_n38859_, new_n38860_, new_n38861_, new_n38862_, new_n38863_,
    new_n38864_, new_n38865_, new_n38866_, new_n38867_, new_n38868_,
    new_n38869_, new_n38870_, new_n38871_, new_n38872_, new_n38873_,
    new_n38874_, new_n38875_, new_n38876_, new_n38877_, new_n38878_,
    new_n38879_, new_n38880_, new_n38881_, new_n38882_, new_n38883_,
    new_n38884_, new_n38885_, new_n38886_, new_n38887_, new_n38888_,
    new_n38889_, new_n38890_, new_n38891_, new_n38892_, new_n38893_,
    new_n38894_, new_n38895_, new_n38896_, new_n38897_, new_n38898_,
    new_n38899_, new_n38900_, new_n38901_, new_n38902_, new_n38903_,
    new_n38904_, new_n38905_, new_n38906_, new_n38907_, new_n38908_,
    new_n38909_, new_n38910_, new_n38911_, new_n38912_, new_n38913_,
    new_n38914_, new_n38915_, new_n38916_, new_n38917_, new_n38918_,
    new_n38919_, new_n38920_, new_n38921_, new_n38922_, new_n38923_,
    new_n38924_, new_n38925_, new_n38926_, new_n38927_, new_n38928_,
    new_n38929_, new_n38930_, new_n38931_, new_n38932_, new_n38933_,
    new_n38934_, new_n38935_, new_n38936_, new_n38937_, new_n38938_,
    new_n38939_, new_n38940_, new_n38941_, new_n38942_, new_n38943_,
    new_n38944_, new_n38945_, new_n38946_, new_n38947_, new_n38948_,
    new_n38949_, new_n38950_, new_n38951_, new_n38952_, new_n38953_,
    new_n38954_, new_n38955_, new_n38956_, new_n38957_, new_n38958_,
    new_n38959_, new_n38960_, new_n38961_, new_n38962_, new_n38963_,
    new_n38964_, new_n38965_, new_n38966_, new_n38967_, new_n38968_,
    new_n38969_, new_n38970_, new_n38971_, new_n38972_, new_n38973_,
    new_n38974_, new_n38975_, new_n38976_, new_n38977_, new_n38978_,
    new_n38979_, new_n38980_, new_n38981_, new_n38982_, new_n38983_,
    new_n38984_, new_n38985_, new_n38986_, new_n38987_, new_n38988_,
    new_n38989_, new_n38990_, new_n38991_, new_n38992_, new_n38993_,
    new_n38994_, new_n38995_, new_n38996_, new_n38997_, new_n38998_,
    new_n38999_, new_n39000_, new_n39001_, new_n39002_, new_n39003_,
    new_n39004_, new_n39005_, new_n39006_, new_n39007_, new_n39008_,
    new_n39009_, new_n39010_, new_n39011_, new_n39012_, new_n39013_,
    new_n39014_, new_n39015_, new_n39016_, new_n39017_, new_n39018_,
    new_n39019_, new_n39020_, new_n39021_, new_n39022_, new_n39023_,
    new_n39024_, new_n39025_, new_n39026_, new_n39027_, new_n39028_,
    new_n39029_, new_n39030_, new_n39031_, new_n39032_, new_n39033_,
    new_n39034_, new_n39035_, new_n39036_, new_n39037_, new_n39038_,
    new_n39039_, new_n39040_, new_n39041_, new_n39042_, new_n39043_,
    new_n39044_, new_n39045_, new_n39046_, new_n39047_, new_n39048_,
    new_n39049_, new_n39050_, new_n39051_, new_n39052_, new_n39053_,
    new_n39054_, new_n39055_, new_n39056_, new_n39057_, new_n39058_,
    new_n39059_, new_n39060_, new_n39061_, new_n39062_, new_n39063_,
    new_n39064_, new_n39065_, new_n39066_, new_n39067_, new_n39068_,
    new_n39069_, new_n39070_, new_n39071_, new_n39072_, new_n39073_,
    new_n39074_, new_n39075_, new_n39076_, new_n39077_, new_n39078_,
    new_n39079_, new_n39080_, new_n39081_, new_n39082_, new_n39083_,
    new_n39084_, new_n39085_, new_n39086_, new_n39087_, new_n39088_,
    new_n39089_, new_n39090_, new_n39091_, new_n39092_, new_n39093_,
    new_n39094_, new_n39095_, new_n39096_, new_n39097_, new_n39098_,
    new_n39099_, new_n39100_, new_n39101_, new_n39102_, new_n39103_,
    new_n39104_, new_n39105_, new_n39106_, new_n39107_, new_n39108_,
    new_n39109_, new_n39110_, new_n39111_, new_n39112_, new_n39113_,
    new_n39114_, new_n39115_, new_n39116_, new_n39117_, new_n39118_,
    new_n39119_, new_n39120_, new_n39121_, new_n39122_, new_n39123_,
    new_n39124_, new_n39125_, new_n39126_, new_n39127_, new_n39128_,
    new_n39129_, new_n39130_, new_n39131_, new_n39132_, new_n39133_,
    new_n39134_, new_n39135_, new_n39136_, new_n39137_, new_n39138_,
    new_n39139_, new_n39140_, new_n39141_, new_n39142_, new_n39143_,
    new_n39144_, new_n39145_, new_n39146_, new_n39147_, new_n39148_,
    new_n39149_, new_n39150_, new_n39151_, new_n39152_, new_n39153_,
    new_n39154_, new_n39155_, new_n39156_, new_n39157_, new_n39158_,
    new_n39159_, new_n39160_, new_n39161_, new_n39162_, new_n39163_,
    new_n39164_, new_n39165_, new_n39166_, new_n39167_, new_n39168_,
    new_n39169_, new_n39170_, new_n39171_, new_n39172_, new_n39173_,
    new_n39174_, new_n39175_, new_n39176_, new_n39177_, new_n39178_,
    new_n39179_, new_n39180_, new_n39181_, new_n39182_, new_n39183_,
    new_n39184_, new_n39185_, new_n39186_, new_n39187_, new_n39188_,
    new_n39189_, new_n39190_, new_n39191_, new_n39192_, new_n39193_,
    new_n39194_, new_n39195_, new_n39196_, new_n39197_, new_n39198_,
    new_n39199_, new_n39200_, new_n39201_, new_n39202_, new_n39203_,
    new_n39204_, new_n39205_, new_n39206_, new_n39207_, new_n39208_,
    new_n39209_, new_n39210_, new_n39211_, new_n39212_, new_n39213_,
    new_n39214_, new_n39215_, new_n39216_, new_n39217_, new_n39218_,
    new_n39219_, new_n39220_, new_n39221_, new_n39222_, new_n39223_,
    new_n39224_, new_n39225_, new_n39226_, new_n39227_, new_n39228_,
    new_n39229_, new_n39230_, new_n39231_, new_n39232_, new_n39233_,
    new_n39234_, new_n39235_, new_n39236_, new_n39237_, new_n39238_,
    new_n39239_, new_n39240_, new_n39241_, new_n39242_, new_n39243_,
    new_n39244_, new_n39245_, new_n39246_, new_n39247_, new_n39248_,
    new_n39249_, new_n39250_, new_n39251_, new_n39252_, new_n39253_,
    new_n39254_, new_n39255_, new_n39256_, new_n39257_, new_n39258_,
    new_n39259_, new_n39260_, new_n39261_, new_n39262_, new_n39263_,
    new_n39264_, new_n39265_, new_n39266_, new_n39267_, new_n39268_,
    new_n39269_, new_n39270_, new_n39271_, new_n39272_, new_n39273_,
    new_n39274_, new_n39275_, new_n39276_, new_n39277_, new_n39278_,
    new_n39279_, new_n39280_, new_n39281_, new_n39282_, new_n39283_,
    new_n39284_, new_n39285_, new_n39286_, new_n39287_, new_n39288_,
    new_n39289_, new_n39290_, new_n39291_, new_n39292_, new_n39293_,
    new_n39294_, new_n39295_, new_n39296_, new_n39297_, new_n39298_,
    new_n39299_, new_n39300_, new_n39301_, new_n39302_, new_n39303_,
    new_n39304_, new_n39305_, new_n39306_, new_n39307_, new_n39308_,
    new_n39309_, new_n39310_, new_n39311_, new_n39312_, new_n39313_,
    new_n39314_, new_n39315_, new_n39316_, new_n39317_, new_n39318_,
    new_n39319_, new_n39320_, new_n39321_, new_n39322_, new_n39323_,
    new_n39324_, new_n39325_, new_n39326_, new_n39327_, new_n39328_,
    new_n39329_, new_n39330_, new_n39331_, new_n39332_, new_n39333_,
    new_n39334_, new_n39335_, new_n39336_, new_n39337_, new_n39338_,
    new_n39339_, new_n39340_, new_n39341_, new_n39342_, new_n39343_,
    new_n39344_, new_n39345_, new_n39346_, new_n39347_, new_n39348_,
    new_n39349_, new_n39350_, new_n39351_, new_n39352_, new_n39353_,
    new_n39354_, new_n39355_, new_n39356_, new_n39357_, new_n39358_,
    new_n39359_, new_n39360_, new_n39361_, new_n39362_, new_n39363_,
    new_n39364_, new_n39365_, new_n39366_, new_n39367_, new_n39368_,
    new_n39369_, new_n39370_, new_n39371_, new_n39372_, new_n39373_,
    new_n39374_, new_n39375_, new_n39376_, new_n39377_, new_n39378_,
    new_n39379_, new_n39380_, new_n39381_, new_n39382_, new_n39383_,
    new_n39384_, new_n39385_, new_n39386_, new_n39387_, new_n39388_,
    new_n39389_, new_n39390_, new_n39391_, new_n39392_, new_n39393_,
    new_n39394_, new_n39395_, new_n39396_, new_n39397_, new_n39398_,
    new_n39399_, new_n39400_, new_n39401_, new_n39402_, new_n39403_,
    new_n39404_, new_n39405_, new_n39406_, new_n39407_, new_n39408_,
    new_n39409_, new_n39410_, new_n39411_, new_n39412_, new_n39413_,
    new_n39414_, new_n39415_, new_n39416_, new_n39417_, new_n39418_,
    new_n39419_, new_n39420_, new_n39421_, new_n39422_, new_n39423_,
    new_n39424_, new_n39425_, new_n39426_, new_n39427_, new_n39428_,
    new_n39429_, new_n39430_, new_n39431_, new_n39432_, new_n39433_,
    new_n39434_, new_n39435_, new_n39436_, new_n39437_, new_n39438_,
    new_n39439_, new_n39440_, new_n39441_, new_n39442_, new_n39443_,
    new_n39444_, new_n39445_, new_n39446_, new_n39447_, new_n39448_,
    new_n39449_, new_n39450_, new_n39451_, new_n39452_, new_n39453_,
    new_n39454_, new_n39455_, new_n39456_, new_n39457_, new_n39458_,
    new_n39459_, new_n39460_, new_n39461_, new_n39462_, new_n39463_,
    new_n39464_, new_n39465_, new_n39466_, new_n39467_, new_n39468_,
    new_n39469_, new_n39470_, new_n39471_, new_n39472_, new_n39473_,
    new_n39474_, new_n39475_, new_n39476_, new_n39477_, new_n39478_,
    new_n39479_, new_n39480_, new_n39481_, new_n39482_, new_n39483_,
    new_n39484_, new_n39485_, new_n39486_, new_n39487_, new_n39488_,
    new_n39489_, new_n39490_, new_n39491_, new_n39492_, new_n39493_,
    new_n39494_, new_n39495_, new_n39496_, new_n39497_, new_n39498_,
    new_n39499_, new_n39500_, new_n39501_, new_n39502_, new_n39503_,
    new_n39504_, new_n39505_, new_n39506_, new_n39507_, new_n39508_,
    new_n39509_, new_n39510_, new_n39511_, new_n39512_, new_n39513_,
    new_n39514_, new_n39515_, new_n39516_, new_n39517_, new_n39518_,
    new_n39519_, new_n39520_, new_n39521_, new_n39522_, new_n39523_,
    new_n39524_, new_n39525_, new_n39526_, new_n39527_, new_n39528_,
    new_n39529_, new_n39530_, new_n39531_, new_n39532_, new_n39533_,
    new_n39534_, new_n39535_, new_n39536_, new_n39537_, new_n39538_,
    new_n39539_, new_n39540_, new_n39541_, new_n39542_, new_n39543_,
    new_n39544_, new_n39545_, new_n39546_, new_n39547_, new_n39548_,
    new_n39549_, new_n39550_, new_n39551_, new_n39552_, new_n39553_,
    new_n39554_, new_n39555_, new_n39556_, new_n39557_, new_n39558_,
    new_n39559_, new_n39560_, new_n39561_, new_n39562_, new_n39563_,
    new_n39564_, new_n39565_, new_n39566_, new_n39567_, new_n39568_,
    new_n39569_, new_n39570_, new_n39571_, new_n39572_, new_n39573_,
    new_n39574_, new_n39575_, new_n39576_, new_n39577_, new_n39578_,
    new_n39579_, new_n39580_, new_n39581_, new_n39582_, new_n39583_,
    new_n39584_, new_n39585_, new_n39586_, new_n39587_, new_n39588_,
    new_n39589_, new_n39590_, new_n39591_, new_n39592_, new_n39593_,
    new_n39594_, new_n39595_, new_n39596_, new_n39597_, new_n39598_,
    new_n39599_, new_n39600_, new_n39601_, new_n39602_, new_n39603_,
    new_n39604_, new_n39605_, new_n39606_, new_n39607_, new_n39608_,
    new_n39609_, new_n39610_, new_n39611_, new_n39612_, new_n39613_,
    new_n39614_, new_n39615_, new_n39616_, new_n39617_, new_n39618_,
    new_n39619_, new_n39620_, new_n39621_, new_n39622_, new_n39623_,
    new_n39624_, new_n39625_, new_n39626_, new_n39627_, new_n39628_,
    new_n39629_, new_n39630_, new_n39631_, new_n39632_, new_n39633_,
    new_n39634_, new_n39635_, new_n39636_, new_n39637_, new_n39638_,
    new_n39639_, new_n39640_, new_n39641_, new_n39642_, new_n39643_,
    new_n39644_, new_n39645_, new_n39646_, new_n39647_, new_n39648_,
    new_n39649_, new_n39650_, new_n39651_, new_n39652_, new_n39653_,
    new_n39654_, new_n39655_, new_n39656_, new_n39657_, new_n39658_,
    new_n39659_, new_n39660_, new_n39661_, new_n39662_, new_n39663_,
    new_n39664_, new_n39665_, new_n39666_, new_n39667_, new_n39668_,
    new_n39669_, new_n39670_, new_n39671_, new_n39672_, new_n39673_,
    new_n39674_, new_n39675_, new_n39676_, new_n39677_, new_n39678_,
    new_n39679_, new_n39680_, new_n39681_, new_n39682_, new_n39683_,
    new_n39684_, new_n39685_, new_n39686_, new_n39687_, new_n39688_,
    new_n39689_, new_n39690_, new_n39691_, new_n39692_, new_n39693_,
    new_n39694_, new_n39695_, new_n39696_, new_n39697_, new_n39698_,
    new_n39699_, new_n39700_, new_n39701_, new_n39702_, new_n39703_,
    new_n39704_, new_n39705_, new_n39706_, new_n39707_, new_n39708_,
    new_n39709_, new_n39710_, new_n39711_, new_n39712_, new_n39713_,
    new_n39714_, new_n39715_, new_n39716_, new_n39717_, new_n39718_,
    new_n39719_, new_n39720_, new_n39721_, new_n39722_, new_n39723_,
    new_n39724_, new_n39725_, new_n39726_, new_n39727_, new_n39728_,
    new_n39729_, new_n39730_, new_n39731_, new_n39732_, new_n39733_,
    new_n39734_, new_n39735_, new_n39736_, new_n39737_, new_n39738_,
    new_n39739_, new_n39740_, new_n39741_, new_n39742_, new_n39743_,
    new_n39744_, new_n39745_, new_n39746_, new_n39747_, new_n39748_,
    new_n39749_, new_n39750_, new_n39751_, new_n39752_, new_n39753_,
    new_n39754_, new_n39755_, new_n39756_, new_n39757_, new_n39758_,
    new_n39759_, new_n39760_, new_n39761_, new_n39762_, new_n39763_,
    new_n39764_, new_n39765_, new_n39766_, new_n39767_, new_n39768_,
    new_n39769_, new_n39770_, new_n39771_, new_n39772_, new_n39773_,
    new_n39774_, new_n39775_, new_n39776_, new_n39777_, new_n39778_,
    new_n39779_, new_n39780_, new_n39781_, new_n39782_, new_n39783_,
    new_n39784_, new_n39785_, new_n39786_, new_n39787_, new_n39788_,
    new_n39789_, new_n39790_, new_n39791_, new_n39792_, new_n39793_,
    new_n39794_, new_n39795_, new_n39796_, new_n39797_, new_n39798_,
    new_n39799_, new_n39800_, new_n39801_, new_n39802_, new_n39803_,
    new_n39804_, new_n39805_, new_n39806_, new_n39807_, new_n39808_,
    new_n39809_, new_n39810_, new_n39811_, new_n39812_, new_n39813_,
    new_n39814_, new_n39815_, new_n39816_, new_n39817_, new_n39818_,
    new_n39819_, new_n39820_, new_n39821_, new_n39822_, new_n39823_,
    new_n39824_, new_n39825_, new_n39826_, new_n39827_, new_n39828_,
    new_n39829_, new_n39830_, new_n39831_, new_n39832_, new_n39833_,
    new_n39834_, new_n39835_, new_n39836_, new_n39837_, new_n39838_,
    new_n39839_, new_n39840_, new_n39841_, new_n39842_, new_n39843_,
    new_n39844_, new_n39845_, new_n39846_, new_n39847_, new_n39848_,
    new_n39849_, new_n39850_, new_n39851_, new_n39852_, new_n39853_,
    new_n39854_, new_n39855_, new_n39856_, new_n39857_, new_n39858_,
    new_n39859_, new_n39860_, new_n39861_, new_n39862_, new_n39863_,
    new_n39864_, new_n39865_, new_n39866_, new_n39867_, new_n39868_,
    new_n39869_, new_n39870_, new_n39871_, new_n39872_, new_n39873_,
    new_n39874_, new_n39875_, new_n39876_, new_n39877_, new_n39878_,
    new_n39879_, new_n39880_, new_n39881_, new_n39882_, new_n39883_,
    new_n39884_, new_n39885_, new_n39886_, new_n39887_, new_n39888_,
    new_n39889_, new_n39890_, new_n39891_, new_n39892_, new_n39893_,
    new_n39894_, new_n39895_, new_n39896_, new_n39897_, new_n39898_,
    new_n39899_, new_n39900_, new_n39901_, new_n39902_, new_n39903_,
    new_n39904_, new_n39905_, new_n39906_, new_n39907_, new_n39908_,
    new_n39909_, new_n39910_, new_n39911_, new_n39912_, new_n39913_,
    new_n39914_, new_n39915_, new_n39916_, new_n39917_, new_n39918_,
    new_n39919_, new_n39920_, new_n39921_, new_n39922_, new_n39923_,
    new_n39924_, new_n39925_, new_n39926_, new_n39927_, new_n39928_,
    new_n39929_, new_n39930_, new_n39931_, new_n39932_, new_n39933_,
    new_n39934_, new_n39935_, new_n39936_, new_n39937_, new_n39938_,
    new_n39939_, new_n39940_, new_n39941_, new_n39942_, new_n39943_,
    new_n39944_, new_n39945_, new_n39946_, new_n39947_, new_n39948_,
    new_n39949_, new_n39950_, new_n39951_, new_n39952_, new_n39953_,
    new_n39954_, new_n39955_, new_n39956_, new_n39957_, new_n39958_,
    new_n39959_, new_n39960_, new_n39961_, new_n39962_, new_n39963_,
    new_n39964_, new_n39965_, new_n39966_, new_n39967_, new_n39968_,
    new_n39969_, new_n39970_, new_n39971_, new_n39972_, new_n39973_,
    new_n39974_, new_n39975_, new_n39976_, new_n39977_, new_n39978_,
    new_n39979_, new_n39980_, new_n39981_, new_n39982_, new_n39983_,
    new_n39984_, new_n39985_, new_n39986_, new_n39987_, new_n39988_,
    new_n39989_, new_n39990_, new_n39991_, new_n39992_, new_n39993_,
    new_n39994_, new_n39995_, new_n39996_, new_n39997_, new_n39998_,
    new_n39999_, new_n40000_, new_n40001_, new_n40002_, new_n40003_,
    new_n40004_, new_n40005_, new_n40006_, new_n40007_, new_n40008_,
    new_n40009_, new_n40010_, new_n40011_, new_n40012_, new_n40013_,
    new_n40014_, new_n40015_, new_n40016_, new_n40017_, new_n40018_,
    new_n40019_, new_n40020_, new_n40021_, new_n40022_, new_n40023_,
    new_n40024_, new_n40025_, new_n40026_, new_n40027_, new_n40028_,
    new_n40029_, new_n40030_, new_n40031_, new_n40032_, new_n40033_,
    new_n40034_, new_n40035_, new_n40036_, new_n40037_, new_n40038_,
    new_n40039_, new_n40040_, new_n40041_, new_n40042_, new_n40043_,
    new_n40044_, new_n40045_, new_n40046_, new_n40047_, new_n40048_,
    new_n40049_, new_n40050_, new_n40051_, new_n40052_, new_n40053_,
    new_n40054_, new_n40055_, new_n40056_, new_n40057_, new_n40058_,
    new_n40059_, new_n40060_, new_n40061_, new_n40062_, new_n40063_,
    new_n40064_, new_n40065_, new_n40066_, new_n40067_, new_n40068_,
    new_n40069_, new_n40070_, new_n40071_, new_n40072_, new_n40073_,
    new_n40074_, new_n40075_, new_n40076_, new_n40077_, new_n40078_,
    new_n40079_, new_n40080_, new_n40081_, new_n40082_, new_n40083_,
    new_n40084_, new_n40085_, new_n40086_, new_n40087_, new_n40088_,
    new_n40089_, new_n40090_, new_n40091_, new_n40092_, new_n40093_,
    new_n40094_, new_n40095_, new_n40096_, new_n40097_, new_n40098_,
    new_n40099_, new_n40100_, new_n40101_, new_n40102_, new_n40103_,
    new_n40104_, new_n40105_, new_n40106_, new_n40107_, new_n40108_,
    new_n40109_, new_n40110_, new_n40111_, new_n40112_, new_n40113_,
    new_n40114_, new_n40115_, new_n40116_, new_n40117_, new_n40118_,
    new_n40119_, new_n40120_, new_n40121_, new_n40122_, new_n40123_,
    new_n40124_, new_n40125_, new_n40126_, new_n40127_, new_n40128_,
    new_n40129_, new_n40130_, new_n40131_, new_n40132_, new_n40133_,
    new_n40134_, new_n40135_, new_n40136_, new_n40137_, new_n40138_,
    new_n40139_, new_n40140_, new_n40141_, new_n40142_, new_n40143_,
    new_n40144_, new_n40145_, new_n40146_, new_n40147_, new_n40148_,
    new_n40149_, new_n40150_, new_n40151_, new_n40152_, new_n40153_,
    new_n40154_, new_n40155_, new_n40156_, new_n40157_, new_n40158_,
    new_n40159_, new_n40160_, new_n40161_, new_n40162_, new_n40163_,
    new_n40164_, new_n40165_, new_n40166_, new_n40167_, new_n40168_,
    new_n40169_, new_n40170_, new_n40171_, new_n40172_, new_n40173_,
    new_n40174_, new_n40175_, new_n40176_, new_n40177_, new_n40178_,
    new_n40179_, new_n40180_, new_n40181_, new_n40182_, new_n40183_,
    new_n40184_, new_n40185_, new_n40186_, new_n40187_, new_n40188_,
    new_n40189_, new_n40190_, new_n40191_, new_n40192_, new_n40193_,
    new_n40194_, new_n40195_, new_n40196_, new_n40197_, new_n40198_,
    new_n40199_, new_n40200_, new_n40201_, new_n40202_, new_n40203_,
    new_n40204_, new_n40205_, new_n40206_, new_n40207_, new_n40208_,
    new_n40209_, new_n40210_, new_n40211_, new_n40212_, new_n40213_,
    new_n40214_, new_n40215_, new_n40216_, new_n40217_, new_n40218_,
    new_n40219_, new_n40220_, new_n40221_, new_n40222_, new_n40223_,
    new_n40224_, new_n40225_, new_n40226_, new_n40227_, new_n40228_,
    new_n40229_, new_n40230_, new_n40231_, new_n40232_, new_n40233_,
    new_n40234_, new_n40235_, new_n40236_, new_n40237_, new_n40238_,
    new_n40239_, new_n40240_, new_n40241_, new_n40242_, new_n40243_,
    new_n40244_, new_n40245_, new_n40246_, new_n40247_, new_n40248_,
    new_n40249_, new_n40250_, new_n40251_, new_n40252_, new_n40253_,
    new_n40254_, new_n40255_, new_n40256_, new_n40257_, new_n40258_,
    new_n40259_, new_n40260_, new_n40261_, new_n40262_, new_n40263_,
    new_n40264_, new_n40265_, new_n40266_, new_n40267_, new_n40268_,
    new_n40269_, new_n40270_, new_n40271_, new_n40272_, new_n40273_,
    new_n40274_, new_n40275_, new_n40276_, new_n40277_, new_n40278_,
    new_n40279_, new_n40280_, new_n40281_, new_n40282_, new_n40283_,
    new_n40284_, new_n40285_, new_n40286_, new_n40287_, new_n40288_,
    new_n40289_, new_n40290_, new_n40291_, new_n40292_, new_n40293_,
    new_n40294_, new_n40295_, new_n40296_, new_n40297_, new_n40298_,
    new_n40299_, new_n40300_, new_n40301_, new_n40302_, new_n40303_,
    new_n40304_, new_n40305_, new_n40306_, new_n40307_, new_n40308_,
    new_n40309_, new_n40310_, new_n40311_, new_n40312_, new_n40313_,
    new_n40314_, new_n40315_, new_n40316_, new_n40317_, new_n40318_,
    new_n40319_, new_n40320_, new_n40321_, new_n40322_, new_n40323_,
    new_n40324_, new_n40325_, new_n40326_, new_n40327_, new_n40328_,
    new_n40329_, new_n40330_, new_n40331_, new_n40332_, new_n40333_,
    new_n40334_, new_n40335_, new_n40336_, new_n40337_, new_n40338_,
    new_n40339_, new_n40340_, new_n40341_, new_n40342_, new_n40343_,
    new_n40344_, new_n40345_, new_n40346_, new_n40347_, new_n40348_,
    new_n40349_, new_n40350_, new_n40351_, new_n40352_, new_n40353_,
    new_n40354_, new_n40355_, new_n40356_, new_n40357_, new_n40358_,
    new_n40359_, new_n40360_, new_n40361_, new_n40362_, new_n40363_,
    new_n40364_, new_n40365_, new_n40366_, new_n40367_, new_n40368_,
    new_n40369_, new_n40370_, new_n40371_, new_n40372_, new_n40373_,
    new_n40374_, new_n40375_, new_n40376_, new_n40377_, new_n40378_,
    new_n40379_, new_n40380_, new_n40381_, new_n40382_, new_n40383_,
    new_n40384_, new_n40385_, new_n40386_, new_n40387_, new_n40388_,
    new_n40389_, new_n40390_, new_n40391_, new_n40392_, new_n40393_,
    new_n40394_, new_n40395_, new_n40396_, new_n40397_, new_n40398_,
    new_n40399_, new_n40400_, new_n40401_, new_n40402_, new_n40403_,
    new_n40404_, new_n40405_, new_n40406_, new_n40407_, new_n40408_,
    new_n40409_, new_n40410_, new_n40411_, new_n40412_, new_n40413_,
    new_n40414_, new_n40415_, new_n40416_, new_n40417_, new_n40418_,
    new_n40419_, new_n40420_, new_n40421_, new_n40422_, new_n40423_,
    new_n40424_, new_n40425_, new_n40426_, new_n40427_, new_n40428_,
    new_n40429_, new_n40430_, new_n40431_, new_n40432_, new_n40433_,
    new_n40434_, new_n40435_, new_n40436_, new_n40437_, new_n40438_,
    new_n40439_, new_n40440_, new_n40441_, new_n40442_, new_n40443_,
    new_n40444_, new_n40445_, new_n40446_, new_n40447_, new_n40448_,
    new_n40449_, new_n40450_, new_n40451_, new_n40452_, new_n40453_,
    new_n40454_, new_n40455_, new_n40456_, new_n40457_, new_n40458_,
    new_n40459_, new_n40460_, new_n40461_, new_n40462_, new_n40463_,
    new_n40464_, new_n40465_, new_n40466_, new_n40467_, new_n40468_,
    new_n40469_, new_n40470_, new_n40471_, new_n40472_, new_n40473_,
    new_n40474_, new_n40475_, new_n40476_, new_n40477_, new_n40478_,
    new_n40479_, new_n40480_, new_n40481_, new_n40482_, new_n40483_,
    new_n40484_, new_n40485_, new_n40486_, new_n40487_, new_n40488_,
    new_n40489_, new_n40490_, new_n40491_, new_n40492_, new_n40493_,
    new_n40494_, new_n40495_, new_n40496_, new_n40497_, new_n40498_,
    new_n40499_, new_n40500_, new_n40501_, new_n40502_, new_n40503_,
    new_n40504_, new_n40505_, new_n40506_, new_n40507_, new_n40508_,
    new_n40509_, new_n40510_, new_n40511_, new_n40512_, new_n40513_,
    new_n40514_, new_n40515_, new_n40516_, new_n40517_, new_n40518_,
    new_n40519_, new_n40520_, new_n40521_, new_n40522_, new_n40523_,
    new_n40524_, new_n40525_, new_n40526_, new_n40527_, new_n40528_,
    new_n40529_, new_n40530_, new_n40531_, new_n40532_, new_n40533_,
    new_n40534_, new_n40535_, new_n40536_, new_n40537_, new_n40538_,
    new_n40539_, new_n40540_, new_n40541_, new_n40542_, new_n40543_,
    new_n40544_, new_n40545_, new_n40546_, new_n40547_, new_n40548_,
    new_n40549_, new_n40550_, new_n40551_, new_n40552_, new_n40553_,
    new_n40554_, new_n40555_, new_n40556_, new_n40557_, new_n40558_,
    new_n40559_, new_n40560_, new_n40561_, new_n40562_, new_n40563_,
    new_n40564_, new_n40565_, new_n40566_, new_n40567_, new_n40568_,
    new_n40569_, new_n40570_, new_n40571_, new_n40572_, new_n40573_,
    new_n40574_, new_n40575_, new_n40576_, new_n40577_, new_n40578_,
    new_n40579_, new_n40580_, new_n40581_, new_n40582_, new_n40583_,
    new_n40584_, new_n40585_, new_n40586_, new_n40587_, new_n40588_,
    new_n40589_, new_n40590_, new_n40591_, new_n40592_, new_n40593_,
    new_n40594_, new_n40595_, new_n40596_, new_n40597_, new_n40598_,
    new_n40599_, new_n40600_, new_n40601_, new_n40602_, new_n40603_,
    new_n40604_, new_n40605_, new_n40606_, new_n40607_, new_n40608_,
    new_n40609_, new_n40610_, new_n40611_, new_n40612_, new_n40613_,
    new_n40614_, new_n40615_, new_n40616_, new_n40617_, new_n40618_,
    new_n40619_, new_n40620_, new_n40621_, new_n40622_, new_n40623_,
    new_n40624_, new_n40625_, new_n40626_, new_n40627_, new_n40628_,
    new_n40629_, new_n40630_, new_n40631_, new_n40632_, new_n40633_,
    new_n40634_, new_n40635_, new_n40636_, new_n40637_, new_n40638_,
    new_n40639_, new_n40640_, new_n40641_, new_n40642_, new_n40643_,
    new_n40644_, new_n40645_, new_n40646_, new_n40647_, new_n40648_,
    new_n40649_, new_n40650_, new_n40651_, new_n40652_, new_n40653_,
    new_n40654_, new_n40655_, new_n40656_, new_n40657_, new_n40658_,
    new_n40659_, new_n40660_, new_n40661_, new_n40662_, new_n40663_,
    new_n40664_, new_n40665_, new_n40666_, new_n40667_, new_n40668_,
    new_n40669_, new_n40670_, new_n40671_, new_n40672_, new_n40673_,
    new_n40674_, new_n40675_, new_n40676_, new_n40677_, new_n40678_,
    new_n40679_, new_n40680_, new_n40681_, new_n40682_, new_n40683_,
    new_n40684_, new_n40685_, new_n40686_, new_n40687_, new_n40688_,
    new_n40689_, new_n40690_, new_n40691_, new_n40692_, new_n40693_,
    new_n40694_, new_n40695_, new_n40696_, new_n40697_, new_n40698_,
    new_n40699_, new_n40700_, new_n40701_, new_n40702_, new_n40703_,
    new_n40704_, new_n40705_, new_n40706_, new_n40707_, new_n40708_,
    new_n40709_, new_n40710_, new_n40711_, new_n40712_, new_n40713_,
    new_n40714_, new_n40715_, new_n40716_, new_n40717_, new_n40718_,
    new_n40719_, new_n40720_, new_n40721_, new_n40722_, new_n40723_,
    new_n40724_, new_n40725_, new_n40726_, new_n40727_, new_n40728_,
    new_n40729_, new_n40730_, new_n40731_, new_n40732_, new_n40733_,
    new_n40734_, new_n40735_, new_n40736_, new_n40737_, new_n40738_,
    new_n40739_, new_n40740_, new_n40741_, new_n40742_, new_n40743_,
    new_n40744_, new_n40745_, new_n40746_, new_n40747_, new_n40748_,
    new_n40749_, new_n40750_, new_n40751_, new_n40752_, new_n40753_,
    new_n40754_, new_n40755_, new_n40756_, new_n40757_, new_n40758_,
    new_n40759_, new_n40760_, new_n40761_, new_n40762_, new_n40763_,
    new_n40764_, new_n40765_, new_n40766_, new_n40767_, new_n40768_,
    new_n40769_, new_n40770_, new_n40771_, new_n40772_, new_n40773_,
    new_n40774_, new_n40775_, new_n40776_, new_n40777_, new_n40778_,
    new_n40779_, new_n40780_, new_n40781_, new_n40782_, new_n40783_,
    new_n40784_, new_n40785_, new_n40786_, new_n40787_, new_n40788_,
    new_n40789_, new_n40790_, new_n40791_, new_n40792_, new_n40793_,
    new_n40794_, new_n40795_, new_n40796_, new_n40797_, new_n40798_,
    new_n40799_, new_n40800_, new_n40801_, new_n40802_, new_n40803_,
    new_n40804_, new_n40805_, new_n40806_, new_n40807_, new_n40808_,
    new_n40809_, new_n40810_, new_n40811_, new_n40812_, new_n40813_,
    new_n40814_, new_n40815_, new_n40816_, new_n40817_, new_n40818_,
    new_n40819_, new_n40820_, new_n40821_, new_n40822_, new_n40823_,
    new_n40824_, new_n40825_, new_n40826_, new_n40827_, new_n40828_,
    new_n40829_, new_n40830_, new_n40831_, new_n40832_, new_n40833_,
    new_n40834_, new_n40835_, new_n40836_, new_n40837_, new_n40838_,
    new_n40839_, new_n40840_, new_n40841_, new_n40842_, new_n40843_,
    new_n40844_, new_n40845_, new_n40846_, new_n40847_, new_n40848_,
    new_n40849_, new_n40850_, new_n40851_, new_n40852_, new_n40853_,
    new_n40854_, new_n40855_, new_n40856_, new_n40857_, new_n40858_,
    new_n40859_, new_n40860_, new_n40861_, new_n40862_, new_n40863_,
    new_n40864_, new_n40865_, new_n40866_, new_n40867_, new_n40868_,
    new_n40869_, new_n40870_, new_n40871_, new_n40872_, new_n40873_,
    new_n40874_, new_n40875_, new_n40876_, new_n40877_, new_n40878_,
    new_n40879_, new_n40880_, new_n40881_, new_n40882_, new_n40883_,
    new_n40884_, new_n40885_, new_n40886_, new_n40887_, new_n40888_,
    new_n40889_, new_n40890_, new_n40891_, new_n40892_, new_n40893_,
    new_n40894_, new_n40895_, new_n40896_, new_n40897_, new_n40898_,
    new_n40899_, new_n40900_, new_n40901_, new_n40902_, new_n40903_,
    new_n40904_, new_n40905_, new_n40906_, new_n40907_, new_n40908_,
    new_n40909_, new_n40910_, new_n40911_, new_n40912_, new_n40913_,
    new_n40914_, new_n40915_, new_n40916_, new_n40917_, new_n40918_,
    new_n40919_, new_n40920_, new_n40921_, new_n40922_, new_n40923_,
    new_n40924_, new_n40925_, new_n40926_, new_n40927_, new_n40928_,
    new_n40929_, new_n40930_, new_n40931_, new_n40932_, new_n40933_,
    new_n40934_, new_n40935_, new_n40936_, new_n40937_, new_n40938_,
    new_n40939_, new_n40940_, new_n40941_, new_n40942_, new_n40943_,
    new_n40944_, new_n40945_, new_n40946_, new_n40947_, new_n40948_,
    new_n40949_, new_n40950_, new_n40951_, new_n40952_, new_n40953_,
    new_n40954_, new_n40955_, new_n40956_, new_n40957_, new_n40958_,
    new_n40959_, new_n40960_, new_n40961_, new_n40962_, new_n40963_,
    new_n40964_, new_n40965_, new_n40966_, new_n40967_, new_n40968_,
    new_n40969_, new_n40970_, new_n40971_, new_n40972_, new_n40973_,
    new_n40974_, new_n40975_, new_n40976_, new_n40977_, new_n40978_,
    new_n40979_, new_n40980_, new_n40981_, new_n40982_, new_n40983_,
    new_n40984_, new_n40985_, new_n40986_, new_n40987_, new_n40988_,
    new_n40989_, new_n40990_, new_n40991_, new_n40992_, new_n40993_,
    new_n40994_, new_n40995_, new_n40996_, new_n40997_, new_n40998_,
    new_n40999_, new_n41000_, new_n41001_, new_n41002_, new_n41003_,
    new_n41004_, new_n41005_, new_n41006_, new_n41007_, new_n41008_,
    new_n41009_, new_n41010_, new_n41011_, new_n41012_, new_n41013_,
    new_n41014_, new_n41015_, new_n41016_, new_n41017_, new_n41018_,
    new_n41019_, new_n41020_, new_n41021_, new_n41022_, new_n41023_,
    new_n41024_, new_n41025_, new_n41026_, new_n41027_, new_n41028_,
    new_n41029_, new_n41030_, new_n41031_, new_n41032_, new_n41033_,
    new_n41034_, new_n41035_, new_n41036_, new_n41037_, new_n41038_,
    new_n41039_, new_n41040_, new_n41041_, new_n41042_, new_n41043_,
    new_n41044_, new_n41045_, new_n41046_, new_n41047_, new_n41048_,
    new_n41049_, new_n41050_, new_n41051_, new_n41052_, new_n41053_,
    new_n41054_, new_n41055_, new_n41056_, new_n41057_, new_n41058_,
    new_n41059_, new_n41060_, new_n41061_, new_n41062_, new_n41063_,
    new_n41064_, new_n41065_, new_n41066_, new_n41067_, new_n41068_,
    new_n41069_, new_n41070_, new_n41071_, new_n41072_, new_n41073_,
    new_n41074_, new_n41075_, new_n41076_, new_n41077_, new_n41078_,
    new_n41079_, new_n41080_, new_n41081_, new_n41082_, new_n41083_,
    new_n41084_, new_n41085_, new_n41086_, new_n41087_, new_n41088_,
    new_n41089_, new_n41090_, new_n41091_, new_n41092_, new_n41093_,
    new_n41094_, new_n41095_, new_n41096_, new_n41097_, new_n41098_,
    new_n41099_, new_n41100_, new_n41101_, new_n41102_, new_n41103_,
    new_n41104_, new_n41105_, new_n41106_, new_n41107_, new_n41108_,
    new_n41109_, new_n41110_, new_n41111_, new_n41112_, new_n41113_,
    new_n41114_, new_n41115_, new_n41116_, new_n41117_, new_n41118_,
    new_n41119_, new_n41120_, new_n41121_, new_n41122_, new_n41123_,
    new_n41124_, new_n41125_, new_n41126_, new_n41127_, new_n41128_,
    new_n41129_, new_n41130_, new_n41131_, new_n41132_, new_n41133_,
    new_n41134_, new_n41135_, new_n41136_, new_n41137_, new_n41138_,
    new_n41139_, new_n41140_, new_n41141_, new_n41142_, new_n41143_,
    new_n41144_, new_n41145_, new_n41146_, new_n41147_, new_n41148_,
    new_n41149_, new_n41150_, new_n41151_, new_n41152_, new_n41153_,
    new_n41154_, new_n41155_, new_n41156_, new_n41157_, new_n41158_,
    new_n41159_, new_n41160_, new_n41161_, new_n41162_, new_n41163_,
    new_n41164_, new_n41165_, new_n41166_, new_n41167_, new_n41168_,
    new_n41169_, new_n41170_, new_n41171_, new_n41172_, new_n41173_,
    new_n41174_, new_n41175_, new_n41176_, new_n41177_, new_n41178_,
    new_n41179_, new_n41180_, new_n41181_, new_n41182_, new_n41183_,
    new_n41184_, new_n41185_, new_n41186_, new_n41187_, new_n41188_,
    new_n41189_, new_n41190_, new_n41191_, new_n41192_, new_n41193_,
    new_n41194_, new_n41195_, new_n41196_, new_n41197_, new_n41198_,
    new_n41199_, new_n41200_, new_n41201_, new_n41202_, new_n41203_,
    new_n41204_, new_n41205_, new_n41206_, new_n41207_, new_n41208_,
    new_n41209_, new_n41210_, new_n41211_, new_n41212_, new_n41213_,
    new_n41214_, new_n41215_, new_n41216_, new_n41217_, new_n41218_,
    new_n41219_, new_n41220_, new_n41221_, new_n41222_, new_n41223_,
    new_n41224_, new_n41225_, new_n41226_, new_n41227_, new_n41228_,
    new_n41229_, new_n41230_, new_n41231_, new_n41232_, new_n41233_,
    new_n41234_, new_n41235_, new_n41236_, new_n41237_, new_n41238_,
    new_n41239_, new_n41240_, new_n41241_, new_n41242_, new_n41243_,
    new_n41244_, new_n41245_, new_n41246_, new_n41247_, new_n41248_,
    new_n41249_, new_n41250_, new_n41251_, new_n41252_, new_n41253_,
    new_n41254_, new_n41255_, new_n41256_, new_n41257_, new_n41258_,
    new_n41259_, new_n41260_, new_n41261_, new_n41262_, new_n41263_,
    new_n41264_, new_n41265_, new_n41266_, new_n41267_, new_n41268_,
    new_n41269_, new_n41270_, new_n41271_, new_n41272_, new_n41273_,
    new_n41274_, new_n41275_, new_n41276_, new_n41277_, new_n41278_,
    new_n41279_, new_n41280_, new_n41281_, new_n41282_, new_n41283_,
    new_n41284_, new_n41285_, new_n41286_, new_n41287_, new_n41288_,
    new_n41289_, new_n41290_, new_n41291_, new_n41292_, new_n41293_,
    new_n41294_, new_n41295_, new_n41296_, new_n41297_, new_n41298_,
    new_n41299_, new_n41300_, new_n41301_, new_n41302_, new_n41303_,
    new_n41304_, new_n41305_, new_n41306_, new_n41307_, new_n41308_,
    new_n41309_, new_n41310_, new_n41311_, new_n41312_, new_n41313_,
    new_n41314_, new_n41315_, new_n41316_, new_n41317_, new_n41318_,
    new_n41319_, new_n41320_, new_n41321_, new_n41322_, new_n41323_,
    new_n41324_, new_n41325_, new_n41326_, new_n41327_, new_n41328_,
    new_n41329_, new_n41330_, new_n41331_, new_n41332_, new_n41333_,
    new_n41334_, new_n41335_, new_n41336_, new_n41337_, new_n41338_,
    new_n41339_, new_n41340_, new_n41341_, new_n41342_, new_n41343_,
    new_n41344_, new_n41345_, new_n41346_, new_n41347_, new_n41348_,
    new_n41349_, new_n41350_, new_n41351_, new_n41352_, new_n41353_,
    new_n41354_, new_n41355_, new_n41356_, new_n41357_, new_n41358_,
    new_n41359_, new_n41360_, new_n41361_, new_n41362_, new_n41363_,
    new_n41364_, new_n41365_, new_n41366_, new_n41367_, new_n41368_,
    new_n41369_, new_n41370_, new_n41371_, new_n41372_, new_n41373_,
    new_n41374_, new_n41375_, new_n41376_, new_n41377_, new_n41378_,
    new_n41379_, new_n41380_, new_n41381_, new_n41382_, new_n41383_,
    new_n41384_, new_n41385_, new_n41386_, new_n41387_, new_n41388_,
    new_n41389_, new_n41390_, new_n41391_, new_n41392_, new_n41393_,
    new_n41394_, new_n41395_, new_n41396_, new_n41397_, new_n41398_,
    new_n41399_, new_n41400_, new_n41401_, new_n41402_, new_n41403_,
    new_n41404_, new_n41405_, new_n41406_, new_n41407_, new_n41408_,
    new_n41409_, new_n41410_, new_n41411_, new_n41412_, new_n41413_,
    new_n41414_, new_n41415_, new_n41416_, new_n41417_, new_n41418_,
    new_n41419_, new_n41420_, new_n41421_, new_n41422_, new_n41423_,
    new_n41424_, new_n41425_, new_n41426_, new_n41427_, new_n41428_,
    new_n41429_, new_n41430_, new_n41431_, new_n41432_, new_n41433_,
    new_n41434_, new_n41435_, new_n41436_, new_n41437_, new_n41438_,
    new_n41439_, new_n41440_, new_n41441_, new_n41442_, new_n41443_,
    new_n41444_, new_n41445_, new_n41446_, new_n41447_, new_n41448_,
    new_n41449_, new_n41450_, new_n41451_, new_n41452_, new_n41453_,
    new_n41454_, new_n41455_, new_n41456_, new_n41457_, new_n41458_,
    new_n41459_, new_n41460_, new_n41461_, new_n41462_, new_n41463_,
    new_n41464_, new_n41465_, new_n41466_, new_n41467_, new_n41468_,
    new_n41469_, new_n41470_, new_n41471_, new_n41472_, new_n41473_,
    new_n41474_, new_n41475_, new_n41476_, new_n41477_, new_n41478_,
    new_n41479_, new_n41480_, new_n41481_, new_n41482_, new_n41483_,
    new_n41484_, new_n41485_, new_n41486_, new_n41487_, new_n41488_,
    new_n41489_, new_n41490_, new_n41491_, new_n41492_, new_n41493_,
    new_n41494_, new_n41495_, new_n41496_, new_n41497_, new_n41498_,
    new_n41499_, new_n41500_, new_n41501_, new_n41502_, new_n41503_,
    new_n41504_, new_n41505_, new_n41506_, new_n41507_, new_n41508_,
    new_n41509_, new_n41510_, new_n41511_, new_n41512_, new_n41513_,
    new_n41514_, new_n41515_, new_n41516_, new_n41517_, new_n41518_,
    new_n41519_, new_n41520_, new_n41521_, new_n41522_, new_n41523_,
    new_n41524_, new_n41525_, new_n41526_, new_n41527_, new_n41528_,
    new_n41529_, new_n41530_, new_n41531_, new_n41532_, new_n41533_,
    new_n41534_, new_n41535_, new_n41536_, new_n41537_, new_n41538_,
    new_n41539_, new_n41540_, new_n41541_, new_n41542_, new_n41543_,
    new_n41544_, new_n41545_, new_n41546_, new_n41547_, new_n41548_,
    new_n41549_, new_n41550_, new_n41551_, new_n41552_, new_n41553_,
    new_n41554_, new_n41555_, new_n41556_, new_n41557_, new_n41558_,
    new_n41559_, new_n41560_, new_n41561_, new_n41562_, new_n41563_,
    new_n41564_, new_n41565_, new_n41566_, new_n41567_, new_n41568_,
    new_n41569_, new_n41570_, new_n41571_, new_n41572_, new_n41573_,
    new_n41574_, new_n41575_, new_n41576_, new_n41577_, new_n41578_,
    new_n41579_, new_n41580_, new_n41581_, new_n41582_, new_n41583_,
    new_n41584_, new_n41585_, new_n41586_, new_n41587_, new_n41588_,
    new_n41589_, new_n41590_, new_n41591_, new_n41592_, new_n41593_,
    new_n41594_, new_n41595_, new_n41596_, new_n41597_, new_n41598_,
    new_n41599_, new_n41600_, new_n41601_, new_n41602_, new_n41603_,
    new_n41604_, new_n41605_, new_n41606_, new_n41607_, new_n41608_,
    new_n41609_, new_n41610_, new_n41611_, new_n41612_, new_n41613_,
    new_n41614_, new_n41615_, new_n41616_, new_n41617_, new_n41618_,
    new_n41619_, new_n41620_, new_n41621_, new_n41622_, new_n41623_,
    new_n41624_, new_n41625_, new_n41626_, new_n41627_, new_n41628_,
    new_n41629_, new_n41630_, new_n41631_, new_n41632_, new_n41633_,
    new_n41634_, new_n41635_, new_n41636_, new_n41637_, new_n41638_,
    new_n41639_, new_n41640_, new_n41641_, new_n41642_, new_n41643_,
    new_n41644_, new_n41645_, new_n41646_, new_n41647_, new_n41648_,
    new_n41649_, new_n41650_, new_n41651_, new_n41652_, new_n41653_,
    new_n41654_, new_n41655_, new_n41656_, new_n41657_, new_n41658_,
    new_n41659_, new_n41660_, new_n41661_, new_n41662_, new_n41663_,
    new_n41664_, new_n41665_, new_n41666_, new_n41667_, new_n41668_,
    new_n41669_, new_n41670_, new_n41671_, new_n41672_, new_n41673_,
    new_n41674_, new_n41675_, new_n41676_, new_n41677_, new_n41678_,
    new_n41679_, new_n41680_, new_n41681_, new_n41682_, new_n41683_,
    new_n41684_, new_n41685_, new_n41686_, new_n41687_, new_n41688_,
    new_n41689_, new_n41690_, new_n41691_, new_n41692_, new_n41693_,
    new_n41694_, new_n41695_, new_n41696_, new_n41697_, new_n41698_,
    new_n41699_, new_n41700_, new_n41701_, new_n41702_, new_n41703_,
    new_n41704_, new_n41705_, new_n41706_, new_n41707_, new_n41708_,
    new_n41709_, new_n41710_, new_n41711_, new_n41712_, new_n41713_,
    new_n41714_, new_n41715_, new_n41716_, new_n41717_, new_n41718_,
    new_n41719_, new_n41720_, new_n41721_, new_n41722_, new_n41723_,
    new_n41724_, new_n41725_, new_n41726_, new_n41727_, new_n41728_,
    new_n41729_, new_n41730_, new_n41731_, new_n41732_, new_n41733_,
    new_n41734_, new_n41735_, new_n41736_, new_n41737_, new_n41738_,
    new_n41739_, new_n41740_, new_n41741_, new_n41742_, new_n41743_,
    new_n41744_, new_n41745_, new_n41746_, new_n41747_, new_n41748_,
    new_n41749_, new_n41750_, new_n41751_, new_n41752_, new_n41753_,
    new_n41754_, new_n41755_, new_n41756_, new_n41757_, new_n41758_,
    new_n41759_, new_n41760_, new_n41761_, new_n41762_, new_n41763_,
    new_n41764_, new_n41765_, new_n41766_, new_n41767_, new_n41768_,
    new_n41769_, new_n41770_, new_n41771_, new_n41772_, new_n41773_,
    new_n41774_, new_n41775_, new_n41776_, new_n41777_, new_n41778_,
    new_n41779_, new_n41780_, new_n41781_, new_n41782_, new_n41783_,
    new_n41784_, new_n41785_, new_n41786_, new_n41787_, new_n41788_,
    new_n41789_, new_n41790_, new_n41791_, new_n41792_, new_n41793_,
    new_n41794_, new_n41795_, new_n41796_, new_n41797_, new_n41798_,
    new_n41799_, new_n41800_, new_n41801_, new_n41802_, new_n41803_,
    new_n41804_, new_n41805_, new_n41806_, new_n41807_, new_n41808_,
    new_n41809_, new_n41810_, new_n41811_, new_n41812_, new_n41813_,
    new_n41814_, new_n41815_, new_n41816_, new_n41817_, new_n41818_,
    new_n41819_, new_n41820_, new_n41821_, new_n41822_, new_n41823_,
    new_n41824_, new_n41825_, new_n41826_, new_n41827_, new_n41828_,
    new_n41829_, new_n41830_, new_n41831_, new_n41832_, new_n41833_,
    new_n41834_, new_n41835_, new_n41836_, new_n41837_, new_n41838_,
    new_n41839_, new_n41840_, new_n41841_, new_n41842_, new_n41843_,
    new_n41844_, new_n41845_, new_n41846_, new_n41847_, new_n41848_,
    new_n41849_, new_n41850_, new_n41851_, new_n41852_, new_n41853_,
    new_n41854_, new_n41855_, new_n41856_, new_n41857_, new_n41858_,
    new_n41859_, new_n41860_, new_n41861_, new_n41862_, new_n41863_,
    new_n41864_, new_n41865_, new_n41866_, new_n41867_, new_n41868_,
    new_n41869_, new_n41870_, new_n41871_, new_n41872_, new_n41873_,
    new_n41874_, new_n41875_, new_n41876_, new_n41877_, new_n41878_,
    new_n41879_, new_n41880_, new_n41881_, new_n41882_, new_n41883_,
    new_n41884_, new_n41885_, new_n41886_, new_n41887_, new_n41888_,
    new_n41889_, new_n41890_, new_n41891_, new_n41892_, new_n41893_,
    new_n41894_, new_n41895_, new_n41896_, new_n41897_, new_n41898_,
    new_n41899_, new_n41900_, new_n41901_, new_n41902_, new_n41903_,
    new_n41904_, new_n41905_, new_n41906_, new_n41907_, new_n41908_,
    new_n41909_, new_n41910_, new_n41911_, new_n41912_, new_n41913_,
    new_n41914_, new_n41915_, new_n41916_, new_n41917_, new_n41918_,
    new_n41919_, new_n41920_, new_n41921_, new_n41922_, new_n41923_,
    new_n41924_, new_n41925_, new_n41926_, new_n41927_, new_n41928_,
    new_n41929_, new_n41930_, new_n41931_, new_n41932_, new_n41933_,
    new_n41934_, new_n41935_, new_n41936_, new_n41937_, new_n41938_,
    new_n41939_, new_n41940_, new_n41941_, new_n41942_, new_n41943_,
    new_n41944_, new_n41945_, new_n41946_, new_n41947_, new_n41948_,
    new_n41949_, new_n41950_, new_n41951_, new_n41952_, new_n41953_,
    new_n41954_, new_n41955_, new_n41956_, new_n41957_, new_n41958_,
    new_n41959_, new_n41960_, new_n41961_, new_n41962_, new_n41963_,
    new_n41964_, new_n41965_, new_n41966_, new_n41967_, new_n41968_,
    new_n41969_, new_n41970_, new_n41971_, new_n41972_, new_n41973_,
    new_n41974_, new_n41975_, new_n41976_, new_n41977_, new_n41978_,
    new_n41979_, new_n41980_, new_n41981_, new_n41982_, new_n41983_,
    new_n41984_, new_n41985_, new_n41986_, new_n41987_, new_n41988_,
    new_n41989_, new_n41990_, new_n41991_, new_n41992_, new_n41993_,
    new_n41994_, new_n41995_, new_n41996_, new_n41997_, new_n41998_,
    new_n41999_, new_n42000_, new_n42001_, new_n42002_, new_n42003_,
    new_n42004_, new_n42005_, new_n42006_, new_n42007_, new_n42008_,
    new_n42009_, new_n42010_, new_n42011_, new_n42012_, new_n42013_,
    new_n42014_, new_n42015_, new_n42016_, new_n42017_, new_n42018_,
    new_n42019_, new_n42020_, new_n42021_, new_n42022_, new_n42023_,
    new_n42024_, new_n42025_, new_n42026_, new_n42027_, new_n42028_,
    new_n42029_, new_n42030_, new_n42031_, new_n42032_, new_n42033_,
    new_n42034_, new_n42035_, new_n42036_, new_n42037_, new_n42038_,
    new_n42039_, new_n42040_, new_n42041_, new_n42042_, new_n42043_,
    new_n42044_, new_n42045_, new_n42046_, new_n42047_, new_n42048_,
    new_n42049_, new_n42050_, new_n42051_, new_n42052_, new_n42053_,
    new_n42054_, new_n42055_, new_n42056_, new_n42057_, new_n42058_,
    new_n42059_, new_n42060_, new_n42061_, new_n42062_, new_n42063_,
    new_n42064_, new_n42065_, new_n42066_, new_n42067_, new_n42068_,
    new_n42069_, new_n42070_, new_n42071_, new_n42072_, new_n42073_,
    new_n42074_, new_n42075_, new_n42076_, new_n42077_, new_n42078_,
    new_n42079_, new_n42080_, new_n42081_, new_n42082_, new_n42083_,
    new_n42084_, new_n42085_, new_n42086_, new_n42087_, new_n42088_,
    new_n42089_, new_n42090_, new_n42091_, new_n42092_, new_n42093_,
    new_n42094_, new_n42095_, new_n42096_, new_n42097_, new_n42098_,
    new_n42099_, new_n42100_, new_n42101_, new_n42102_, new_n42103_,
    new_n42104_, new_n42105_, new_n42106_, new_n42107_, new_n42108_,
    new_n42109_, new_n42110_, new_n42111_, new_n42112_, new_n42113_,
    new_n42114_, new_n42115_, new_n42116_, new_n42117_, new_n42118_,
    new_n42119_, new_n42120_, new_n42121_, new_n42122_, new_n42123_,
    new_n42124_, new_n42125_, new_n42126_, new_n42127_, new_n42128_,
    new_n42129_, new_n42130_, new_n42131_, new_n42132_, new_n42133_,
    new_n42134_, new_n42135_, new_n42136_, new_n42137_, new_n42138_,
    new_n42139_, new_n42140_, new_n42141_, new_n42142_, new_n42143_,
    new_n42144_, new_n42145_, new_n42146_, new_n42147_, new_n42148_,
    new_n42149_, new_n42150_, new_n42151_, new_n42152_, new_n42153_,
    new_n42154_, new_n42155_, new_n42156_, new_n42157_, new_n42158_,
    new_n42159_, new_n42160_, new_n42161_, new_n42162_, new_n42163_,
    new_n42164_, new_n42165_, new_n42166_, new_n42167_, new_n42168_,
    new_n42169_, new_n42170_, new_n42171_, new_n42172_, new_n42173_,
    new_n42174_, new_n42175_, new_n42176_, new_n42177_, new_n42178_,
    new_n42179_, new_n42180_, new_n42181_, new_n42182_, new_n42183_,
    new_n42184_, new_n42185_, new_n42186_, new_n42187_, new_n42188_,
    new_n42189_, new_n42190_, new_n42191_, new_n42192_, new_n42193_,
    new_n42194_, new_n42195_, new_n42196_, new_n42197_, new_n42198_,
    new_n42199_, new_n42200_, new_n42201_, new_n42202_, new_n42203_,
    new_n42204_, new_n42205_, new_n42206_, new_n42207_, new_n42208_,
    new_n42209_, new_n42210_, new_n42211_, new_n42212_, new_n42213_,
    new_n42214_, new_n42215_, new_n42216_, new_n42217_, new_n42218_,
    new_n42219_, new_n42220_, new_n42221_, new_n42222_, new_n42223_,
    new_n42224_, new_n42225_, new_n42226_, new_n42227_, new_n42228_,
    new_n42229_, new_n42230_, new_n42231_, new_n42232_, new_n42233_,
    new_n42234_, new_n42235_, new_n42236_, new_n42237_, new_n42238_,
    new_n42239_, new_n42240_, new_n42241_, new_n42242_, new_n42243_,
    new_n42244_, new_n42245_, new_n42246_, new_n42247_, new_n42248_,
    new_n42249_, new_n42250_, new_n42251_, new_n42252_, new_n42253_,
    new_n42254_, new_n42255_, new_n42256_, new_n42257_, new_n42258_,
    new_n42259_, new_n42260_, new_n42261_, new_n42262_, new_n42263_,
    new_n42264_, new_n42265_, new_n42266_, new_n42267_, new_n42268_,
    new_n42269_, new_n42270_, new_n42271_, new_n42272_, new_n42273_,
    new_n42274_, new_n42275_, new_n42276_, new_n42277_, new_n42278_,
    new_n42279_, new_n42280_, new_n42281_, new_n42282_, new_n42283_,
    new_n42284_, new_n42285_, new_n42286_, new_n42287_, new_n42288_,
    new_n42289_, new_n42290_, new_n42291_, new_n42292_, new_n42293_,
    new_n42294_, new_n42295_, new_n42296_, new_n42297_, new_n42298_,
    new_n42299_, new_n42300_, new_n42301_, new_n42302_, new_n42303_,
    new_n42304_, new_n42305_, new_n42306_, new_n42307_, new_n42308_,
    new_n42309_, new_n42310_, new_n42311_, new_n42312_, new_n42313_,
    new_n42314_, new_n42315_, new_n42316_, new_n42317_, new_n42318_,
    new_n42319_, new_n42320_, new_n42321_, new_n42322_, new_n42323_,
    new_n42324_, new_n42325_, new_n42326_, new_n42327_, new_n42328_,
    new_n42329_, new_n42330_, new_n42331_, new_n42332_, new_n42333_,
    new_n42334_, new_n42335_, new_n42336_, new_n42337_, new_n42338_,
    new_n42339_, new_n42340_, new_n42341_, new_n42342_, new_n42343_,
    new_n42344_, new_n42345_, new_n42346_, new_n42347_, new_n42348_,
    new_n42349_, new_n42350_, new_n42351_, new_n42352_, new_n42353_,
    new_n42354_, new_n42355_, new_n42356_, new_n42357_, new_n42358_,
    new_n42359_, new_n42360_, new_n42361_, new_n42362_, new_n42363_,
    new_n42364_, new_n42365_, new_n42366_, new_n42367_, new_n42368_,
    new_n42369_, new_n42370_, new_n42371_, new_n42372_, new_n42373_,
    new_n42374_, new_n42375_, new_n42376_, new_n42377_, new_n42378_,
    new_n42379_, new_n42380_, new_n42381_, new_n42382_, new_n42383_,
    new_n42384_, new_n42385_, new_n42386_, new_n42387_, new_n42388_,
    new_n42389_, new_n42390_, new_n42391_, new_n42392_, new_n42393_,
    new_n42394_, new_n42395_, new_n42396_, new_n42397_, new_n42398_,
    new_n42399_, new_n42400_, new_n42401_, new_n42402_, new_n42403_,
    new_n42404_, new_n42405_, new_n42406_, new_n42407_, new_n42408_,
    new_n42409_, new_n42410_, new_n42411_, new_n42412_, new_n42413_,
    new_n42414_, new_n42415_, new_n42416_, new_n42417_, new_n42418_,
    new_n42419_, new_n42420_, new_n42421_, new_n42422_, new_n42423_,
    new_n42424_, new_n42425_, new_n42426_, new_n42427_, new_n42428_,
    new_n42429_, new_n42430_, new_n42431_, new_n42432_, new_n42433_,
    new_n42434_, new_n42435_, new_n42436_, new_n42437_, new_n42438_,
    new_n42439_, new_n42440_, new_n42441_, new_n42442_, new_n42443_,
    new_n42444_, new_n42445_, new_n42446_, new_n42447_, new_n42448_,
    new_n42449_, new_n42450_, new_n42451_, new_n42452_, new_n42453_,
    new_n42454_, new_n42455_, new_n42456_, new_n42457_, new_n42458_,
    new_n42459_, new_n42460_, new_n42461_, new_n42462_, new_n42463_,
    new_n42464_, new_n42465_, new_n42466_, new_n42467_, new_n42468_,
    new_n42469_, new_n42470_, new_n42471_, new_n42472_, new_n42473_,
    new_n42474_, new_n42475_, new_n42476_, new_n42477_, new_n42478_,
    new_n42479_, new_n42480_, new_n42481_, new_n42482_, new_n42483_,
    new_n42484_, new_n42485_, new_n42486_, new_n42487_, new_n42488_,
    new_n42489_, new_n42490_, new_n42491_, new_n42492_, new_n42493_,
    new_n42494_, new_n42495_, new_n42496_, new_n42497_, new_n42498_,
    new_n42499_, new_n42500_, new_n42501_, new_n42502_, new_n42503_,
    new_n42504_, new_n42505_, new_n42506_, new_n42507_, new_n42508_,
    new_n42509_, new_n42510_, new_n42511_, new_n42512_, new_n42513_,
    new_n42514_, new_n42515_, new_n42516_, new_n42517_, new_n42518_,
    new_n42519_, new_n42520_, new_n42521_, new_n42522_, new_n42523_,
    new_n42524_, new_n42525_, new_n42526_, new_n42527_, new_n42528_,
    new_n42529_, new_n42530_, new_n42531_, new_n42532_, new_n42533_,
    new_n42534_, new_n42535_, new_n42536_, new_n42537_, new_n42538_,
    new_n42539_, new_n42540_, new_n42541_, new_n42542_, new_n42543_,
    new_n42544_, new_n42545_, new_n42546_, new_n42547_, new_n42548_,
    new_n42549_, new_n42550_, new_n42551_, new_n42552_, new_n42553_,
    new_n42554_, new_n42555_, new_n42556_, new_n42557_, new_n42558_,
    new_n42559_, new_n42560_, new_n42561_, new_n42562_, new_n42563_,
    new_n42564_, new_n42565_, new_n42566_, new_n42567_, new_n42568_,
    new_n42569_, new_n42570_, new_n42571_, new_n42572_, new_n42573_,
    new_n42574_, new_n42575_, new_n42576_, new_n42577_, new_n42578_,
    new_n42579_, new_n42580_, new_n42581_, new_n42582_, new_n42583_,
    new_n42584_, new_n42585_, new_n42586_, new_n42587_, new_n42588_,
    new_n42589_, new_n42590_, new_n42591_, new_n42592_, new_n42593_,
    new_n42594_, new_n42595_, new_n42596_, new_n42597_, new_n42598_,
    new_n42599_, new_n42600_, new_n42601_, new_n42602_, new_n42603_,
    new_n42604_, new_n42605_, new_n42606_, new_n42607_, new_n42608_,
    new_n42609_, new_n42610_, new_n42611_, new_n42612_, new_n42613_,
    new_n42614_, new_n42615_, new_n42616_, new_n42617_, new_n42618_,
    new_n42619_, new_n42620_, new_n42621_, new_n42622_, new_n42623_,
    new_n42624_, new_n42625_, new_n42626_, new_n42627_, new_n42628_,
    new_n42629_, new_n42630_, new_n42631_, new_n42632_, new_n42633_,
    new_n42634_, new_n42635_, new_n42636_, new_n42637_, new_n42638_,
    new_n42639_, new_n42640_, new_n42641_, new_n42642_, new_n42643_,
    new_n42644_, new_n42645_, new_n42646_, new_n42647_, new_n42648_,
    new_n42649_, new_n42650_, new_n42651_, new_n42652_, new_n42653_,
    new_n42654_, new_n42655_, new_n42656_, new_n42657_, new_n42658_,
    new_n42659_, new_n42660_, new_n42661_, new_n42662_, new_n42663_,
    new_n42664_, new_n42665_, new_n42666_, new_n42667_, new_n42668_,
    new_n42669_, new_n42670_, new_n42671_, new_n42672_, new_n42673_,
    new_n42674_, new_n42675_, new_n42676_, new_n42677_, new_n42678_,
    new_n42679_, new_n42680_, new_n42681_, new_n42682_, new_n42683_,
    new_n42684_, new_n42685_, new_n42686_, new_n42687_, new_n42688_,
    new_n42689_, new_n42690_, new_n42691_, new_n42692_, new_n42693_,
    new_n42694_, new_n42695_, new_n42696_, new_n42697_, new_n42698_,
    new_n42699_, new_n42700_, new_n42701_, new_n42702_, new_n42703_,
    new_n42704_, new_n42705_, new_n42706_, new_n42707_, new_n42708_,
    new_n42709_, new_n42710_, new_n42711_, new_n42712_, new_n42713_,
    new_n42714_, new_n42715_, new_n42716_, new_n42717_, new_n42718_,
    new_n42719_, new_n42720_, new_n42721_, new_n42722_, new_n42723_,
    new_n42724_, new_n42725_, new_n42726_, new_n42727_, new_n42728_,
    new_n42729_, new_n42730_, new_n42731_, new_n42732_, new_n42733_,
    new_n42734_, new_n42735_, new_n42736_, new_n42737_, new_n42738_,
    new_n42739_, new_n42740_, new_n42741_, new_n42742_, new_n42743_,
    new_n42744_, new_n42745_, new_n42746_, new_n42747_, new_n42748_,
    new_n42749_, new_n42750_, new_n42751_, new_n42752_, new_n42753_,
    new_n42754_, new_n42755_, new_n42756_, new_n42757_, new_n42758_,
    new_n42759_, new_n42760_, new_n42761_, new_n42762_, new_n42763_,
    new_n42764_, new_n42765_, new_n42766_, new_n42767_, new_n42768_,
    new_n42769_, new_n42770_, new_n42771_, new_n42772_, new_n42773_,
    new_n42774_, new_n42775_, new_n42776_, new_n42777_, new_n42778_,
    new_n42779_, new_n42780_, new_n42781_, new_n42782_, new_n42783_,
    new_n42784_, new_n42785_, new_n42786_, new_n42787_, new_n42788_,
    new_n42789_, new_n42790_, new_n42791_, new_n42792_, new_n42793_,
    new_n42794_, new_n42795_, new_n42796_, new_n42797_, new_n42798_,
    new_n42799_, new_n42800_, new_n42801_, new_n42802_, new_n42803_,
    new_n42804_, new_n42805_, new_n42806_, new_n42807_, new_n42808_,
    new_n42809_, new_n42810_, new_n42811_, new_n42812_, new_n42813_,
    new_n42814_, new_n42815_, new_n42816_, new_n42817_, new_n42818_,
    new_n42819_, new_n42820_, new_n42821_, new_n42822_, new_n42823_,
    new_n42824_, new_n42825_, new_n42826_, new_n42827_, new_n42828_,
    new_n42829_, new_n42830_, new_n42831_, new_n42832_, new_n42833_,
    new_n42834_, new_n42835_, new_n42836_, new_n42837_, new_n42838_,
    new_n42839_, new_n42840_, new_n42841_, new_n42842_, new_n42843_,
    new_n42844_, new_n42845_, new_n42846_, new_n42847_, new_n42848_,
    new_n42849_, new_n42850_, new_n42851_, new_n42852_, new_n42853_,
    new_n42854_, new_n42855_, new_n42856_, new_n42857_, new_n42858_,
    new_n42859_, new_n42860_, new_n42861_, new_n42862_, new_n42863_,
    new_n42864_, new_n42865_, new_n42866_, new_n42867_, new_n42868_,
    new_n42869_, new_n42870_, new_n42871_, new_n42872_, new_n42873_,
    new_n42874_, new_n42875_, new_n42876_, new_n42877_, new_n42878_,
    new_n42879_, new_n42880_, new_n42881_, new_n42882_, new_n42883_,
    new_n42884_, new_n42885_, new_n42886_, new_n42887_, new_n42888_,
    new_n42889_, new_n42890_, new_n42891_, new_n42892_, new_n42893_,
    new_n42894_, new_n42895_, new_n42896_, new_n42897_, new_n42898_,
    new_n42899_, new_n42900_, new_n42901_, new_n42902_, new_n42903_,
    new_n42904_, new_n42905_, new_n42906_, new_n42907_, new_n42908_,
    new_n42909_, new_n42910_, new_n42911_, new_n42912_, new_n42913_,
    new_n42914_, new_n42915_, new_n42916_, new_n42917_, new_n42918_,
    new_n42919_, new_n42920_, new_n42921_, new_n42922_, new_n42923_,
    new_n42924_, new_n42925_, new_n42926_, new_n42927_, new_n42928_,
    new_n42929_, new_n42930_, new_n42931_, new_n42932_, new_n42933_,
    new_n42934_, new_n42935_, new_n42936_, new_n42937_, new_n42938_,
    new_n42939_, new_n42940_, new_n42941_, new_n42942_, new_n42943_,
    new_n42944_, new_n42945_, new_n42946_, new_n42947_, new_n42948_,
    new_n42949_, new_n42950_, new_n42951_, new_n42952_, new_n42953_,
    new_n42954_, new_n42955_, new_n42956_, new_n42957_, new_n42958_,
    new_n42959_, new_n42960_, new_n42961_, new_n42962_, new_n42963_,
    new_n42964_, new_n42965_, new_n42966_, new_n42967_, new_n42968_,
    new_n42969_, new_n42970_, new_n42971_, new_n42972_, new_n42973_,
    new_n42974_, new_n42975_, new_n42976_, new_n42977_, new_n42978_,
    new_n42979_, new_n42980_, new_n42981_, new_n42982_, new_n42983_,
    new_n42984_, new_n42985_, new_n42986_, new_n42987_, new_n42988_,
    new_n42989_, new_n42990_, new_n42991_, new_n42992_, new_n42993_,
    new_n42994_, new_n42995_, new_n42996_, new_n42997_, new_n42998_,
    new_n42999_, new_n43000_, new_n43001_, new_n43002_, new_n43003_,
    new_n43004_, new_n43005_, new_n43006_, new_n43007_, new_n43008_,
    new_n43009_, new_n43010_, new_n43011_, new_n43012_, new_n43013_,
    new_n43014_, new_n43015_, new_n43016_, new_n43017_, new_n43018_,
    new_n43019_, new_n43020_, new_n43021_, new_n43022_, new_n43023_,
    new_n43024_, new_n43025_, new_n43026_, new_n43027_, new_n43028_,
    new_n43029_, new_n43030_, new_n43031_, new_n43032_, new_n43033_,
    new_n43034_, new_n43035_, new_n43036_, new_n43037_, new_n43038_,
    new_n43039_, new_n43040_, new_n43041_, new_n43042_, new_n43043_,
    new_n43044_, new_n43045_, new_n43046_, new_n43047_, new_n43048_,
    new_n43049_, new_n43050_, new_n43051_, new_n43052_, new_n43053_,
    new_n43054_, new_n43055_, new_n43056_, new_n43057_, new_n43058_,
    new_n43059_, new_n43060_, new_n43061_, new_n43062_, new_n43063_,
    new_n43064_, new_n43065_, new_n43066_, new_n43067_, new_n43068_,
    new_n43069_, new_n43070_, new_n43071_, new_n43072_, new_n43073_,
    new_n43074_, new_n43075_, new_n43076_, new_n43077_, new_n43078_,
    new_n43079_, new_n43080_, new_n43081_, new_n43082_, new_n43083_,
    new_n43084_, new_n43085_, new_n43086_, new_n43087_, new_n43088_,
    new_n43089_, new_n43090_, new_n43091_, new_n43092_, new_n43093_,
    new_n43094_, new_n43095_, new_n43096_, new_n43097_, new_n43098_,
    new_n43099_, new_n43100_, new_n43101_, new_n43102_, new_n43103_,
    new_n43104_, new_n43105_, new_n43106_, new_n43107_, new_n43108_,
    new_n43109_, new_n43110_, new_n43111_, new_n43112_, new_n43113_,
    new_n43114_, new_n43115_, new_n43116_, new_n43117_, new_n43118_,
    new_n43119_, new_n43120_, new_n43121_, new_n43122_, new_n43123_,
    new_n43124_, new_n43125_, new_n43126_, new_n43127_, new_n43128_,
    new_n43129_, new_n43130_, new_n43131_, new_n43132_, new_n43133_,
    new_n43134_, new_n43135_, new_n43136_, new_n43137_, new_n43138_,
    new_n43139_, new_n43140_, new_n43141_, new_n43142_, new_n43143_,
    new_n43144_, new_n43145_, new_n43146_, new_n43147_, new_n43148_,
    new_n43149_, new_n43150_, new_n43151_, new_n43152_, new_n43153_,
    new_n43154_, new_n43155_, new_n43156_, new_n43157_, new_n43158_,
    new_n43159_, new_n43160_, new_n43161_, new_n43162_, new_n43163_,
    new_n43164_, new_n43165_, new_n43166_, new_n43167_, new_n43168_,
    new_n43169_, new_n43170_, new_n43171_, new_n43172_, new_n43173_,
    new_n43174_, new_n43175_, new_n43176_, new_n43177_, new_n43178_,
    new_n43179_, new_n43180_, new_n43181_, new_n43182_, new_n43183_,
    new_n43184_, new_n43185_, new_n43186_, new_n43187_, new_n43188_,
    new_n43189_, new_n43190_, new_n43191_, new_n43192_, new_n43193_,
    new_n43194_, new_n43195_, new_n43196_, new_n43197_, new_n43198_,
    new_n43199_, new_n43200_, new_n43201_, new_n43202_, new_n43203_,
    new_n43204_, new_n43205_, new_n43206_, new_n43207_, new_n43208_,
    new_n43209_, new_n43210_, new_n43211_, new_n43212_, new_n43213_,
    new_n43214_, new_n43215_, new_n43216_, new_n43217_, new_n43218_,
    new_n43219_, new_n43220_, new_n43221_, new_n43222_, new_n43223_,
    new_n43224_, new_n43225_, new_n43226_, new_n43227_, new_n43228_,
    new_n43229_, new_n43230_, new_n43231_, new_n43232_, new_n43233_,
    new_n43234_, new_n43235_, new_n43236_, new_n43237_, new_n43238_,
    new_n43239_, new_n43240_, new_n43241_, new_n43242_, new_n43243_,
    new_n43244_, new_n43245_, new_n43246_, new_n43247_, new_n43248_,
    new_n43249_, new_n43250_, new_n43251_, new_n43252_, new_n43253_,
    new_n43254_, new_n43255_, new_n43256_, new_n43257_, new_n43258_,
    new_n43259_, new_n43260_, new_n43261_, new_n43262_, new_n43263_,
    new_n43264_, new_n43265_, new_n43266_, new_n43267_, new_n43268_,
    new_n43269_, new_n43270_, new_n43271_, new_n43272_, new_n43273_,
    new_n43274_, new_n43275_, new_n43276_, new_n43277_, new_n43278_,
    new_n43279_, new_n43280_, new_n43281_, new_n43282_, new_n43283_,
    new_n43284_, new_n43285_, new_n43286_, new_n43287_, new_n43288_,
    new_n43289_, new_n43290_, new_n43291_, new_n43292_, new_n43293_,
    new_n43294_, new_n43295_, new_n43296_, new_n43297_, new_n43298_,
    new_n43299_, new_n43300_, new_n43301_, new_n43302_, new_n43303_,
    new_n43304_, new_n43305_, new_n43306_, new_n43307_, new_n43308_,
    new_n43309_, new_n43310_, new_n43311_, new_n43312_, new_n43313_,
    new_n43314_, new_n43315_, new_n43316_, new_n43317_, new_n43318_,
    new_n43319_, new_n43320_, new_n43321_, new_n43322_, new_n43323_,
    new_n43324_, new_n43325_, new_n43326_, new_n43327_, new_n43328_,
    new_n43329_, new_n43330_, new_n43331_, new_n43332_, new_n43333_,
    new_n43334_, new_n43335_, new_n43336_, new_n43337_, new_n43338_,
    new_n43339_, new_n43340_, new_n43341_, new_n43342_, new_n43343_,
    new_n43344_, new_n43345_, new_n43346_, new_n43347_, new_n43348_,
    new_n43349_, new_n43350_, new_n43351_, new_n43352_, new_n43353_,
    new_n43354_, new_n43355_, new_n43356_, new_n43357_, new_n43358_,
    new_n43359_, new_n43360_, new_n43361_, new_n43362_, new_n43363_,
    new_n43364_, new_n43365_, new_n43366_, new_n43367_, new_n43368_,
    new_n43369_, new_n43370_, new_n43371_, new_n43372_, new_n43373_,
    new_n43374_, new_n43375_, new_n43376_, new_n43377_, new_n43378_,
    new_n43379_, new_n43380_, new_n43381_, new_n43382_, new_n43383_,
    new_n43384_, new_n43385_, new_n43386_, new_n43387_, new_n43388_,
    new_n43389_, new_n43390_, new_n43391_, new_n43392_, new_n43393_,
    new_n43394_, new_n43395_, new_n43396_, new_n43397_, new_n43398_,
    new_n43399_, new_n43400_, new_n43401_, new_n43402_, new_n43403_,
    new_n43404_, new_n43405_, new_n43406_, new_n43407_, new_n43408_,
    new_n43409_, new_n43410_, new_n43411_, new_n43412_, new_n43413_,
    new_n43414_, new_n43415_, new_n43416_, new_n43417_, new_n43418_,
    new_n43419_, new_n43420_, new_n43421_, new_n43422_, new_n43423_,
    new_n43424_, new_n43425_, new_n43426_, new_n43427_, new_n43428_,
    new_n43429_, new_n43430_, new_n43431_, new_n43432_, new_n43433_,
    new_n43434_, new_n43435_, new_n43436_, new_n43437_, new_n43438_,
    new_n43439_, new_n43440_, new_n43441_, new_n43442_, new_n43443_,
    new_n43444_, new_n43445_, new_n43446_, new_n43447_, new_n43448_,
    new_n43449_, new_n43450_, new_n43451_, new_n43452_, new_n43453_,
    new_n43454_, new_n43455_, new_n43456_, new_n43457_, new_n43458_,
    new_n43459_, new_n43460_, new_n43461_, new_n43462_, new_n43463_,
    new_n43464_, new_n43465_, new_n43466_, new_n43467_, new_n43468_,
    new_n43469_, new_n43470_, new_n43471_, new_n43472_, new_n43473_,
    new_n43474_, new_n43475_, new_n43476_, new_n43477_, new_n43478_,
    new_n43479_, new_n43480_, new_n43481_, new_n43482_, new_n43483_,
    new_n43484_, new_n43485_, new_n43486_, new_n43487_, new_n43488_,
    new_n43489_, new_n43490_, new_n43491_, new_n43492_, new_n43493_,
    new_n43494_, new_n43495_, new_n43496_, new_n43497_, new_n43498_,
    new_n43499_, new_n43500_, new_n43501_, new_n43502_, new_n43503_,
    new_n43504_, new_n43505_, new_n43506_, new_n43507_, new_n43508_,
    new_n43509_, new_n43510_, new_n43511_, new_n43512_, new_n43513_,
    new_n43514_, new_n43515_, new_n43516_, new_n43517_, new_n43518_,
    new_n43519_, new_n43520_, new_n43521_, new_n43522_, new_n43523_,
    new_n43524_, new_n43525_, new_n43526_, new_n43527_, new_n43528_,
    new_n43529_, new_n43530_, new_n43531_, new_n43532_, new_n43533_,
    new_n43534_, new_n43535_, new_n43536_, new_n43537_, new_n43538_,
    new_n43539_, new_n43540_, new_n43541_, new_n43542_, new_n43543_,
    new_n43544_, new_n43545_, new_n43546_, new_n43547_, new_n43548_,
    new_n43549_, new_n43550_, new_n43551_, new_n43552_, new_n43553_,
    new_n43554_, new_n43555_, new_n43556_, new_n43557_, new_n43558_,
    new_n43559_, new_n43560_, new_n43561_, new_n43562_, new_n43563_,
    new_n43564_, new_n43565_, new_n43566_, new_n43567_, new_n43568_,
    new_n43569_, new_n43570_, new_n43571_, new_n43572_, new_n43573_,
    new_n43574_, new_n43575_, new_n43576_, new_n43577_, new_n43578_,
    new_n43579_, new_n43580_, new_n43581_, new_n43582_, new_n43583_,
    new_n43584_, new_n43585_, new_n43586_, new_n43587_, new_n43588_,
    new_n43589_, new_n43590_, new_n43591_, new_n43592_, new_n43593_,
    new_n43594_, new_n43595_, new_n43596_, new_n43597_, new_n43598_,
    new_n43599_, new_n43600_, new_n43601_, new_n43602_, new_n43603_,
    new_n43604_, new_n43605_, new_n43606_, new_n43607_, new_n43608_,
    new_n43609_, new_n43610_, new_n43611_, new_n43612_, new_n43613_,
    new_n43614_, new_n43615_, new_n43616_, new_n43617_, new_n43618_,
    new_n43619_, new_n43620_, new_n43621_, new_n43622_, new_n43623_,
    new_n43624_, new_n43625_, new_n43626_, new_n43627_, new_n43628_,
    new_n43629_, new_n43630_, new_n43631_, new_n43632_, new_n43633_,
    new_n43634_, new_n43635_, new_n43636_, new_n43637_, new_n43638_,
    new_n43639_, new_n43640_, new_n43641_, new_n43642_, new_n43643_,
    new_n43644_, new_n43645_, new_n43646_, new_n43647_, new_n43648_,
    new_n43649_, new_n43650_, new_n43651_, new_n43652_, new_n43653_,
    new_n43654_, new_n43655_, new_n43656_, new_n43657_, new_n43658_,
    new_n43659_, new_n43660_, new_n43661_, new_n43662_, new_n43663_,
    new_n43664_, new_n43665_, new_n43666_, new_n43667_, new_n43668_,
    new_n43669_, new_n43670_, new_n43671_, new_n43672_, new_n43673_,
    new_n43674_, new_n43675_, new_n43676_, new_n43677_, new_n43678_,
    new_n43679_, new_n43680_, new_n43681_, new_n43682_, new_n43683_,
    new_n43684_, new_n43685_, new_n43686_, new_n43687_, new_n43688_,
    new_n43689_, new_n43690_, new_n43691_, new_n43692_, new_n43693_,
    new_n43694_, new_n43695_, new_n43696_, new_n43697_, new_n43698_,
    new_n43699_, new_n43700_, new_n43701_, new_n43702_, new_n43703_,
    new_n43704_, new_n43705_, new_n43706_, new_n43707_, new_n43708_,
    new_n43709_, new_n43710_, new_n43711_, new_n43712_, new_n43713_,
    new_n43714_, new_n43715_, new_n43716_, new_n43717_, new_n43718_,
    new_n43719_, new_n43720_, new_n43721_, new_n43722_, new_n43723_,
    new_n43724_, new_n43725_, new_n43726_, new_n43727_, new_n43728_,
    new_n43729_, new_n43730_, new_n43731_, new_n43732_, new_n43733_,
    new_n43734_, new_n43735_, new_n43736_, new_n43737_, new_n43738_,
    new_n43739_, new_n43740_, new_n43741_, new_n43742_, new_n43743_,
    new_n43744_, new_n43745_, new_n43746_, new_n43747_, new_n43748_,
    new_n43749_, new_n43750_, new_n43751_, new_n43752_, new_n43753_,
    new_n43754_, new_n43755_, new_n43756_, new_n43757_, new_n43758_,
    new_n43759_, new_n43760_, new_n43761_, new_n43762_, new_n43763_,
    new_n43764_, new_n43765_, new_n43766_, new_n43767_, new_n43768_,
    new_n43769_, new_n43770_, new_n43771_, new_n43772_, new_n43773_,
    new_n43774_, new_n43775_, new_n43776_, new_n43777_, new_n43778_,
    new_n43779_, new_n43780_, new_n43781_, new_n43782_, new_n43783_,
    new_n43784_, new_n43785_, new_n43786_, new_n43787_, new_n43788_,
    new_n43789_, new_n43790_, new_n43791_, new_n43792_, new_n43793_,
    new_n43794_, new_n43795_, new_n43796_, new_n43797_, new_n43798_,
    new_n43799_, new_n43800_, new_n43801_, new_n43802_, new_n43803_,
    new_n43804_, new_n43805_, new_n43806_, new_n43807_, new_n43808_,
    new_n43809_, new_n43810_, new_n43811_, new_n43812_, new_n43813_,
    new_n43814_, new_n43815_, new_n43816_, new_n43817_, new_n43818_,
    new_n43819_, new_n43820_, new_n43821_, new_n43822_, new_n43823_,
    new_n43824_, new_n43825_, new_n43826_, new_n43827_, new_n43828_,
    new_n43829_, new_n43830_, new_n43831_, new_n43832_, new_n43833_,
    new_n43834_, new_n43835_, new_n43836_, new_n43837_, new_n43838_,
    new_n43839_, new_n43840_, new_n43841_, new_n43842_, new_n43843_,
    new_n43844_, new_n43845_, new_n43846_, new_n43847_, new_n43848_,
    new_n43849_, new_n43850_, new_n43851_, new_n43852_, new_n43853_,
    new_n43854_, new_n43855_, new_n43856_, new_n43857_, new_n43858_,
    new_n43859_, new_n43860_, new_n43861_, new_n43862_, new_n43863_,
    new_n43864_, new_n43865_, new_n43866_, new_n43867_, new_n43868_,
    new_n43869_, new_n43870_, new_n43871_, new_n43872_, new_n43873_,
    new_n43874_, new_n43875_, new_n43876_, new_n43877_, new_n43878_,
    new_n43879_, new_n43880_, new_n43881_, new_n43882_, new_n43883_,
    new_n43884_, new_n43885_, new_n43886_, new_n43887_, new_n43888_,
    new_n43889_, new_n43890_, new_n43891_, new_n43892_, new_n43893_,
    new_n43894_, new_n43895_, new_n43896_, new_n43897_, new_n43898_,
    new_n43899_, new_n43900_, new_n43901_, new_n43902_, new_n43903_,
    new_n43904_, new_n43905_, new_n43906_, new_n43907_, new_n43908_,
    new_n43909_, new_n43910_, new_n43911_, new_n43912_, new_n43913_,
    new_n43914_, new_n43915_, new_n43916_, new_n43917_, new_n43918_,
    new_n43919_, new_n43920_, new_n43921_, new_n43922_, new_n43923_,
    new_n43924_, new_n43925_, new_n43926_, new_n43927_, new_n43928_,
    new_n43929_, new_n43930_, new_n43931_, new_n43932_, new_n43933_,
    new_n43934_, new_n43935_, new_n43936_, new_n43937_, new_n43938_,
    new_n43939_, new_n43940_, new_n43941_, new_n43942_, new_n43943_,
    new_n43944_, new_n43945_, new_n43946_, new_n43947_, new_n43948_,
    new_n43949_, new_n43950_, new_n43951_, new_n43952_, new_n43953_,
    new_n43954_, new_n43955_, new_n43956_, new_n43957_, new_n43958_,
    new_n43959_, new_n43960_, new_n43961_, new_n43962_, new_n43963_,
    new_n43964_, new_n43965_, new_n43966_, new_n43967_, new_n43968_,
    new_n43969_, new_n43970_, new_n43971_, new_n43972_, new_n43973_,
    new_n43974_, new_n43975_, new_n43976_, new_n43977_, new_n43978_,
    new_n43979_, new_n43980_, new_n43981_, new_n43982_, new_n43983_,
    new_n43984_, new_n43985_, new_n43986_, new_n43987_, new_n43988_,
    new_n43989_, new_n43990_, new_n43991_, new_n43992_, new_n43993_,
    new_n43994_, new_n43995_, new_n43996_, new_n43997_, new_n43998_,
    new_n43999_, new_n44000_, new_n44001_, new_n44002_, new_n44003_,
    new_n44004_, new_n44005_, new_n44006_, new_n44007_, new_n44008_,
    new_n44009_, new_n44010_, new_n44011_, new_n44012_, new_n44013_,
    new_n44014_, new_n44015_, new_n44016_, new_n44017_, new_n44018_,
    new_n44019_, new_n44020_, new_n44021_, new_n44022_, new_n44023_,
    new_n44024_, new_n44025_, new_n44026_, new_n44027_, new_n44028_,
    new_n44029_, new_n44030_, new_n44031_, new_n44032_, new_n44033_,
    new_n44034_, new_n44035_, new_n44036_, new_n44037_, new_n44038_,
    new_n44039_, new_n44040_, new_n44041_, new_n44042_, new_n44043_,
    new_n44044_, new_n44045_, new_n44046_, new_n44047_, new_n44048_,
    new_n44049_, new_n44050_, new_n44051_, new_n44052_, new_n44053_,
    new_n44054_, new_n44055_, new_n44056_, new_n44057_, new_n44058_,
    new_n44059_, new_n44060_, new_n44061_, new_n44062_, new_n44063_,
    new_n44064_, new_n44065_, new_n44066_, new_n44067_, new_n44068_,
    new_n44069_, new_n44070_, new_n44071_, new_n44072_, new_n44073_,
    new_n44074_, new_n44075_, new_n44076_, new_n44077_, new_n44078_,
    new_n44079_, new_n44080_, new_n44081_, new_n44082_, new_n44083_,
    new_n44084_, new_n44085_, new_n44086_, new_n44087_, new_n44088_,
    new_n44089_, new_n44090_, new_n44091_, new_n44092_, new_n44093_,
    new_n44094_, new_n44095_, new_n44096_, new_n44097_, new_n44098_,
    new_n44099_, new_n44100_, new_n44101_, new_n44102_, new_n44103_,
    new_n44104_, new_n44105_, new_n44106_, new_n44107_, new_n44108_,
    new_n44109_, new_n44110_, new_n44111_, new_n44112_, new_n44113_,
    new_n44114_, new_n44115_, new_n44116_, new_n44117_, new_n44118_,
    new_n44119_, new_n44120_, new_n44121_, new_n44122_, new_n44123_,
    new_n44124_, new_n44125_, new_n44126_, new_n44127_, new_n44128_,
    new_n44129_, new_n44130_, new_n44131_, new_n44132_, new_n44133_,
    new_n44134_, new_n44135_, new_n44136_, new_n44137_, new_n44138_,
    new_n44139_, new_n44140_, new_n44141_, new_n44142_, new_n44143_,
    new_n44144_, new_n44145_, new_n44146_, new_n44147_, new_n44148_,
    new_n44149_, new_n44150_, new_n44151_, new_n44152_, new_n44153_,
    new_n44154_, new_n44155_, new_n44156_, new_n44157_, new_n44158_,
    new_n44159_, new_n44160_, new_n44161_, new_n44162_, new_n44163_,
    new_n44164_, new_n44165_, new_n44166_, new_n44167_, new_n44168_,
    new_n44169_, new_n44170_, new_n44171_, new_n44172_, new_n44173_,
    new_n44174_, new_n44175_, new_n44176_, new_n44177_, new_n44178_,
    new_n44179_, new_n44180_, new_n44181_, new_n44182_, new_n44183_,
    new_n44184_, new_n44185_, new_n44186_, new_n44187_, new_n44188_,
    new_n44189_, new_n44190_, new_n44191_, new_n44192_, new_n44193_,
    new_n44194_, new_n44195_, new_n44196_, new_n44197_, new_n44198_,
    new_n44199_, new_n44200_, new_n44201_, new_n44202_, new_n44203_,
    new_n44204_, new_n44205_, new_n44206_, new_n44207_, new_n44208_,
    new_n44209_, new_n44210_, new_n44211_, new_n44212_, new_n44213_,
    new_n44214_, new_n44215_, new_n44216_, new_n44217_, new_n44218_,
    new_n44219_, new_n44220_, new_n44221_, new_n44222_, new_n44223_,
    new_n44224_, new_n44225_, new_n44226_, new_n44227_, new_n44228_,
    new_n44229_, new_n44230_, new_n44231_, new_n44232_, new_n44233_,
    new_n44234_, new_n44235_, new_n44236_, new_n44237_, new_n44238_,
    new_n44239_, new_n44240_, new_n44241_, new_n44242_, new_n44243_,
    new_n44244_, new_n44245_, new_n44246_, new_n44247_, new_n44248_,
    new_n44249_, new_n44250_, new_n44251_, new_n44252_, new_n44253_,
    new_n44254_, new_n44255_, new_n44256_, new_n44257_, new_n44258_,
    new_n44259_, new_n44260_, new_n44261_, new_n44262_, new_n44263_,
    new_n44264_, new_n44265_, new_n44266_, new_n44267_, new_n44268_,
    new_n44269_, new_n44270_, new_n44271_, new_n44272_, new_n44273_,
    new_n44274_, new_n44275_, new_n44276_, new_n44277_, new_n44278_,
    new_n44279_, new_n44280_, new_n44281_, new_n44282_, new_n44283_,
    new_n44284_, new_n44285_, new_n44286_, new_n44287_, new_n44288_,
    new_n44289_, new_n44290_, new_n44291_, new_n44292_, new_n44293_,
    new_n44294_, new_n44295_, new_n44296_, new_n44297_, new_n44298_,
    new_n44299_, new_n44300_, new_n44301_, new_n44302_, new_n44303_,
    new_n44304_, new_n44305_, new_n44306_, new_n44307_, new_n44308_,
    new_n44309_, new_n44310_, new_n44311_, new_n44312_, new_n44313_,
    new_n44314_, new_n44315_, new_n44316_, new_n44317_, new_n44318_,
    new_n44319_, new_n44320_, new_n44321_, new_n44322_, new_n44323_,
    new_n44324_, new_n44325_, new_n44326_, new_n44327_, new_n44328_,
    new_n44329_, new_n44330_, new_n44331_, new_n44332_, new_n44333_,
    new_n44334_, new_n44335_, new_n44336_, new_n44337_, new_n44338_,
    new_n44339_, new_n44340_, new_n44341_, new_n44342_, new_n44343_,
    new_n44344_, new_n44345_, new_n44346_, new_n44347_, new_n44348_,
    new_n44349_, new_n44350_, new_n44351_, new_n44352_, new_n44353_,
    new_n44354_, new_n44355_, new_n44356_, new_n44357_, new_n44358_,
    new_n44359_, new_n44360_, new_n44361_, new_n44362_, new_n44363_,
    new_n44364_, new_n44365_, new_n44366_, new_n44367_, new_n44368_,
    new_n44369_, new_n44370_, new_n44371_, new_n44372_, new_n44373_,
    new_n44374_, new_n44375_, new_n44376_, new_n44377_, new_n44378_,
    new_n44379_, new_n44380_, new_n44381_, new_n44382_, new_n44383_,
    new_n44384_, new_n44385_, new_n44386_, new_n44387_, new_n44388_,
    new_n44389_, new_n44390_, new_n44391_, new_n44392_, new_n44393_,
    new_n44394_, new_n44395_, new_n44396_, new_n44397_, new_n44398_,
    new_n44399_, new_n44400_, new_n44401_, new_n44402_, new_n44403_,
    new_n44404_, new_n44405_, new_n44406_, new_n44407_, new_n44408_,
    new_n44409_, new_n44410_, new_n44411_, new_n44412_, new_n44413_,
    new_n44414_, new_n44415_, new_n44416_, new_n44417_, new_n44418_,
    new_n44419_, new_n44420_, new_n44421_, new_n44422_, new_n44423_,
    new_n44424_, new_n44425_, new_n44426_, new_n44427_, new_n44428_,
    new_n44429_, new_n44430_, new_n44431_, new_n44432_, new_n44433_,
    new_n44434_, new_n44435_, new_n44436_, new_n44437_, new_n44438_,
    new_n44439_, new_n44440_, new_n44441_, new_n44442_, new_n44443_,
    new_n44444_, new_n44445_, new_n44446_, new_n44447_, new_n44448_,
    new_n44449_, new_n44450_, new_n44451_, new_n44452_, new_n44453_,
    new_n44454_, new_n44455_, new_n44456_, new_n44457_, new_n44458_,
    new_n44459_, new_n44460_, new_n44461_, new_n44462_, new_n44463_,
    new_n44464_, new_n44465_, new_n44466_, new_n44467_, new_n44468_,
    new_n44469_, new_n44470_, new_n44471_, new_n44472_, new_n44473_,
    new_n44474_, new_n44475_, new_n44476_, new_n44477_, new_n44478_,
    new_n44479_, new_n44480_, new_n44481_, new_n44482_, new_n44483_,
    new_n44484_, new_n44485_, new_n44486_, new_n44487_, new_n44488_,
    new_n44489_, new_n44490_, new_n44491_, new_n44492_, new_n44493_,
    new_n44494_, new_n44495_, new_n44496_, new_n44497_, new_n44498_,
    new_n44499_, new_n44500_, new_n44501_, new_n44502_, new_n44503_,
    new_n44504_, new_n44505_, new_n44506_, new_n44507_, new_n44508_,
    new_n44509_, new_n44510_, new_n44511_, new_n44512_, new_n44513_,
    new_n44514_, new_n44515_, new_n44516_, new_n44517_, new_n44518_,
    new_n44519_, new_n44520_, new_n44521_, new_n44522_, new_n44523_,
    new_n44524_, new_n44525_, new_n44526_, new_n44527_, new_n44528_,
    new_n44529_, new_n44530_, new_n44531_, new_n44532_, new_n44533_,
    new_n44534_, new_n44535_, new_n44536_, new_n44537_, new_n44538_,
    new_n44539_, new_n44540_, new_n44541_, new_n44542_, new_n44543_,
    new_n44544_, new_n44545_, new_n44546_, new_n44547_, new_n44548_,
    new_n44549_, new_n44550_, new_n44551_, new_n44552_, new_n44553_,
    new_n44554_, new_n44555_, new_n44556_, new_n44557_, new_n44558_,
    new_n44559_, new_n44560_, new_n44561_, new_n44562_, new_n44563_,
    new_n44564_, new_n44565_, new_n44566_, new_n44567_, new_n44568_,
    new_n44569_, new_n44570_, new_n44571_, new_n44572_, new_n44573_,
    new_n44574_, new_n44575_, new_n44576_, new_n44577_, new_n44578_,
    new_n44579_, new_n44580_, new_n44581_, new_n44582_, new_n44583_,
    new_n44584_, new_n44585_, new_n44586_, new_n44587_, new_n44588_,
    new_n44589_, new_n44590_, new_n44591_, new_n44592_, new_n44593_,
    new_n44594_, new_n44595_, new_n44596_, new_n44597_, new_n44598_,
    new_n44599_, new_n44600_, new_n44601_, new_n44602_, new_n44603_,
    new_n44604_, new_n44605_, new_n44606_, new_n44607_, new_n44608_,
    new_n44609_, new_n44610_, new_n44611_, new_n44612_, new_n44613_,
    new_n44614_, new_n44615_, new_n44616_, new_n44617_, new_n44618_,
    new_n44619_, new_n44620_, new_n44621_, new_n44622_, new_n44623_,
    new_n44624_, new_n44625_, new_n44626_, new_n44627_, new_n44628_,
    new_n44629_, new_n44630_, new_n44631_, new_n44632_, new_n44633_,
    new_n44634_, new_n44635_, new_n44636_, new_n44637_, new_n44638_,
    new_n44639_, new_n44640_, new_n44641_, new_n44642_, new_n44643_,
    new_n44644_, new_n44645_, new_n44646_, new_n44647_, new_n44648_,
    new_n44649_, new_n44650_, new_n44651_, new_n44652_, new_n44653_,
    new_n44654_, new_n44655_, new_n44656_, new_n44657_, new_n44658_,
    new_n44659_, new_n44660_, new_n44661_, new_n44662_, new_n44663_,
    new_n44664_, new_n44665_, new_n44666_, new_n44667_, new_n44668_,
    new_n44669_, new_n44670_, new_n44671_, new_n44672_, new_n44673_,
    new_n44674_, new_n44675_, new_n44676_, new_n44677_, new_n44678_,
    new_n44679_, new_n44680_, new_n44681_, new_n44682_, new_n44683_,
    new_n44684_, new_n44685_, new_n44686_, new_n44687_, new_n44688_,
    new_n44689_, new_n44690_, new_n44691_, new_n44692_, new_n44693_,
    new_n44694_, new_n44695_, new_n44696_, new_n44697_, new_n44698_,
    new_n44699_, new_n44700_, new_n44701_, new_n44702_, new_n44703_,
    new_n44704_, new_n44705_, new_n44706_, new_n44707_, new_n44708_,
    new_n44709_, new_n44710_, new_n44711_, new_n44712_, new_n44713_,
    new_n44714_, new_n44715_, new_n44716_, new_n44717_, new_n44718_,
    new_n44719_, new_n44720_, new_n44721_, new_n44722_, new_n44723_,
    new_n44724_, new_n44725_, new_n44726_, new_n44727_, new_n44728_,
    new_n44729_, new_n44730_, new_n44731_, new_n44732_, new_n44733_,
    new_n44734_, new_n44735_, new_n44736_, new_n44737_, new_n44738_,
    new_n44739_, new_n44740_, new_n44741_, new_n44742_, new_n44743_,
    new_n44744_, new_n44745_, new_n44746_, new_n44747_, new_n44748_,
    new_n44749_, new_n44750_, new_n44751_, new_n44752_, new_n44753_,
    new_n44754_, new_n44755_, new_n44756_, new_n44757_, new_n44758_,
    new_n44759_, new_n44760_, new_n44761_, new_n44762_, new_n44763_,
    new_n44764_, new_n44765_, new_n44766_, new_n44767_, new_n44768_,
    new_n44769_, new_n44770_, new_n44771_, new_n44772_, new_n44773_,
    new_n44774_, new_n44775_, new_n44776_, new_n44777_, new_n44778_,
    new_n44779_, new_n44780_, new_n44781_, new_n44782_, new_n44783_,
    new_n44784_, new_n44785_, new_n44786_, new_n44787_, new_n44788_,
    new_n44789_, new_n44790_, new_n44791_, new_n44792_, new_n44793_,
    new_n44794_, new_n44795_, new_n44796_, new_n44797_, new_n44798_,
    new_n44799_, new_n44800_, new_n44801_, new_n44802_, new_n44803_,
    new_n44804_, new_n44805_, new_n44806_, new_n44807_, new_n44808_,
    new_n44809_, new_n44810_, new_n44811_, new_n44812_, new_n44813_,
    new_n44814_, new_n44815_, new_n44816_, new_n44817_, new_n44818_,
    new_n44819_, new_n44820_, new_n44821_, new_n44822_, new_n44823_,
    new_n44824_, new_n44825_, new_n44826_, new_n44827_, new_n44828_,
    new_n44829_, new_n44830_, new_n44831_, new_n44832_, new_n44833_,
    new_n44834_, new_n44835_, new_n44836_, new_n44837_, new_n44838_,
    new_n44839_, new_n44840_, new_n44841_, new_n44842_, new_n44843_,
    new_n44844_, new_n44845_, new_n44846_, new_n44847_, new_n44848_,
    new_n44849_, new_n44850_, new_n44851_, new_n44852_, new_n44853_,
    new_n44854_, new_n44855_, new_n44856_, new_n44857_, new_n44858_,
    new_n44859_, new_n44860_, new_n44861_, new_n44862_, new_n44863_,
    new_n44864_, new_n44865_, new_n44866_, new_n44867_, new_n44868_,
    new_n44869_, new_n44870_, new_n44871_, new_n44872_, new_n44873_,
    new_n44874_, new_n44875_, new_n44876_, new_n44877_, new_n44878_,
    new_n44879_, new_n44880_, new_n44881_, new_n44882_, new_n44883_,
    new_n44884_, new_n44885_, new_n44886_, new_n44887_, new_n44888_,
    new_n44889_, new_n44890_, new_n44891_, new_n44892_, new_n44893_,
    new_n44894_, new_n44895_, new_n44896_, new_n44897_, new_n44898_,
    new_n44899_, new_n44900_, new_n44901_, new_n44902_, new_n44903_,
    new_n44904_, new_n44905_, new_n44906_, new_n44907_, new_n44908_,
    new_n44909_, new_n44910_, new_n44911_, new_n44912_, new_n44913_,
    new_n44914_, new_n44915_, new_n44916_, new_n44917_, new_n44918_,
    new_n44919_, new_n44920_, new_n44921_, new_n44922_, new_n44923_,
    new_n44924_, new_n44925_, new_n44926_, new_n44927_, new_n44928_,
    new_n44929_, new_n44930_, new_n44931_, new_n44932_, new_n44933_,
    new_n44934_, new_n44935_, new_n44936_, new_n44937_, new_n44938_,
    new_n44939_, new_n44940_, new_n44941_, new_n44942_, new_n44943_,
    new_n44944_, new_n44945_, new_n44946_, new_n44947_, new_n44948_,
    new_n44949_, new_n44950_, new_n44951_, new_n44952_, new_n44953_,
    new_n44954_, new_n44955_, new_n44956_, new_n44957_, new_n44958_,
    new_n44959_, new_n44960_, new_n44961_, new_n44962_, new_n44963_,
    new_n44964_, new_n44965_, new_n44966_, new_n44967_, new_n44968_,
    new_n44969_, new_n44970_, new_n44971_, new_n44972_, new_n44973_,
    new_n44974_, new_n44975_, new_n44976_, new_n44977_, new_n44978_,
    new_n44979_, new_n44980_, new_n44981_, new_n44982_, new_n44983_,
    new_n44984_, new_n44985_, new_n44986_, new_n44987_, new_n44988_,
    new_n44989_, new_n44990_, new_n44991_, new_n44992_, new_n44993_,
    new_n44994_, new_n44995_, new_n44996_, new_n44997_, new_n44998_,
    new_n44999_, new_n45000_, new_n45001_, new_n45002_, new_n45003_,
    new_n45004_, new_n45005_, new_n45006_, new_n45007_, new_n45008_,
    new_n45009_, new_n45010_, new_n45011_, new_n45012_, new_n45013_,
    new_n45014_, new_n45015_, new_n45016_, new_n45017_, new_n45018_,
    new_n45019_, new_n45020_, new_n45021_, new_n45022_, new_n45023_,
    new_n45024_, new_n45025_, new_n45026_, new_n45027_, new_n45028_,
    new_n45029_, new_n45030_, new_n45031_, new_n45032_, new_n45033_,
    new_n45034_, new_n45035_, new_n45036_, new_n45037_, new_n45038_,
    new_n45039_, new_n45040_, new_n45041_, new_n45042_, new_n45043_,
    new_n45044_, new_n45045_, new_n45046_, new_n45047_, new_n45048_,
    new_n45049_, new_n45050_, new_n45051_, new_n45052_, new_n45053_,
    new_n45054_, new_n45055_, new_n45056_, new_n45057_, new_n45058_,
    new_n45059_, new_n45060_, new_n45061_, new_n45062_, new_n45063_,
    new_n45064_, new_n45065_, new_n45066_, new_n45067_, new_n45068_,
    new_n45069_, new_n45070_, new_n45071_, new_n45072_, new_n45073_,
    new_n45074_, new_n45075_, new_n45076_, new_n45077_, new_n45078_,
    new_n45079_, new_n45080_, new_n45081_, new_n45082_, new_n45083_,
    new_n45084_, new_n45085_, new_n45086_, new_n45087_, new_n45088_,
    new_n45089_, new_n45090_, new_n45091_, new_n45092_, new_n45093_,
    new_n45094_, new_n45095_, new_n45096_, new_n45097_, new_n45098_,
    new_n45099_, new_n45100_, new_n45101_, new_n45102_, new_n45103_,
    new_n45104_, new_n45105_, new_n45106_, new_n45107_, new_n45108_,
    new_n45109_, new_n45110_, new_n45111_, new_n45112_, new_n45113_,
    new_n45114_, new_n45115_, new_n45116_, new_n45117_, new_n45118_,
    new_n45119_, new_n45120_, new_n45121_, new_n45122_, new_n45123_,
    new_n45124_, new_n45125_, new_n45126_, new_n45127_, new_n45128_,
    new_n45129_, new_n45130_, new_n45131_, new_n45132_, new_n45133_,
    new_n45134_, new_n45135_, new_n45136_, new_n45137_, new_n45138_,
    new_n45139_, new_n45140_, new_n45141_, new_n45142_, new_n45143_,
    new_n45144_, new_n45145_, new_n45146_, new_n45147_, new_n45148_,
    new_n45149_, new_n45150_, new_n45151_, new_n45152_, new_n45153_,
    new_n45154_, new_n45155_, new_n45156_, new_n45157_, new_n45158_,
    new_n45159_, new_n45160_, new_n45161_, new_n45162_, new_n45163_,
    new_n45164_, new_n45165_, new_n45166_, new_n45167_, new_n45168_,
    new_n45169_, new_n45170_, new_n45171_, new_n45172_, new_n45173_,
    new_n45174_, new_n45175_, new_n45176_, new_n45177_, new_n45178_,
    new_n45179_, new_n45180_, new_n45181_, new_n45182_, new_n45183_,
    new_n45184_, new_n45185_, new_n45186_, new_n45187_, new_n45188_,
    new_n45189_, new_n45190_, new_n45191_, new_n45192_, new_n45193_,
    new_n45194_, new_n45195_, new_n45196_, new_n45197_, new_n45198_,
    new_n45199_, new_n45200_, new_n45201_, new_n45202_, new_n45203_,
    new_n45204_, new_n45205_, new_n45206_, new_n45207_, new_n45208_,
    new_n45209_, new_n45210_, new_n45211_, new_n45212_, new_n45213_,
    new_n45214_, new_n45215_, new_n45216_, new_n45217_, new_n45218_,
    new_n45219_, new_n45220_, new_n45221_, new_n45222_, new_n45223_,
    new_n45224_, new_n45225_, new_n45226_, new_n45227_, new_n45228_,
    new_n45229_, new_n45230_, new_n45231_, new_n45232_, new_n45233_,
    new_n45234_, new_n45235_, new_n45236_, new_n45237_, new_n45238_,
    new_n45239_, new_n45240_, new_n45241_, new_n45242_, new_n45243_,
    new_n45244_, new_n45245_, new_n45246_, new_n45247_, new_n45248_,
    new_n45249_, new_n45250_, new_n45251_, new_n45252_, new_n45253_,
    new_n45254_, new_n45255_, new_n45256_, new_n45257_, new_n45258_,
    new_n45259_, new_n45260_, new_n45261_, new_n45262_, new_n45263_,
    new_n45264_, new_n45265_, new_n45266_, new_n45267_, new_n45268_,
    new_n45269_, new_n45270_, new_n45271_, new_n45272_, new_n45273_,
    new_n45274_, new_n45275_, new_n45276_, new_n45277_, new_n45278_,
    new_n45279_, new_n45280_, new_n45281_, new_n45282_, new_n45283_,
    new_n45284_, new_n45285_, new_n45286_, new_n45287_, new_n45288_,
    new_n45289_, new_n45290_, new_n45291_, new_n45292_, new_n45293_,
    new_n45294_, new_n45295_, new_n45296_, new_n45297_, new_n45298_,
    new_n45299_, new_n45300_, new_n45301_, new_n45302_, new_n45303_,
    new_n45304_, new_n45305_, new_n45306_, new_n45307_, new_n45308_,
    new_n45309_, new_n45310_, new_n45311_, new_n45312_, new_n45313_,
    new_n45314_, new_n45315_, new_n45316_, new_n45317_, new_n45318_,
    new_n45319_, new_n45320_, new_n45321_, new_n45322_, new_n45323_,
    new_n45324_, new_n45325_, new_n45326_, new_n45327_, new_n45328_,
    new_n45329_, new_n45330_, new_n45331_, new_n45332_, new_n45333_,
    new_n45334_, new_n45335_, new_n45336_, new_n45337_, new_n45338_,
    new_n45339_, new_n45340_, new_n45341_, new_n45342_, new_n45343_,
    new_n45344_, new_n45345_, new_n45346_, new_n45347_, new_n45348_,
    new_n45349_, new_n45350_, new_n45351_, new_n45352_, new_n45353_,
    new_n45354_, new_n45355_, new_n45356_, new_n45357_, new_n45358_,
    new_n45359_, new_n45360_, new_n45361_, new_n45362_, new_n45363_,
    new_n45364_, new_n45365_, new_n45366_, new_n45367_, new_n45368_,
    new_n45369_, new_n45370_, new_n45371_, new_n45372_, new_n45373_,
    new_n45374_, new_n45375_, new_n45376_, new_n45377_, new_n45378_,
    new_n45379_, new_n45380_, new_n45381_, new_n45382_, new_n45383_,
    new_n45384_, new_n45385_, new_n45386_, new_n45387_, new_n45388_,
    new_n45389_, new_n45390_, new_n45391_, new_n45392_, new_n45393_,
    new_n45394_, new_n45395_, new_n45396_, new_n45397_, new_n45398_,
    new_n45399_, new_n45400_, new_n45401_, new_n45402_, new_n45403_,
    new_n45404_, new_n45405_, new_n45406_, new_n45407_, new_n45408_,
    new_n45409_, new_n45410_, new_n45411_, new_n45412_, new_n45413_,
    new_n45414_, new_n45415_, new_n45416_, new_n45417_, new_n45418_,
    new_n45419_, new_n45420_, new_n45421_, new_n45422_, new_n45423_,
    new_n45424_, new_n45425_, new_n45426_, new_n45427_, new_n45428_,
    new_n45429_, new_n45430_, new_n45431_, new_n45432_, new_n45433_,
    new_n45434_, new_n45435_, new_n45436_, new_n45437_, new_n45438_,
    new_n45439_, new_n45440_, new_n45441_, new_n45442_, new_n45443_,
    new_n45444_, new_n45445_, new_n45446_, new_n45447_, new_n45448_,
    new_n45449_, new_n45450_, new_n45451_, new_n45452_, new_n45453_,
    new_n45454_, new_n45455_, new_n45456_, new_n45457_, new_n45458_,
    new_n45459_, new_n45460_, new_n45461_, new_n45462_, new_n45463_,
    new_n45464_, new_n45465_, new_n45466_, new_n45467_, new_n45468_,
    new_n45469_, new_n45470_, new_n45471_, new_n45472_, new_n45473_,
    new_n45474_, new_n45475_, new_n45476_, new_n45477_, new_n45478_,
    new_n45479_, new_n45480_, new_n45481_, new_n45482_, new_n45483_,
    new_n45484_, new_n45485_, new_n45486_, new_n45487_, new_n45488_,
    new_n45489_, new_n45490_, new_n45491_, new_n45492_, new_n45493_,
    new_n45494_, new_n45495_, new_n45496_, new_n45497_, new_n45498_,
    new_n45499_, new_n45500_, new_n45501_, new_n45502_, new_n45503_,
    new_n45504_, new_n45505_, new_n45506_, new_n45507_, new_n45508_,
    new_n45509_, new_n45510_, new_n45511_, new_n45512_, new_n45513_,
    new_n45514_, new_n45515_, new_n45516_, new_n45517_, new_n45518_,
    new_n45519_, new_n45520_, new_n45521_, new_n45522_, new_n45523_,
    new_n45524_, new_n45525_, new_n45526_, new_n45527_, new_n45528_,
    new_n45529_, new_n45530_, new_n45531_, new_n45532_, new_n45533_,
    new_n45534_, new_n45535_, new_n45536_, new_n45537_, new_n45538_,
    new_n45539_, new_n45540_, new_n45541_, new_n45542_, new_n45543_,
    new_n45544_, new_n45545_, new_n45546_, new_n45547_, new_n45548_,
    new_n45549_, new_n45550_, new_n45551_, new_n45552_, new_n45553_,
    new_n45554_, new_n45555_, new_n45556_, new_n45557_, new_n45558_,
    new_n45559_, new_n45560_, new_n45561_, new_n45562_, new_n45563_,
    new_n45564_, new_n45565_, new_n45566_, new_n45567_, new_n45568_,
    new_n45569_, new_n45570_, new_n45571_, new_n45572_, new_n45573_,
    new_n45574_, new_n45575_, new_n45576_, new_n45577_, new_n45578_,
    new_n45579_, new_n45580_, new_n45581_, new_n45582_, new_n45583_,
    new_n45584_, new_n45585_, new_n45586_, new_n45587_, new_n45588_,
    new_n45589_, new_n45590_, new_n45591_, new_n45592_, new_n45593_,
    new_n45594_, new_n45595_, new_n45596_, new_n45597_, new_n45598_,
    new_n45599_, new_n45600_, new_n45601_, new_n45602_, new_n45603_,
    new_n45604_, new_n45605_, new_n45606_, new_n45607_, new_n45608_,
    new_n45609_, new_n45610_, new_n45611_, new_n45612_, new_n45613_,
    new_n45614_, new_n45615_, new_n45616_, new_n45617_, new_n45618_,
    new_n45619_, new_n45620_, new_n45621_, new_n45622_, new_n45623_,
    new_n45624_, new_n45625_, new_n45626_, new_n45627_, new_n45628_,
    new_n45629_, new_n45630_, new_n45631_, new_n45632_, new_n45633_,
    new_n45634_, new_n45635_, new_n45636_, new_n45637_, new_n45638_,
    new_n45639_, new_n45640_, new_n45641_, new_n45642_, new_n45643_,
    new_n45644_, new_n45645_, new_n45646_, new_n45647_, new_n45648_,
    new_n45649_, new_n45650_, new_n45651_, new_n45652_, new_n45653_,
    new_n45654_, new_n45655_, new_n45656_, new_n45657_, new_n45658_,
    new_n45659_, new_n45660_, new_n45661_, new_n45662_, new_n45663_,
    new_n45664_, new_n45665_, new_n45666_, new_n45667_, new_n45668_,
    new_n45669_, new_n45670_, new_n45671_, new_n45672_, new_n45673_,
    new_n45674_, new_n45675_, new_n45676_, new_n45677_, new_n45678_,
    new_n45679_, new_n45680_, new_n45681_, new_n45682_, new_n45683_,
    new_n45684_, new_n45685_, new_n45686_, new_n45687_, new_n45688_,
    new_n45689_, new_n45690_, new_n45691_, new_n45692_, new_n45693_,
    new_n45694_, new_n45695_, new_n45696_, new_n45697_, new_n45698_,
    new_n45699_, new_n45700_, new_n45701_, new_n45702_, new_n45703_,
    new_n45704_, new_n45705_, new_n45706_, new_n45707_, new_n45708_,
    new_n45709_, new_n45710_, new_n45711_, new_n45712_, new_n45713_,
    new_n45714_, new_n45715_, new_n45716_, new_n45717_, new_n45718_,
    new_n45719_, new_n45720_, new_n45721_, new_n45722_, new_n45723_,
    new_n45724_, new_n45725_, new_n45726_, new_n45727_, new_n45728_,
    new_n45729_, new_n45730_, new_n45731_, new_n45732_, new_n45733_,
    new_n45734_, new_n45735_, new_n45736_, new_n45737_, new_n45738_,
    new_n45739_, new_n45740_, new_n45741_, new_n45742_, new_n45743_,
    new_n45744_, new_n45745_, new_n45746_, new_n45747_, new_n45748_,
    new_n45749_, new_n45750_, new_n45751_, new_n45752_, new_n45753_,
    new_n45754_, new_n45755_, new_n45756_, new_n45757_, new_n45758_,
    new_n45759_, new_n45760_, new_n45761_, new_n45762_, new_n45763_,
    new_n45764_, new_n45765_, new_n45766_, new_n45767_, new_n45768_,
    new_n45769_, new_n45770_, new_n45771_, new_n45772_, new_n45773_,
    new_n45774_, new_n45775_, new_n45776_, new_n45777_, new_n45778_,
    new_n45779_, new_n45780_, new_n45781_, new_n45782_, new_n45783_,
    new_n45784_, new_n45785_, new_n45786_, new_n45787_, new_n45788_,
    new_n45789_, new_n45790_, new_n45791_, new_n45792_, new_n45793_,
    new_n45794_, new_n45795_, new_n45796_, new_n45797_, new_n45798_,
    new_n45799_, new_n45800_, new_n45801_, new_n45802_, new_n45803_,
    new_n45804_, new_n45805_, new_n45806_, new_n45807_, new_n45808_,
    new_n45809_, new_n45810_, new_n45811_, new_n45812_, new_n45813_,
    new_n45814_, new_n45815_, new_n45816_, new_n45817_, new_n45818_,
    new_n45819_, new_n45820_, new_n45821_, new_n45822_, new_n45823_,
    new_n45824_, new_n45825_, new_n45826_, new_n45827_, new_n45828_,
    new_n45829_, new_n45830_, new_n45831_, new_n45832_, new_n45833_,
    new_n45834_, new_n45835_, new_n45836_, new_n45837_, new_n45838_,
    new_n45839_, new_n45840_, new_n45841_, new_n45842_, new_n45843_,
    new_n45844_, new_n45845_, new_n45846_, new_n45847_, new_n45848_,
    new_n45849_, new_n45850_, new_n45851_, new_n45852_, new_n45853_,
    new_n45854_, new_n45855_, new_n45856_, new_n45857_, new_n45858_,
    new_n45859_, new_n45860_, new_n45861_, new_n45862_, new_n45863_,
    new_n45864_, new_n45865_, new_n45866_, new_n45867_, new_n45868_,
    new_n45869_, new_n45870_, new_n45871_, new_n45872_, new_n45873_,
    new_n45874_, new_n45875_, new_n45876_, new_n45877_, new_n45878_,
    new_n45879_, new_n45880_, new_n45881_, new_n45882_, new_n45883_,
    new_n45884_, new_n45885_, new_n45886_, new_n45887_, new_n45888_,
    new_n45889_, new_n45890_, new_n45891_, new_n45892_, new_n45893_,
    new_n45894_, new_n45895_, new_n45896_, new_n45897_, new_n45898_,
    new_n45899_, new_n45900_, new_n45901_, new_n45902_, new_n45903_,
    new_n45904_, new_n45905_, new_n45906_, new_n45907_, new_n45908_,
    new_n45909_, new_n45910_, new_n45911_, new_n45912_, new_n45913_,
    new_n45914_, new_n45915_, new_n45916_, new_n45917_, new_n45918_,
    new_n45919_, new_n45920_, new_n45921_, new_n45922_, new_n45923_,
    new_n45924_, new_n45925_, new_n45926_, new_n45927_, new_n45928_,
    new_n45929_, new_n45930_, new_n45931_, new_n45932_, new_n45933_,
    new_n45934_, new_n45935_, new_n45936_, new_n45937_, new_n45938_,
    new_n45939_, new_n45940_, new_n45941_, new_n45942_, new_n45943_,
    new_n45944_, new_n45945_, new_n45946_, new_n45947_, new_n45948_,
    new_n45949_, new_n45950_, new_n45951_, new_n45952_, new_n45953_,
    new_n45954_, new_n45955_, new_n45956_, new_n45957_, new_n45958_,
    new_n45959_, new_n45960_, new_n45961_, new_n45962_, new_n45963_,
    new_n45964_, new_n45965_, new_n45966_, new_n45967_, new_n45968_,
    new_n45969_, new_n45970_, new_n45971_, new_n45972_, new_n45973_,
    new_n45974_, new_n45975_, new_n45976_, new_n45977_, new_n45978_,
    new_n45979_, new_n45980_, new_n45981_, new_n45982_, new_n45983_,
    new_n45984_, new_n45985_, new_n45986_, new_n45987_, new_n45988_,
    new_n45989_, new_n45990_, new_n45991_, new_n45992_, new_n45993_,
    new_n45994_, new_n45995_, new_n45996_, new_n45997_, new_n45998_,
    new_n45999_, new_n46000_, new_n46001_, new_n46002_, new_n46003_,
    new_n46004_, new_n46005_, new_n46006_, new_n46007_, new_n46008_,
    new_n46009_, new_n46010_, new_n46011_, new_n46012_, new_n46013_,
    new_n46014_, new_n46015_, new_n46016_, new_n46017_, new_n46018_,
    new_n46019_, new_n46020_, new_n46021_, new_n46022_, new_n46023_,
    new_n46024_, new_n46025_, new_n46026_, new_n46027_, new_n46028_,
    new_n46029_, new_n46030_, new_n46031_, new_n46032_, new_n46033_,
    new_n46034_, new_n46035_, new_n46036_, new_n46037_, new_n46038_,
    new_n46039_, new_n46040_, new_n46041_, new_n46042_, new_n46043_,
    new_n46044_, new_n46045_, new_n46046_, new_n46047_, new_n46048_,
    new_n46049_, new_n46050_, new_n46051_, new_n46052_, new_n46053_,
    new_n46054_, new_n46055_, new_n46056_, new_n46057_, new_n46058_,
    new_n46059_, new_n46060_, new_n46061_, new_n46062_, new_n46063_,
    new_n46064_, new_n46065_, new_n46066_, new_n46067_, new_n46068_,
    new_n46069_, new_n46070_, new_n46071_, new_n46072_, new_n46073_,
    new_n46074_, new_n46075_, new_n46076_, new_n46077_, new_n46078_,
    new_n46079_, new_n46080_, new_n46081_, new_n46082_, new_n46083_,
    new_n46084_, new_n46085_, new_n46086_, new_n46087_, new_n46088_,
    new_n46089_, new_n46090_, new_n46091_, new_n46092_, new_n46093_,
    new_n46094_, new_n46095_, new_n46096_, new_n46097_, new_n46098_,
    new_n46099_, new_n46100_, new_n46101_, new_n46102_, new_n46103_,
    new_n46104_, new_n46105_, new_n46106_, new_n46107_, new_n46108_,
    new_n46109_, new_n46110_, new_n46111_, new_n46112_, new_n46113_,
    new_n46114_, new_n46115_, new_n46116_, new_n46117_, new_n46118_,
    new_n46119_, new_n46120_, new_n46121_, new_n46122_, new_n46123_,
    new_n46124_, new_n46125_, new_n46126_, new_n46127_, new_n46128_,
    new_n46129_, new_n46130_, new_n46131_, new_n46132_, new_n46133_,
    new_n46134_, new_n46135_, new_n46136_, new_n46137_, new_n46138_,
    new_n46139_, new_n46140_, new_n46141_, new_n46142_, new_n46143_,
    new_n46144_, new_n46145_, new_n46146_, new_n46147_, new_n46148_,
    new_n46149_, new_n46150_, new_n46151_, new_n46152_, new_n46153_,
    new_n46154_, new_n46155_, new_n46156_, new_n46157_, new_n46158_,
    new_n46159_, new_n46160_, new_n46161_, new_n46162_, new_n46163_,
    new_n46164_, new_n46165_, new_n46166_, new_n46167_, new_n46168_,
    new_n46169_, new_n46170_, new_n46171_, new_n46172_, new_n46173_,
    new_n46174_, new_n46175_, new_n46176_, new_n46177_, new_n46178_,
    new_n46179_, new_n46180_, new_n46181_, new_n46182_, new_n46183_,
    new_n46184_, new_n46185_, new_n46186_, new_n46187_, new_n46188_,
    new_n46189_, new_n46190_, new_n46191_, new_n46192_, new_n46193_,
    new_n46194_, new_n46195_, new_n46196_, new_n46197_, new_n46198_,
    new_n46199_, new_n46200_, new_n46201_, new_n46202_, new_n46203_,
    new_n46204_, new_n46205_, new_n46206_, new_n46207_, new_n46208_,
    new_n46209_, new_n46210_, new_n46211_, new_n46212_, new_n46213_,
    new_n46214_, new_n46215_, new_n46216_, new_n46217_, new_n46218_,
    new_n46219_, new_n46220_, new_n46221_, new_n46222_, new_n46223_,
    new_n46224_, new_n46225_, new_n46226_, new_n46227_, new_n46228_,
    new_n46229_, new_n46230_, new_n46231_, new_n46232_, new_n46233_,
    new_n46234_, new_n46235_, new_n46236_, new_n46237_, new_n46238_,
    new_n46239_, new_n46240_, new_n46241_, new_n46242_, new_n46243_,
    new_n46244_, new_n46245_, new_n46246_, new_n46247_, new_n46248_,
    new_n46249_, new_n46250_, new_n46251_, new_n46252_, new_n46253_,
    new_n46254_, new_n46255_, new_n46256_, new_n46257_, new_n46258_,
    new_n46259_, new_n46260_, new_n46261_, new_n46262_, new_n46263_,
    new_n46264_, new_n46265_, new_n46266_, new_n46267_, new_n46268_,
    new_n46269_, new_n46270_, new_n46271_, new_n46272_, new_n46273_,
    new_n46274_, new_n46275_, new_n46276_, new_n46277_, new_n46278_,
    new_n46279_, new_n46280_, new_n46281_, new_n46282_, new_n46283_,
    new_n46284_, new_n46285_, new_n46286_, new_n46287_, new_n46288_,
    new_n46289_, new_n46290_, new_n46291_, new_n46292_, new_n46293_,
    new_n46294_, new_n46295_, new_n46296_, new_n46297_, new_n46298_,
    new_n46299_, new_n46300_, new_n46301_, new_n46302_, new_n46303_,
    new_n46304_, new_n46305_, new_n46306_, new_n46307_, new_n46308_,
    new_n46309_, new_n46310_, new_n46311_, new_n46312_, new_n46313_,
    new_n46314_, new_n46315_, new_n46316_, new_n46317_, new_n46318_,
    new_n46319_, new_n46320_, new_n46321_, new_n46322_, new_n46323_,
    new_n46324_, new_n46325_, new_n46326_, new_n46327_, new_n46328_,
    new_n46329_, new_n46330_, new_n46331_, new_n46332_, new_n46333_,
    new_n46334_, new_n46335_, new_n46336_, new_n46337_, new_n46338_,
    new_n46339_, new_n46340_, new_n46341_, new_n46342_, new_n46343_,
    new_n46344_, new_n46345_, new_n46346_, new_n46347_, new_n46348_,
    new_n46349_, new_n46350_, new_n46351_, new_n46352_, new_n46353_,
    new_n46354_, new_n46355_, new_n46356_, new_n46357_, new_n46358_,
    new_n46359_, new_n46360_, new_n46361_, new_n46362_, new_n46363_,
    new_n46364_, new_n46365_, new_n46366_, new_n46367_, new_n46368_,
    new_n46369_, new_n46370_, new_n46371_, new_n46372_, new_n46373_,
    new_n46374_, new_n46375_, new_n46376_, new_n46377_, new_n46378_,
    new_n46379_, new_n46380_, new_n46381_, new_n46382_, new_n46383_,
    new_n46384_, new_n46385_, new_n46386_, new_n46387_, new_n46388_,
    new_n46389_, new_n46390_, new_n46391_, new_n46392_, new_n46393_,
    new_n46394_, new_n46395_, new_n46396_, new_n46397_, new_n46398_,
    new_n46399_, new_n46400_, new_n46401_, new_n46402_, new_n46403_,
    new_n46404_, new_n46405_, new_n46406_, new_n46407_, new_n46408_,
    new_n46409_, new_n46410_, new_n46411_, new_n46412_, new_n46413_,
    new_n46414_, new_n46415_, new_n46416_, new_n46417_, new_n46418_,
    new_n46419_, new_n46420_, new_n46421_, new_n46422_, new_n46423_,
    new_n46424_, new_n46425_, new_n46426_, new_n46427_, new_n46428_,
    new_n46429_, new_n46430_, new_n46431_, new_n46432_, new_n46433_,
    new_n46434_, new_n46435_, new_n46436_, new_n46437_, new_n46438_,
    new_n46439_, new_n46440_, new_n46441_, new_n46442_, new_n46443_,
    new_n46444_, new_n46445_, new_n46446_, new_n46447_, new_n46448_,
    new_n46449_, new_n46450_, new_n46451_, new_n46452_, new_n46453_,
    new_n46454_, new_n46455_, new_n46456_, new_n46457_, new_n46458_,
    new_n46459_, new_n46460_, new_n46461_, new_n46462_, new_n46463_,
    new_n46464_, new_n46465_, new_n46466_, new_n46467_, new_n46468_,
    new_n46469_, new_n46470_, new_n46471_, new_n46472_, new_n46473_,
    new_n46474_, new_n46475_, new_n46476_, new_n46477_, new_n46478_,
    new_n46479_, new_n46480_, new_n46481_, new_n46482_, new_n46483_,
    new_n46484_, new_n46485_, new_n46486_, new_n46487_, new_n46488_,
    new_n46489_, new_n46490_, new_n46491_, new_n46492_, new_n46493_,
    new_n46494_, new_n46495_, new_n46496_, new_n46497_, new_n46498_,
    new_n46499_, new_n46500_, new_n46501_, new_n46502_, new_n46503_,
    new_n46504_, new_n46505_, new_n46506_, new_n46507_, new_n46508_,
    new_n46509_, new_n46510_, new_n46511_, new_n46512_, new_n46513_,
    new_n46514_, new_n46515_, new_n46516_, new_n46517_, new_n46518_,
    new_n46519_, new_n46520_, new_n46521_, new_n46522_, new_n46523_,
    new_n46524_, new_n46525_, new_n46526_, new_n46527_, new_n46528_,
    new_n46529_, new_n46530_, new_n46531_, new_n46532_, new_n46533_,
    new_n46534_, new_n46535_, new_n46536_, new_n46537_, new_n46538_,
    new_n46539_, new_n46540_, new_n46541_, new_n46542_, new_n46543_,
    new_n46544_, new_n46545_, new_n46546_, new_n46547_, new_n46548_,
    new_n46549_, new_n46550_, new_n46551_, new_n46552_, new_n46553_,
    new_n46554_, new_n46555_, new_n46556_, new_n46557_, new_n46558_,
    new_n46559_, new_n46560_, new_n46561_, new_n46562_, new_n46563_,
    new_n46564_, new_n46565_, new_n46566_, new_n46567_, new_n46568_,
    new_n46569_, new_n46570_, new_n46571_, new_n46572_, new_n46573_,
    new_n46574_, new_n46575_, new_n46576_, new_n46577_, new_n46578_,
    new_n46579_, new_n46580_, new_n46581_, new_n46582_, new_n46583_,
    new_n46584_, new_n46585_, new_n46586_, new_n46587_, new_n46588_,
    new_n46589_, new_n46590_, new_n46591_, new_n46592_, new_n46593_,
    new_n46594_, new_n46595_, new_n46596_, new_n46597_, new_n46598_,
    new_n46599_, new_n46600_, new_n46601_, new_n46602_, new_n46603_,
    new_n46604_, new_n46605_, new_n46606_, new_n46607_, new_n46608_,
    new_n46609_, new_n46610_, new_n46611_, new_n46612_, new_n46613_,
    new_n46614_, new_n46615_, new_n46616_, new_n46617_, new_n46618_,
    new_n46619_, new_n46620_, new_n46621_, new_n46622_, new_n46623_,
    new_n46624_, new_n46625_, new_n46626_, new_n46627_, new_n46628_,
    new_n46629_, new_n46630_, new_n46631_, new_n46632_, new_n46633_,
    new_n46634_, new_n46635_, new_n46636_, new_n46637_, new_n46638_,
    new_n46639_, new_n46640_, new_n46641_, new_n46642_, new_n46643_,
    new_n46644_, new_n46645_, new_n46646_, new_n46647_, new_n46648_,
    new_n46649_, new_n46650_, new_n46651_, new_n46652_, new_n46653_,
    new_n46654_, new_n46655_, new_n46656_, new_n46657_, new_n46658_,
    new_n46659_, new_n46660_, new_n46661_, new_n46662_, new_n46663_,
    new_n46664_, new_n46665_, new_n46666_, new_n46667_, new_n46668_,
    new_n46669_, new_n46670_, new_n46671_, new_n46672_, new_n46673_,
    new_n46674_, new_n46675_, new_n46676_, new_n46677_, new_n46678_,
    new_n46679_, new_n46680_, new_n46681_, new_n46682_, new_n46683_,
    new_n46684_, new_n46685_, new_n46686_, new_n46687_, new_n46688_,
    new_n46689_, new_n46690_, new_n46691_, new_n46692_, new_n46693_,
    new_n46694_, new_n46695_, new_n46696_, new_n46697_, new_n46698_,
    new_n46699_, new_n46700_, new_n46701_, new_n46702_, new_n46703_,
    new_n46704_, new_n46705_, new_n46706_, new_n46707_, new_n46708_,
    new_n46709_, new_n46710_, new_n46711_, new_n46712_, new_n46713_,
    new_n46714_, new_n46715_, new_n46716_, new_n46717_, new_n46718_,
    new_n46719_, new_n46720_, new_n46721_, new_n46722_, new_n46723_,
    new_n46724_, new_n46725_, new_n46726_, new_n46727_, new_n46728_,
    new_n46729_, new_n46730_, new_n46731_, new_n46732_, new_n46733_,
    new_n46734_, new_n46735_, new_n46736_, new_n46737_, new_n46738_,
    new_n46739_, new_n46740_, new_n46741_, new_n46742_, new_n46743_,
    new_n46744_, new_n46745_, new_n46746_, new_n46747_, new_n46748_,
    new_n46749_, new_n46750_, new_n46751_, new_n46752_, new_n46753_,
    new_n46754_, new_n46755_, new_n46756_, new_n46757_, new_n46758_,
    new_n46759_, new_n46760_, new_n46761_, new_n46762_, new_n46763_,
    new_n46764_, new_n46765_, new_n46766_, new_n46767_, new_n46768_,
    new_n46769_, new_n46770_, new_n46771_, new_n46772_, new_n46773_,
    new_n46774_, new_n46775_, new_n46776_, new_n46777_, new_n46778_,
    new_n46779_, new_n46780_, new_n46781_, new_n46782_, new_n46783_,
    new_n46784_, new_n46785_, new_n46786_, new_n46787_, new_n46788_,
    new_n46789_, new_n46790_, new_n46791_, new_n46792_, new_n46793_,
    new_n46794_, new_n46795_, new_n46796_, new_n46797_, new_n46798_,
    new_n46799_, new_n46800_, new_n46801_, new_n46802_, new_n46803_,
    new_n46804_, new_n46805_, new_n46806_, new_n46807_, new_n46808_,
    new_n46809_, new_n46810_, new_n46811_, new_n46812_, new_n46813_,
    new_n46814_, new_n46815_, new_n46816_, new_n46817_, new_n46818_,
    new_n46819_, new_n46820_, new_n46821_, new_n46822_, new_n46823_,
    new_n46824_, new_n46825_, new_n46826_, new_n46827_, new_n46828_,
    new_n46829_, new_n46830_, new_n46831_, new_n46832_, new_n46833_,
    new_n46834_, new_n46835_, new_n46836_, new_n46837_, new_n46838_,
    new_n46839_, new_n46840_, new_n46841_, new_n46842_, new_n46843_,
    new_n46844_, new_n46845_, new_n46846_, new_n46847_, new_n46848_,
    new_n46849_, new_n46850_, new_n46851_, new_n46852_, new_n46853_,
    new_n46854_, new_n46855_, new_n46856_, new_n46857_, new_n46858_,
    new_n46859_, new_n46860_, new_n46861_, new_n46862_, new_n46863_,
    new_n46864_, new_n46865_, new_n46866_, new_n46867_, new_n46868_,
    new_n46869_, new_n46870_, new_n46871_, new_n46872_, new_n46873_,
    new_n46874_, new_n46875_, new_n46876_, new_n46877_, new_n46878_,
    new_n46879_, new_n46880_, new_n46881_, new_n46882_, new_n46883_,
    new_n46884_, new_n46885_, new_n46886_, new_n46887_, new_n46888_,
    new_n46889_, new_n46890_, new_n46891_, new_n46892_, new_n46893_,
    new_n46894_, new_n46895_, new_n46896_, new_n46897_, new_n46898_,
    new_n46899_, new_n46900_, new_n46901_, new_n46902_, new_n46903_,
    new_n46904_, new_n46905_, new_n46906_, new_n46907_, new_n46908_,
    new_n46909_, new_n46910_, new_n46911_, new_n46912_, new_n46913_,
    new_n46914_, new_n46915_, new_n46916_, new_n46917_, new_n46918_,
    new_n46919_, new_n46920_, new_n46921_, new_n46922_, new_n46923_,
    new_n46924_, new_n46925_, new_n46926_, new_n46927_, new_n46928_,
    new_n46929_, new_n46930_, new_n46931_, new_n46932_, new_n46933_,
    new_n46934_, new_n46935_, new_n46936_, new_n46937_, new_n46938_,
    new_n46939_, new_n46940_, new_n46941_, new_n46942_, new_n46943_,
    new_n46944_, new_n46945_, new_n46946_, new_n46947_, new_n46948_,
    new_n46949_, new_n46950_, new_n46951_, new_n46952_, new_n46953_,
    new_n46954_, new_n46955_, new_n46956_, new_n46957_, new_n46958_,
    new_n46959_, new_n46960_, new_n46961_, new_n46962_, new_n46963_,
    new_n46964_, new_n46965_, new_n46966_, new_n46967_, new_n46968_,
    new_n46969_, new_n46970_, new_n46971_, new_n46972_, new_n46973_,
    new_n46974_, new_n46975_, new_n46976_, new_n46977_, new_n46978_,
    new_n46979_, new_n46980_, new_n46981_, new_n46982_, new_n46983_,
    new_n46984_, new_n46985_, new_n46986_, new_n46987_, new_n46988_,
    new_n46989_, new_n46990_, new_n46991_, new_n46992_, new_n46993_,
    new_n46994_, new_n46995_, new_n46996_, new_n46997_, new_n46998_,
    new_n46999_, new_n47000_, new_n47001_, new_n47002_, new_n47003_,
    new_n47004_, new_n47005_, new_n47006_, new_n47007_, new_n47008_,
    new_n47009_, new_n47010_, new_n47011_, new_n47012_, new_n47013_,
    new_n47014_, new_n47015_, new_n47016_, new_n47017_, new_n47018_,
    new_n47019_, new_n47020_, new_n47021_, new_n47022_, new_n47023_,
    new_n47024_, new_n47025_, new_n47026_, new_n47027_, new_n47028_,
    new_n47029_, new_n47030_, new_n47031_, new_n47032_, new_n47033_,
    new_n47034_, new_n47035_, new_n47036_, new_n47037_, new_n47038_,
    new_n47039_, new_n47040_, new_n47041_, new_n47042_, new_n47043_,
    new_n47044_, new_n47045_, new_n47046_, new_n47047_, new_n47048_,
    new_n47049_, new_n47050_, new_n47051_, new_n47052_, new_n47053_,
    new_n47054_, new_n47055_, new_n47056_, new_n47057_, new_n47058_,
    new_n47059_, new_n47060_, new_n47061_, new_n47062_, new_n47063_,
    new_n47064_, new_n47065_, new_n47066_, new_n47067_, new_n47068_,
    new_n47069_, new_n47070_, new_n47071_, new_n47072_, new_n47073_,
    new_n47074_, new_n47075_, new_n47076_, new_n47077_, new_n47078_,
    new_n47079_, new_n47080_, new_n47081_, new_n47082_, new_n47083_,
    new_n47084_, new_n47085_, new_n47086_, new_n47087_, new_n47088_,
    new_n47089_, new_n47090_, new_n47091_, new_n47092_, new_n47093_,
    new_n47094_, new_n47095_, new_n47096_, new_n47097_, new_n47098_,
    new_n47099_, new_n47100_, new_n47101_, new_n47102_, new_n47103_,
    new_n47104_, new_n47105_, new_n47106_, new_n47107_, new_n47108_,
    new_n47109_, new_n47110_, new_n47111_, new_n47112_, new_n47113_,
    new_n47114_, new_n47115_, new_n47116_, new_n47117_, new_n47118_,
    new_n47119_, new_n47120_, new_n47121_, new_n47122_, new_n47123_,
    new_n47124_, new_n47125_, new_n47126_, new_n47127_, new_n47128_,
    new_n47129_, new_n47130_, new_n47131_, new_n47132_, new_n47133_,
    new_n47134_, new_n47135_, new_n47136_, new_n47137_, new_n47138_,
    new_n47139_, new_n47140_, new_n47141_, new_n47142_, new_n47143_,
    new_n47144_, new_n47145_, new_n47146_, new_n47147_, new_n47148_,
    new_n47149_, new_n47150_, new_n47151_, new_n47152_, new_n47153_,
    new_n47154_, new_n47155_, new_n47156_, new_n47157_, new_n47158_,
    new_n47159_, new_n47160_, new_n47161_, new_n47162_, new_n47163_,
    new_n47164_, new_n47165_, new_n47166_, new_n47167_, new_n47168_,
    new_n47169_, new_n47170_, new_n47171_, new_n47172_, new_n47173_,
    new_n47174_, new_n47175_, new_n47176_, new_n47177_, new_n47178_,
    new_n47179_, new_n47180_, new_n47181_, new_n47182_, new_n47183_,
    new_n47184_, new_n47185_, new_n47186_, new_n47187_, new_n47188_,
    new_n47189_, new_n47190_, new_n47191_, new_n47192_, new_n47193_,
    new_n47194_, new_n47195_, new_n47196_, new_n47197_, new_n47198_,
    new_n47199_, new_n47200_, new_n47201_, new_n47202_, new_n47203_,
    new_n47204_, new_n47205_, new_n47206_, new_n47207_, new_n47208_,
    new_n47209_, new_n47210_, new_n47211_, new_n47212_, new_n47213_,
    new_n47214_, new_n47215_, new_n47216_, new_n47217_, new_n47218_,
    new_n47219_, new_n47220_, new_n47221_, new_n47222_, new_n47223_,
    new_n47224_, new_n47225_, new_n47226_, new_n47227_, new_n47228_,
    new_n47229_, new_n47230_, new_n47231_, new_n47232_, new_n47233_,
    new_n47234_, new_n47235_, new_n47236_, new_n47237_, new_n47238_,
    new_n47239_, new_n47240_, new_n47241_, new_n47242_, new_n47243_,
    new_n47244_, new_n47245_, new_n47246_, new_n47247_, new_n47248_,
    new_n47249_, new_n47250_, new_n47251_, new_n47252_, new_n47253_,
    new_n47254_, new_n47255_, new_n47256_, new_n47257_, new_n47258_,
    new_n47259_, new_n47260_, new_n47261_, new_n47262_, new_n47263_,
    new_n47264_, new_n47265_, new_n47266_, new_n47267_, new_n47268_,
    new_n47269_, new_n47270_, new_n47271_, new_n47272_, new_n47273_,
    new_n47274_, new_n47275_, new_n47276_, new_n47277_, new_n47278_,
    new_n47279_, new_n47280_, new_n47281_, new_n47282_, new_n47283_,
    new_n47284_, new_n47285_, new_n47286_, new_n47287_, new_n47288_,
    new_n47289_, new_n47290_, new_n47291_, new_n47292_, new_n47293_,
    new_n47294_, new_n47295_, new_n47296_, new_n47297_, new_n47298_,
    new_n47299_, new_n47300_, new_n47301_, new_n47302_, new_n47303_,
    new_n47304_, new_n47305_, new_n47306_, new_n47307_, new_n47308_,
    new_n47309_, new_n47310_, new_n47311_, new_n47312_, new_n47313_,
    new_n47314_, new_n47315_, new_n47316_, new_n47317_, new_n47318_,
    new_n47319_, new_n47320_, new_n47321_, new_n47322_, new_n47323_,
    new_n47324_, new_n47325_, new_n47326_, new_n47327_, new_n47328_,
    new_n47329_, new_n47330_, new_n47331_, new_n47332_, new_n47333_,
    new_n47334_, new_n47335_, new_n47336_, new_n47337_, new_n47338_,
    new_n47339_, new_n47340_, new_n47341_, new_n47342_, new_n47343_,
    new_n47344_, new_n47345_, new_n47346_, new_n47347_, new_n47348_,
    new_n47349_, new_n47350_, new_n47351_, new_n47352_, new_n47353_,
    new_n47354_, new_n47355_, new_n47356_, new_n47357_, new_n47358_,
    new_n47359_, new_n47360_, new_n47361_, new_n47362_, new_n47363_,
    new_n47364_, new_n47365_, new_n47366_, new_n47367_, new_n47368_,
    new_n47369_, new_n47370_, new_n47371_, new_n47372_, new_n47373_,
    new_n47374_, new_n47375_, new_n47376_, new_n47377_, new_n47378_,
    new_n47379_, new_n47380_, new_n47381_, new_n47382_, new_n47383_,
    new_n47384_, new_n47385_, new_n47386_, new_n47387_, new_n47388_,
    new_n47389_, new_n47390_, new_n47391_, new_n47392_, new_n47393_,
    new_n47394_, new_n47395_, new_n47396_, new_n47397_, new_n47398_,
    new_n47399_, new_n47400_, new_n47401_, new_n47402_, new_n47403_,
    new_n47404_, new_n47405_, new_n47406_, new_n47407_, new_n47408_,
    new_n47409_, new_n47410_, new_n47411_, new_n47412_, new_n47413_,
    new_n47414_, new_n47415_, new_n47416_, new_n47417_, new_n47418_,
    new_n47419_, new_n47420_, new_n47421_, new_n47422_, new_n47423_,
    new_n47424_, new_n47425_, new_n47426_, new_n47427_, new_n47428_,
    new_n47429_, new_n47430_, new_n47431_, new_n47432_, new_n47433_,
    new_n47434_, new_n47435_, new_n47436_, new_n47437_, new_n47438_,
    new_n47439_, new_n47440_, new_n47441_, new_n47442_, new_n47443_,
    new_n47444_, new_n47445_, new_n47446_, new_n47447_, new_n47448_,
    new_n47449_, new_n47450_, new_n47451_, new_n47452_, new_n47453_,
    new_n47454_, new_n47455_, new_n47456_, new_n47457_, new_n47458_,
    new_n47459_, new_n47460_, new_n47461_, new_n47462_, new_n47463_,
    new_n47464_, new_n47465_, new_n47466_, new_n47467_, new_n47468_,
    new_n47469_, new_n47470_, new_n47471_, new_n47472_, new_n47473_,
    new_n47474_, new_n47475_, new_n47476_, new_n47477_, new_n47478_,
    new_n47479_, new_n47480_, new_n47481_, new_n47482_, new_n47483_,
    new_n47484_, new_n47485_, new_n47486_, new_n47487_, new_n47488_,
    new_n47489_, new_n47490_, new_n47491_, new_n47492_, new_n47493_,
    new_n47494_, new_n47495_, new_n47496_, new_n47497_, new_n47498_,
    new_n47499_, new_n47500_, new_n47501_, new_n47502_, new_n47503_,
    new_n47504_, new_n47505_, new_n47506_, new_n47507_, new_n47508_,
    new_n47509_, new_n47510_, new_n47511_, new_n47512_, new_n47513_,
    new_n47514_, new_n47515_, new_n47516_, new_n47517_, new_n47518_,
    new_n47519_, new_n47520_, new_n47521_, new_n47522_, new_n47523_,
    new_n47524_, new_n47525_, new_n47526_, new_n47527_, new_n47528_,
    new_n47529_, new_n47530_, new_n47531_, new_n47532_, new_n47533_,
    new_n47534_, new_n47535_, new_n47536_, new_n47537_, new_n47538_,
    new_n47539_, new_n47540_, new_n47541_, new_n47542_, new_n47543_,
    new_n47544_, new_n47545_, new_n47546_, new_n47547_, new_n47548_,
    new_n47549_, new_n47550_, new_n47551_, new_n47552_, new_n47553_,
    new_n47554_, new_n47555_, new_n47556_, new_n47557_, new_n47558_,
    new_n47559_, new_n47560_, new_n47561_, new_n47562_, new_n47563_,
    new_n47564_, new_n47565_, new_n47566_, new_n47567_, new_n47568_,
    new_n47569_, new_n47570_, new_n47571_, new_n47572_, new_n47573_,
    new_n47574_, new_n47575_, new_n47576_, new_n47577_, new_n47578_,
    new_n47579_, new_n47580_, new_n47581_, new_n47582_, new_n47583_,
    new_n47584_, new_n47585_, new_n47586_, new_n47587_, new_n47588_,
    new_n47589_, new_n47590_, new_n47591_, new_n47592_, new_n47593_,
    new_n47594_, new_n47595_, new_n47596_, new_n47597_, new_n47598_,
    new_n47599_, new_n47600_, new_n47601_, new_n47602_, new_n47603_,
    new_n47604_, new_n47605_, new_n47606_, new_n47607_, new_n47608_,
    new_n47609_, new_n47610_, new_n47611_, new_n47612_, new_n47613_,
    new_n47614_, new_n47615_, new_n47616_, new_n47617_, new_n47618_,
    new_n47619_, new_n47620_, new_n47621_, new_n47622_, new_n47623_,
    new_n47624_, new_n47625_, new_n47626_, new_n47627_, new_n47628_,
    new_n47629_, new_n47630_, new_n47631_, new_n47632_, new_n47633_,
    new_n47634_, new_n47635_, new_n47636_, new_n47637_, new_n47638_,
    new_n47639_, new_n47640_, new_n47641_, new_n47642_, new_n47643_,
    new_n47644_, new_n47645_, new_n47646_, new_n47647_, new_n47648_,
    new_n47649_, new_n47650_, new_n47651_, new_n47652_, new_n47653_,
    new_n47654_, new_n47655_, new_n47656_, new_n47657_, new_n47658_,
    new_n47659_, new_n47660_, new_n47661_, new_n47662_, new_n47663_,
    new_n47664_, new_n47665_, new_n47666_, new_n47667_, new_n47668_,
    new_n47669_, new_n47670_, new_n47671_, new_n47672_, new_n47673_,
    new_n47674_, new_n47675_, new_n47676_, new_n47677_, new_n47678_,
    new_n47679_, new_n47680_, new_n47681_, new_n47682_, new_n47683_,
    new_n47684_, new_n47685_, new_n47686_, new_n47687_, new_n47688_,
    new_n47689_, new_n47690_, new_n47691_, new_n47692_, new_n47693_,
    new_n47694_, new_n47695_, new_n47696_, new_n47697_, new_n47698_,
    new_n47699_, new_n47700_, new_n47701_, new_n47702_, new_n47703_,
    new_n47704_, new_n47705_, new_n47706_, new_n47707_, new_n47708_,
    new_n47709_, new_n47710_, new_n47711_, new_n47712_, new_n47713_,
    new_n47714_, new_n47715_, new_n47716_, new_n47717_, new_n47718_,
    new_n47719_, new_n47720_, new_n47721_, new_n47722_, new_n47723_,
    new_n47724_, new_n47725_, new_n47726_, new_n47727_, new_n47728_,
    new_n47729_, new_n47730_, new_n47731_, new_n47732_, new_n47733_,
    new_n47734_, new_n47735_, new_n47736_, new_n47737_, new_n47738_,
    new_n47739_, new_n47740_, new_n47741_, new_n47742_, new_n47743_,
    new_n47744_, new_n47745_, new_n47746_, new_n47747_, new_n47748_,
    new_n47749_, new_n47750_, new_n47751_, new_n47752_, new_n47753_,
    new_n47754_, new_n47755_, new_n47756_, new_n47757_, new_n47758_,
    new_n47759_, new_n47760_, new_n47761_, new_n47762_, new_n47763_,
    new_n47764_, new_n47765_, new_n47766_, new_n47767_, new_n47768_,
    new_n47769_, new_n47770_, new_n47771_, new_n47772_, new_n47773_,
    new_n47774_, new_n47775_, new_n47776_, new_n47777_, new_n47778_,
    new_n47779_, new_n47780_, new_n47781_, new_n47782_, new_n47783_,
    new_n47784_, new_n47785_, new_n47786_, new_n47787_, new_n47788_,
    new_n47789_, new_n47790_, new_n47791_, new_n47792_, new_n47793_,
    new_n47794_, new_n47795_, new_n47796_, new_n47797_, new_n47798_,
    new_n47799_, new_n47800_, new_n47801_, new_n47802_, new_n47803_,
    new_n47804_, new_n47805_, new_n47806_, new_n47807_, new_n47808_,
    new_n47809_, new_n47810_, new_n47811_, new_n47812_, new_n47813_,
    new_n47814_, new_n47815_, new_n47816_, new_n47817_, new_n47818_,
    new_n47819_, new_n47820_, new_n47821_, new_n47822_, new_n47823_,
    new_n47824_, new_n47825_, new_n47826_, new_n47827_, new_n47828_,
    new_n47829_, new_n47830_, new_n47831_, new_n47832_, new_n47833_,
    new_n47834_, new_n47835_, new_n47836_, new_n47837_, new_n47838_,
    new_n47839_, new_n47840_, new_n47841_, new_n47842_, new_n47843_,
    new_n47844_, new_n47845_, new_n47846_, new_n47847_, new_n47848_,
    new_n47849_, new_n47850_, new_n47851_, new_n47852_, new_n47853_,
    new_n47854_, new_n47855_, new_n47856_, new_n47857_, new_n47858_,
    new_n47859_, new_n47860_, new_n47861_, new_n47862_, new_n47863_,
    new_n47864_, new_n47865_, new_n47866_, new_n47867_, new_n47868_,
    new_n47869_, new_n47870_, new_n47871_, new_n47872_, new_n47873_,
    new_n47874_, new_n47875_, new_n47876_, new_n47877_, new_n47878_,
    new_n47879_, new_n47880_, new_n47881_, new_n47882_, new_n47883_,
    new_n47884_, new_n47885_, new_n47886_, new_n47887_, new_n47888_,
    new_n47889_, new_n47890_, new_n47891_, new_n47892_, new_n47893_,
    new_n47894_, new_n47895_, new_n47896_, new_n47897_, new_n47898_,
    new_n47899_, new_n47900_, new_n47901_, new_n47902_, new_n47903_,
    new_n47904_, new_n47905_, new_n47906_, new_n47907_, new_n47908_,
    new_n47909_, new_n47910_, new_n47911_, new_n47912_, new_n47913_,
    new_n47914_, new_n47915_, new_n47916_, new_n47917_, new_n47918_,
    new_n47919_, new_n47920_, new_n47921_, new_n47922_, new_n47923_,
    new_n47924_, new_n47925_, new_n47926_, new_n47927_, new_n47928_,
    new_n47929_, new_n47930_, new_n47931_, new_n47932_, new_n47933_,
    new_n47934_, new_n47935_, new_n47936_, new_n47937_, new_n47938_,
    new_n47939_, new_n47940_, new_n47941_, new_n47942_, new_n47943_,
    new_n47944_, new_n47945_, new_n47946_, new_n47947_, new_n47948_,
    new_n47949_, new_n47950_, new_n47951_, new_n47952_, new_n47953_,
    new_n47954_, new_n47955_, new_n47956_, new_n47957_, new_n47958_,
    new_n47959_, new_n47960_, new_n47961_, new_n47962_, new_n47963_,
    new_n47964_, new_n47965_, new_n47966_, new_n47967_, new_n47968_,
    new_n47969_, new_n47970_, new_n47971_, new_n47972_, new_n47973_,
    new_n47974_, new_n47975_, new_n47976_, new_n47977_, new_n47978_,
    new_n47979_, new_n47980_, new_n47981_, new_n47982_, new_n47983_,
    new_n47984_, new_n47985_, new_n47986_, new_n47987_, new_n47988_,
    new_n47989_, new_n47990_, new_n47991_, new_n47992_, new_n47993_,
    new_n47994_, new_n47995_, new_n47996_, new_n47997_, new_n47998_,
    new_n47999_, new_n48000_, new_n48001_, new_n48002_, new_n48003_,
    new_n48004_, new_n48005_, new_n48006_, new_n48007_, new_n48008_,
    new_n48009_, new_n48010_, new_n48011_, new_n48012_, new_n48013_,
    new_n48014_, new_n48015_, new_n48016_, new_n48017_, new_n48018_,
    new_n48019_, new_n48020_, new_n48021_, new_n48022_, new_n48023_,
    new_n48024_, new_n48025_, new_n48026_, new_n48027_, new_n48028_,
    new_n48029_, new_n48030_, new_n48031_, new_n48032_, new_n48033_,
    new_n48034_, new_n48035_, new_n48036_, new_n48037_, new_n48038_,
    new_n48039_, new_n48040_, new_n48041_, new_n48042_, new_n48043_,
    new_n48044_, new_n48045_, new_n48046_, new_n48047_, new_n48048_,
    new_n48049_, new_n48050_, new_n48051_, new_n48052_, new_n48053_,
    new_n48054_, new_n48055_, new_n48056_, new_n48057_, new_n48058_,
    new_n48059_, new_n48060_, new_n48061_, new_n48062_, new_n48063_,
    new_n48064_, new_n48065_, new_n48066_, new_n48067_, new_n48068_,
    new_n48069_, new_n48070_, new_n48071_, new_n48072_, new_n48073_,
    new_n48074_, new_n48075_, new_n48076_, new_n48077_, new_n48078_,
    new_n48079_, new_n48080_, new_n48081_, new_n48082_, new_n48083_,
    new_n48084_, new_n48085_, new_n48086_, new_n48087_, new_n48088_,
    new_n48089_, new_n48090_, new_n48091_, new_n48092_, new_n48093_,
    new_n48094_, new_n48095_, new_n48096_, new_n48097_, new_n48098_,
    new_n48099_, new_n48100_, new_n48101_, new_n48102_, new_n48103_,
    new_n48104_, new_n48105_, new_n48106_, new_n48107_, new_n48108_,
    new_n48109_, new_n48110_, new_n48111_, new_n48112_, new_n48113_,
    new_n48114_, new_n48115_, new_n48116_, new_n48117_, new_n48118_,
    new_n48119_, new_n48120_, new_n48121_, new_n48122_, new_n48123_,
    new_n48124_, new_n48125_, new_n48126_, new_n48127_, new_n48128_,
    new_n48129_, new_n48130_, new_n48131_, new_n48132_, new_n48133_,
    new_n48134_, new_n48135_, new_n48136_, new_n48137_, new_n48138_,
    new_n48139_, new_n48140_, new_n48141_, new_n48142_, new_n48143_,
    new_n48144_, new_n48145_, new_n48146_, new_n48147_, new_n48148_,
    new_n48149_, new_n48150_, new_n48151_, new_n48152_, new_n48153_,
    new_n48154_, new_n48155_, new_n48156_, new_n48157_, new_n48158_,
    new_n48159_, new_n48160_, new_n48161_, new_n48162_, new_n48163_,
    new_n48164_, new_n48165_, new_n48166_, new_n48167_, new_n48168_,
    new_n48169_, new_n48170_, new_n48171_, new_n48172_, new_n48173_,
    new_n48174_, new_n48175_, new_n48176_, new_n48177_, new_n48178_,
    new_n48179_, new_n48180_, new_n48181_, new_n48182_, new_n48183_,
    new_n48184_, new_n48185_, new_n48186_, new_n48187_, new_n48188_,
    new_n48189_, new_n48190_, new_n48191_, new_n48192_, new_n48193_,
    new_n48194_, new_n48195_, new_n48196_, new_n48197_, new_n48198_,
    new_n48199_, new_n48200_, new_n48201_, new_n48202_, new_n48203_,
    new_n48204_, new_n48205_, new_n48206_, new_n48207_, new_n48208_,
    new_n48209_, new_n48210_, new_n48211_, new_n48212_, new_n48213_,
    new_n48214_, new_n48215_, new_n48216_, new_n48217_, new_n48218_,
    new_n48219_, new_n48220_, new_n48221_, new_n48222_, new_n48223_,
    new_n48224_, new_n48225_, new_n48226_, new_n48227_, new_n48228_,
    new_n48229_, new_n48230_, new_n48231_, new_n48232_, new_n48233_,
    new_n48234_, new_n48235_, new_n48236_, new_n48237_, new_n48238_,
    new_n48239_, new_n48240_, new_n48241_, new_n48242_, new_n48243_,
    new_n48244_, new_n48245_, new_n48246_, new_n48247_, new_n48248_,
    new_n48249_, new_n48250_, new_n48251_, new_n48252_, new_n48253_,
    new_n48254_, new_n48255_, new_n48256_, new_n48257_, new_n48258_,
    new_n48259_, new_n48260_, new_n48261_, new_n48262_, new_n48263_,
    new_n48264_, new_n48265_, new_n48266_, new_n48267_, new_n48268_,
    new_n48269_, new_n48270_, new_n48271_, new_n48272_, new_n48273_,
    new_n48274_, new_n48275_, new_n48276_, new_n48277_, new_n48278_,
    new_n48279_, new_n48280_, new_n48281_, new_n48282_, new_n48283_,
    new_n48284_, new_n48285_, new_n48286_, new_n48287_, new_n48288_,
    new_n48289_, new_n48290_, new_n48291_, new_n48292_, new_n48293_,
    new_n48294_, new_n48295_, new_n48296_, new_n48297_, new_n48298_,
    new_n48299_, new_n48300_, new_n48301_, new_n48302_, new_n48303_,
    new_n48304_, new_n48305_, new_n48306_, new_n48307_, new_n48308_,
    new_n48309_, new_n48310_, new_n48311_, new_n48312_, new_n48313_,
    new_n48314_, new_n48315_, new_n48316_, new_n48317_, new_n48318_,
    new_n48319_, new_n48320_, new_n48321_, new_n48322_, new_n48323_,
    new_n48324_, new_n48325_, new_n48326_, new_n48327_, new_n48328_,
    new_n48329_, new_n48330_, new_n48331_, new_n48332_, new_n48333_,
    new_n48334_, new_n48335_, new_n48336_, new_n48337_, new_n48338_,
    new_n48339_, new_n48340_, new_n48341_, new_n48342_, new_n48343_,
    new_n48344_, new_n48345_, new_n48346_, new_n48347_, new_n48348_,
    new_n48349_, new_n48350_, new_n48351_, new_n48352_, new_n48353_,
    new_n48354_, new_n48355_, new_n48356_, new_n48357_, new_n48358_,
    new_n48359_, new_n48360_, new_n48361_, new_n48362_, new_n48363_,
    new_n48364_, new_n48365_, new_n48366_, new_n48367_, new_n48368_,
    new_n48369_, new_n48370_, new_n48371_, new_n48372_, new_n48373_,
    new_n48374_, new_n48375_, new_n48376_, new_n48377_, new_n48378_,
    new_n48379_, new_n48380_, new_n48381_, new_n48382_, new_n48383_,
    new_n48384_, new_n48385_, new_n48386_, new_n48387_, new_n48388_,
    new_n48389_, new_n48390_, new_n48391_, new_n48392_, new_n48393_,
    new_n48394_, new_n48395_, new_n48396_, new_n48397_, new_n48398_,
    new_n48399_, new_n48400_, new_n48401_, new_n48402_, new_n48403_,
    new_n48404_, new_n48405_, new_n48406_, new_n48407_, new_n48408_,
    new_n48409_, new_n48410_, new_n48411_, new_n48412_, new_n48413_,
    new_n48414_, new_n48415_, new_n48416_, new_n48417_, new_n48418_,
    new_n48419_, new_n48420_, new_n48421_, new_n48422_, new_n48423_,
    new_n48424_, new_n48425_, new_n48426_, new_n48427_, new_n48428_,
    new_n48429_, new_n48430_, new_n48431_, new_n48432_, new_n48433_,
    new_n48434_, new_n48435_, new_n48436_, new_n48437_, new_n48438_,
    new_n48439_, new_n48440_, new_n48441_, new_n48442_, new_n48443_,
    new_n48444_, new_n48445_, new_n48446_, new_n48447_, new_n48448_,
    new_n48449_, new_n48450_, new_n48451_, new_n48452_, new_n48453_,
    new_n48454_, new_n48455_, new_n48456_, new_n48457_, new_n48458_,
    new_n48459_, new_n48460_, new_n48461_, new_n48462_, new_n48463_,
    new_n48464_, new_n48465_, new_n48466_, new_n48467_, new_n48468_,
    new_n48469_, new_n48470_, new_n48471_, new_n48472_, new_n48473_,
    new_n48474_, new_n48475_, new_n48476_, new_n48477_, new_n48478_,
    new_n48479_, new_n48480_, new_n48481_, new_n48482_, new_n48483_,
    new_n48484_, new_n48485_, new_n48486_, new_n48487_, new_n48488_,
    new_n48489_, new_n48490_, new_n48491_, new_n48492_, new_n48493_,
    new_n48494_, new_n48495_, new_n48496_, new_n48497_, new_n48498_,
    new_n48499_, new_n48500_, new_n48501_, new_n48502_, new_n48503_,
    new_n48504_, new_n48505_, new_n48506_, new_n48507_, new_n48508_,
    new_n48509_, new_n48510_, new_n48511_, new_n48512_, new_n48513_,
    new_n48514_, new_n48515_, new_n48516_, new_n48517_, new_n48518_,
    new_n48519_, new_n48520_, new_n48521_, new_n48522_, new_n48523_,
    new_n48524_, new_n48525_, new_n48526_, new_n48527_, new_n48528_,
    new_n48529_, new_n48530_, new_n48531_, new_n48532_, new_n48533_,
    new_n48534_, new_n48535_, new_n48536_, new_n48537_, new_n48538_,
    new_n48539_, new_n48540_, new_n48541_, new_n48542_, new_n48543_,
    new_n48544_, new_n48545_, new_n48546_, new_n48547_, new_n48548_,
    new_n48549_, new_n48550_, new_n48551_, new_n48552_, new_n48553_,
    new_n48554_, new_n48555_, new_n48556_, new_n48557_, new_n48558_,
    new_n48559_, new_n48560_, new_n48561_, new_n48562_, new_n48563_,
    new_n48564_, new_n48565_, new_n48566_, new_n48567_, new_n48568_,
    new_n48569_, new_n48570_, new_n48571_, new_n48572_, new_n48573_,
    new_n48574_, new_n48575_, new_n48576_, new_n48577_, new_n48578_,
    new_n48579_, new_n48580_, new_n48581_, new_n48582_, new_n48583_,
    new_n48584_, new_n48585_, new_n48586_, new_n48587_, new_n48588_,
    new_n48589_, new_n48590_, new_n48591_, new_n48592_, new_n48593_,
    new_n48594_, new_n48595_, new_n48596_, new_n48597_, new_n48598_,
    new_n48599_, new_n48600_, new_n48601_, new_n48602_, new_n48603_,
    new_n48604_, new_n48605_, new_n48606_, new_n48607_, new_n48608_,
    new_n48609_, new_n48610_, new_n48611_, new_n48612_, new_n48613_,
    new_n48614_, new_n48615_, new_n48616_, new_n48617_, new_n48618_,
    new_n48619_, new_n48620_, new_n48621_, new_n48622_, new_n48623_,
    new_n48624_, new_n48625_, new_n48626_, new_n48627_, new_n48628_,
    new_n48629_, new_n48630_, new_n48631_, new_n48632_, new_n48633_,
    new_n48634_, new_n48635_, new_n48636_, new_n48637_, new_n48638_,
    new_n48639_, new_n48640_, new_n48641_, new_n48642_, new_n48643_,
    new_n48644_, new_n48645_, new_n48646_, new_n48647_, new_n48648_,
    new_n48649_, new_n48650_, new_n48651_, new_n48652_, new_n48653_,
    new_n48654_, new_n48655_, new_n48656_, new_n48657_, new_n48658_,
    new_n48659_, new_n48660_, new_n48661_, new_n48662_, new_n48663_,
    new_n48664_, new_n48665_, new_n48666_, new_n48667_, new_n48668_,
    new_n48669_, new_n48670_, new_n48671_, new_n48672_, new_n48673_,
    new_n48674_, new_n48675_, new_n48676_, new_n48677_, new_n48678_,
    new_n48679_, new_n48680_, new_n48681_, new_n48682_, new_n48683_,
    new_n48684_, new_n48685_, new_n48686_, new_n48687_, new_n48688_,
    new_n48689_, new_n48690_, new_n48691_, new_n48692_, new_n48693_,
    new_n48694_, new_n48695_, new_n48696_, new_n48697_, new_n48698_,
    new_n48699_, new_n48700_, new_n48701_, new_n48702_, new_n48703_,
    new_n48704_, new_n48705_, new_n48706_, new_n48707_, new_n48708_,
    new_n48709_, new_n48710_, new_n48711_, new_n48712_, new_n48713_,
    new_n48714_, new_n48715_, new_n48716_, new_n48717_, new_n48718_,
    new_n48719_, new_n48720_, new_n48721_, new_n48722_, new_n48723_,
    new_n48724_, new_n48725_, new_n48726_, new_n48727_, new_n48728_,
    new_n48729_, new_n48730_, new_n48731_, new_n48732_, new_n48733_,
    new_n48734_, new_n48735_, new_n48736_, new_n48737_, new_n48738_,
    new_n48739_, new_n48740_, new_n48741_, new_n48742_, new_n48743_,
    new_n48744_, new_n48745_, new_n48746_, new_n48747_, new_n48748_,
    new_n48749_, new_n48750_, new_n48751_, new_n48752_, new_n48753_,
    new_n48754_, new_n48755_, new_n48756_, new_n48757_, new_n48758_,
    new_n48759_, new_n48760_, new_n48761_, new_n48762_, new_n48763_,
    new_n48764_, new_n48765_, new_n48766_, new_n48767_, new_n48768_,
    new_n48769_, new_n48770_, new_n48771_, new_n48772_, new_n48773_,
    new_n48774_, new_n48775_, new_n48776_, new_n48777_, new_n48778_,
    new_n48779_, new_n48780_, new_n48781_, new_n48782_, new_n48783_,
    new_n48784_, new_n48785_, new_n48786_, new_n48787_, new_n48788_,
    new_n48789_, new_n48790_, new_n48791_, new_n48792_, new_n48793_,
    new_n48794_, new_n48795_, new_n48796_, new_n48797_, new_n48798_,
    new_n48799_, new_n48800_, new_n48801_, new_n48802_, new_n48803_,
    new_n48804_, new_n48805_, new_n48806_, new_n48807_, new_n48808_,
    new_n48809_, new_n48810_, new_n48811_, new_n48812_, new_n48813_,
    new_n48814_, new_n48815_, new_n48816_, new_n48817_, new_n48818_,
    new_n48819_, new_n48820_, new_n48821_, new_n48822_, new_n48823_,
    new_n48824_, new_n48825_, new_n48826_, new_n48827_, new_n48828_,
    new_n48829_, new_n48830_, new_n48831_, new_n48832_, new_n48833_,
    new_n48834_, new_n48835_, new_n48836_, new_n48837_, new_n48838_,
    new_n48839_, new_n48840_, new_n48841_, new_n48842_, new_n48843_,
    new_n48844_, new_n48845_, new_n48846_, new_n48847_, new_n48848_,
    new_n48849_, new_n48850_, new_n48851_, new_n48852_, new_n48853_,
    new_n48854_, new_n48855_, new_n48856_, new_n48857_, new_n48858_,
    new_n48859_, new_n48860_, new_n48861_, new_n48862_, new_n48863_,
    new_n48864_, new_n48865_, new_n48866_, new_n48867_, new_n48868_,
    new_n48869_, new_n48870_, new_n48871_, new_n48872_, new_n48873_,
    new_n48874_, new_n48875_, new_n48876_, new_n48877_, new_n48878_,
    new_n48879_, new_n48880_, new_n48881_, new_n48882_, new_n48883_,
    new_n48884_, new_n48885_, new_n48886_, new_n48887_, new_n48888_,
    new_n48889_, new_n48890_, new_n48891_, new_n48892_, new_n48893_,
    new_n48894_, new_n48895_, new_n48896_, new_n48897_, new_n48898_,
    new_n48899_, new_n48900_, new_n48901_, new_n48902_, new_n48903_,
    new_n48904_, new_n48905_, new_n48906_, new_n48907_, new_n48908_,
    new_n48909_, new_n48910_, new_n48911_, new_n48912_, new_n48913_,
    new_n48914_, new_n48915_, new_n48916_, new_n48917_, new_n48918_,
    new_n48919_, new_n48920_, new_n48921_, new_n48922_, new_n48923_,
    new_n48924_, new_n48925_, new_n48926_, new_n48927_, new_n48928_,
    new_n48929_, new_n48930_, new_n48931_, new_n48932_, new_n48933_,
    new_n48934_, new_n48935_, new_n48936_, new_n48937_, new_n48938_,
    new_n48939_, new_n48940_, new_n48941_, new_n48942_, new_n48943_,
    new_n48944_, new_n48945_, new_n48946_, new_n48947_, new_n48948_,
    new_n48949_, new_n48950_, new_n48951_, new_n48952_, new_n48953_,
    new_n48954_, new_n48955_, new_n48956_, new_n48957_, new_n48958_,
    new_n48959_, new_n48960_, new_n48961_, new_n48962_, new_n48963_,
    new_n48964_, new_n48965_, new_n48966_, new_n48967_, new_n48968_,
    new_n48969_, new_n48970_, new_n48971_, new_n48972_, new_n48973_,
    new_n48974_, new_n48975_, new_n48976_, new_n48977_, new_n48978_,
    new_n48979_, new_n48980_, new_n48981_, new_n48982_, new_n48983_,
    new_n48984_, new_n48985_, new_n48986_, new_n48987_, new_n48988_,
    new_n48989_, new_n48990_, new_n48991_, new_n48992_, new_n48993_,
    new_n48994_, new_n48995_, new_n48996_, new_n48997_, new_n48998_,
    new_n48999_, new_n49000_, new_n49001_, new_n49002_, new_n49003_,
    new_n49004_, new_n49005_, new_n49006_, new_n49007_, new_n49008_,
    new_n49009_, new_n49010_, new_n49011_, new_n49012_, new_n49013_,
    new_n49014_, new_n49015_, new_n49016_, new_n49017_, new_n49018_,
    new_n49019_, new_n49020_, new_n49021_, new_n49022_, new_n49023_,
    new_n49024_, new_n49025_, new_n49026_, new_n49027_, new_n49028_,
    new_n49029_, new_n49030_, new_n49031_, new_n49032_, new_n49033_,
    new_n49034_, new_n49035_, new_n49036_, new_n49037_, new_n49038_,
    new_n49039_, new_n49040_, new_n49041_, new_n49042_, new_n49043_,
    new_n49044_, new_n49045_, new_n49046_, new_n49047_, new_n49048_,
    new_n49049_, new_n49050_, new_n49051_, new_n49052_, new_n49053_,
    new_n49054_, new_n49055_, new_n49056_, new_n49057_, new_n49058_,
    new_n49059_, new_n49060_, new_n49061_, new_n49062_, new_n49063_,
    new_n49064_, new_n49065_, new_n49066_, new_n49067_, new_n49068_,
    new_n49069_, new_n49070_, new_n49071_, new_n49072_, new_n49073_,
    new_n49074_, new_n49075_, new_n49076_, new_n49077_, new_n49078_,
    new_n49079_, new_n49080_, new_n49081_, new_n49082_, new_n49083_,
    new_n49084_, new_n49085_, new_n49086_, new_n49087_, new_n49088_,
    new_n49089_, new_n49090_, new_n49091_, new_n49092_, new_n49093_,
    new_n49094_, new_n49095_, new_n49096_, new_n49097_, new_n49098_,
    new_n49099_, new_n49100_, new_n49101_, new_n49102_, new_n49103_,
    new_n49104_, new_n49105_, new_n49106_, new_n49107_, new_n49108_,
    new_n49109_, new_n49110_, new_n49111_, new_n49112_, new_n49113_,
    new_n49114_, new_n49115_, new_n49116_, new_n49117_, new_n49118_,
    new_n49119_, new_n49120_, new_n49121_, new_n49122_, new_n49123_,
    new_n49124_, new_n49125_, new_n49126_, new_n49127_, new_n49128_,
    new_n49129_, new_n49130_, new_n49131_, new_n49132_, new_n49133_,
    new_n49134_, new_n49135_, new_n49136_, new_n49137_, new_n49138_,
    new_n49139_, new_n49140_, new_n49141_, new_n49142_, new_n49143_,
    new_n49144_, new_n49145_, new_n49146_, new_n49147_, new_n49148_,
    new_n49149_, new_n49150_, new_n49151_, new_n49152_, new_n49153_,
    new_n49154_, new_n49155_, new_n49156_, new_n49157_, new_n49158_,
    new_n49159_, new_n49160_, new_n49161_, new_n49162_, new_n49163_,
    new_n49164_, new_n49165_, new_n49166_, new_n49167_, new_n49168_,
    new_n49169_, new_n49170_, new_n49171_, new_n49172_, new_n49173_,
    new_n49174_, new_n49175_, new_n49176_, new_n49177_, new_n49178_,
    new_n49179_, new_n49180_, new_n49181_, new_n49182_, new_n49183_,
    new_n49184_, new_n49185_, new_n49186_, new_n49187_, new_n49188_,
    new_n49189_, new_n49190_, new_n49191_, new_n49192_, new_n49193_,
    new_n49194_, new_n49195_, new_n49196_, new_n49197_, new_n49198_,
    new_n49199_, new_n49200_, new_n49201_, new_n49202_, new_n49203_,
    new_n49204_, new_n49205_, new_n49206_, new_n49207_, new_n49208_,
    new_n49209_, new_n49210_, new_n49211_, new_n49212_, new_n49213_,
    new_n49214_, new_n49215_, new_n49216_, new_n49217_, new_n49218_,
    new_n49219_, new_n49220_, new_n49221_, new_n49222_, new_n49223_,
    new_n49224_, new_n49225_, new_n49226_, new_n49227_, new_n49228_,
    new_n49229_, new_n49230_, new_n49231_, new_n49232_, new_n49233_,
    new_n49234_, new_n49235_, new_n49236_, new_n49237_, new_n49238_,
    new_n49239_, new_n49240_, new_n49241_, new_n49242_, new_n49243_,
    new_n49244_, new_n49245_, new_n49246_, new_n49247_, new_n49248_,
    new_n49249_, new_n49250_, new_n49251_, new_n49252_, new_n49253_,
    new_n49254_, new_n49255_, new_n49256_, new_n49257_, new_n49258_,
    new_n49259_, new_n49260_, new_n49261_, new_n49262_, new_n49263_,
    new_n49264_, new_n49265_, new_n49266_, new_n49267_, new_n49268_,
    new_n49269_, new_n49270_, new_n49271_, new_n49272_, new_n49273_,
    new_n49274_, new_n49275_, new_n49276_, new_n49277_, new_n49278_,
    new_n49279_, new_n49280_, new_n49281_, new_n49282_, new_n49283_,
    new_n49284_, new_n49285_, new_n49286_, new_n49287_, new_n49288_,
    new_n49289_, new_n49290_, new_n49291_, new_n49292_, new_n49293_,
    new_n49294_, new_n49295_, new_n49296_, new_n49297_, new_n49298_,
    new_n49299_, new_n49300_, new_n49301_, new_n49302_, new_n49303_,
    new_n49304_, new_n49305_, new_n49306_, new_n49307_, new_n49308_,
    new_n49309_, new_n49310_, new_n49311_, new_n49312_, new_n49313_,
    new_n49314_, new_n49315_, new_n49316_, new_n49317_, new_n49318_,
    new_n49319_, new_n49320_, new_n49321_, new_n49322_, new_n49323_,
    new_n49324_, new_n49325_, new_n49326_, new_n49327_, new_n49328_,
    new_n49329_, new_n49330_, new_n49331_, new_n49332_, new_n49333_,
    new_n49334_, new_n49335_, new_n49336_, new_n49337_, new_n49338_,
    new_n49339_, new_n49340_, new_n49341_, new_n49342_, new_n49343_,
    new_n49344_, new_n49345_, new_n49346_, new_n49347_, new_n49348_,
    new_n49349_, new_n49350_, new_n49351_, new_n49352_, new_n49353_,
    new_n49354_, new_n49355_, new_n49356_, new_n49357_, new_n49358_,
    new_n49359_, new_n49360_, new_n49361_, new_n49362_, new_n49363_,
    new_n49364_, new_n49365_, new_n49366_, new_n49367_, new_n49368_,
    new_n49369_, new_n49370_, new_n49371_, new_n49372_, new_n49373_,
    new_n49374_, new_n49375_, new_n49376_, new_n49377_, new_n49378_,
    new_n49379_, new_n49380_, new_n49381_, new_n49382_, new_n49383_,
    new_n49384_, new_n49385_, new_n49386_, new_n49387_, new_n49388_,
    new_n49389_, new_n49390_, new_n49391_, new_n49392_, new_n49393_,
    new_n49394_, new_n49395_, new_n49396_, new_n49397_, new_n49398_,
    new_n49399_, new_n49400_, new_n49401_, new_n49402_, new_n49403_,
    new_n49404_, new_n49405_, new_n49406_, new_n49407_, new_n49408_,
    new_n49409_, new_n49410_, new_n49411_, new_n49412_, new_n49413_,
    new_n49414_, new_n49415_, new_n49416_, new_n49417_, new_n49418_,
    new_n49419_, new_n49420_, new_n49421_, new_n49422_, new_n49423_,
    new_n49424_, new_n49425_, new_n49426_, new_n49427_, new_n49428_,
    new_n49429_, new_n49430_, new_n49431_, new_n49432_, new_n49433_,
    new_n49434_, new_n49435_, new_n49436_, new_n49437_, new_n49438_,
    new_n49439_, new_n49440_, new_n49441_, new_n49442_, new_n49443_,
    new_n49444_, new_n49445_, new_n49446_, new_n49447_, new_n49448_,
    new_n49449_, new_n49450_, new_n49451_, new_n49452_, new_n49453_,
    new_n49454_, new_n49455_, new_n49456_, new_n49457_, new_n49458_,
    new_n49459_, new_n49460_, new_n49461_, new_n49462_, new_n49463_,
    new_n49464_, new_n49465_, new_n49466_, new_n49467_, new_n49468_,
    new_n49469_, new_n49470_, new_n49471_, new_n49472_, new_n49473_,
    new_n49474_, new_n49475_, new_n49476_, new_n49477_, new_n49478_,
    new_n49479_, new_n49480_, new_n49481_, new_n49482_, new_n49483_,
    new_n49484_, new_n49485_, new_n49486_, new_n49487_, new_n49488_,
    new_n49489_, new_n49490_, new_n49491_, new_n49492_, new_n49493_,
    new_n49494_, new_n49495_, new_n49496_, new_n49497_, new_n49498_,
    new_n49499_, new_n49500_, new_n49501_, new_n49502_, new_n49503_,
    new_n49504_, new_n49505_, new_n49506_, new_n49507_, new_n49508_,
    new_n49509_, new_n49510_, new_n49511_, new_n49512_, new_n49513_,
    new_n49514_, new_n49515_, new_n49516_, new_n49517_, new_n49518_,
    new_n49519_, new_n49520_, new_n49521_, new_n49522_, new_n49523_,
    new_n49524_, new_n49525_, new_n49526_, new_n49527_, new_n49528_,
    new_n49529_, new_n49530_, new_n49531_, new_n49532_, new_n49533_,
    new_n49534_, new_n49535_, new_n49536_, new_n49537_, new_n49538_,
    new_n49539_, new_n49540_, new_n49541_, new_n49542_, new_n49543_,
    new_n49544_, new_n49545_, new_n49546_, new_n49547_, new_n49548_,
    new_n49549_, new_n49550_, new_n49551_, new_n49552_, new_n49553_,
    new_n49554_, new_n49555_, new_n49556_, new_n49557_, new_n49558_,
    new_n49559_, new_n49560_, new_n49561_, new_n49562_, new_n49563_,
    new_n49564_, new_n49565_, new_n49566_, new_n49567_, new_n49568_,
    new_n49569_, new_n49570_, new_n49571_, new_n49572_, new_n49573_,
    new_n49574_, new_n49575_, new_n49576_, new_n49577_, new_n49578_,
    new_n49579_, new_n49580_, new_n49581_, new_n49582_, new_n49583_,
    new_n49584_, new_n49585_, new_n49586_, new_n49587_, new_n49588_,
    new_n49589_, new_n49590_, new_n49591_, new_n49592_, new_n49593_,
    new_n49594_, new_n49595_, new_n49596_, new_n49597_, new_n49598_,
    new_n49599_, new_n49600_, new_n49601_, new_n49602_, new_n49603_,
    new_n49604_, new_n49605_, new_n49606_, new_n49607_, new_n49608_,
    new_n49609_, new_n49610_, new_n49611_, new_n49612_, new_n49613_,
    new_n49614_, new_n49615_, new_n49616_, new_n49617_, new_n49618_,
    new_n49619_, new_n49620_, new_n49621_, new_n49622_, new_n49623_,
    new_n49624_, new_n49625_, new_n49626_, new_n49627_, new_n49628_,
    new_n49629_, new_n49630_, new_n49631_, new_n49632_, new_n49633_,
    new_n49634_, new_n49635_, new_n49636_, new_n49637_, new_n49638_,
    new_n49639_, new_n49640_, new_n49641_, new_n49642_, new_n49643_,
    new_n49644_, new_n49645_, new_n49646_, new_n49647_, new_n49648_,
    new_n49649_, new_n49650_, new_n49651_, new_n49652_, new_n49653_,
    new_n49654_, new_n49655_, new_n49656_, new_n49657_, new_n49658_,
    new_n49659_, new_n49660_, new_n49661_, new_n49662_, new_n49663_,
    new_n49664_, new_n49665_, new_n49666_, new_n49667_, new_n49668_,
    new_n49669_, new_n49670_, new_n49671_, new_n49672_, new_n49673_,
    new_n49674_, new_n49675_, new_n49676_, new_n49677_, new_n49678_,
    new_n49679_, new_n49680_, new_n49681_, new_n49682_, new_n49683_,
    new_n49684_, new_n49685_, new_n49686_, new_n49687_, new_n49688_,
    new_n49689_, new_n49690_, new_n49691_, new_n49692_, new_n49693_,
    new_n49694_, new_n49695_, new_n49696_, new_n49697_, new_n49698_,
    new_n49699_, new_n49700_, new_n49701_, new_n49702_, new_n49703_,
    new_n49704_, new_n49705_, new_n49706_, new_n49707_, new_n49708_,
    new_n49709_, new_n49710_, new_n49711_, new_n49712_, new_n49713_,
    new_n49714_, new_n49715_, new_n49716_, new_n49717_, new_n49718_,
    new_n49719_, new_n49720_, new_n49721_, new_n49722_, new_n49723_,
    new_n49724_, new_n49725_, new_n49726_, new_n49727_, new_n49728_,
    new_n49729_, new_n49730_, new_n49731_, new_n49732_, new_n49733_,
    new_n49734_, new_n49735_, new_n49736_, new_n49737_, new_n49738_,
    new_n49739_, new_n49740_, new_n49741_, new_n49742_, new_n49743_,
    new_n49744_, new_n49745_, new_n49746_, new_n49747_, new_n49748_,
    new_n49749_, new_n49750_, new_n49751_, new_n49752_, new_n49753_,
    new_n49754_, new_n49755_, new_n49756_, new_n49757_, new_n49758_,
    new_n49759_, new_n49760_, new_n49761_, new_n49762_, new_n49763_,
    new_n49764_, new_n49765_, new_n49766_, new_n49767_, new_n49768_,
    new_n49769_, new_n49770_, new_n49771_, new_n49772_, new_n49773_,
    new_n49774_, new_n49775_, new_n49776_, new_n49777_, new_n49778_,
    new_n49779_, new_n49780_, new_n49781_, new_n49782_, new_n49783_,
    new_n49784_, new_n49785_, new_n49786_, new_n49787_, new_n49788_,
    new_n49789_, new_n49790_, new_n49791_, new_n49792_, new_n49793_,
    new_n49794_, new_n49795_, new_n49796_, new_n49797_, new_n49798_,
    new_n49799_, new_n49800_, new_n49801_, new_n49802_, new_n49803_,
    new_n49804_, new_n49805_, new_n49806_, new_n49807_, new_n49808_,
    new_n49809_, new_n49810_, new_n49811_, new_n49812_, new_n49813_,
    new_n49814_, new_n49815_, new_n49816_, new_n49817_, new_n49818_,
    new_n49819_, new_n49820_, new_n49821_, new_n49822_, new_n49823_,
    new_n49824_, new_n49825_, new_n49826_, new_n49827_, new_n49828_,
    new_n49829_, new_n49830_, new_n49831_, new_n49832_, new_n49833_,
    new_n49834_, new_n49835_, new_n49836_, new_n49837_, new_n49838_,
    new_n49839_, new_n49840_, new_n49841_, new_n49842_, new_n49843_,
    new_n49844_, new_n49845_, new_n49846_, new_n49847_, new_n49848_,
    new_n49849_, new_n49850_, new_n49851_, new_n49852_, new_n49853_,
    new_n49854_, new_n49855_, new_n49856_, new_n49857_, new_n49858_,
    new_n49859_, new_n49860_, new_n49861_, new_n49862_, new_n49863_,
    new_n49864_, new_n49865_, new_n49866_, new_n49867_, new_n49868_,
    new_n49869_, new_n49870_, new_n49871_, new_n49872_, new_n49873_,
    new_n49874_, new_n49875_, new_n49876_, new_n49877_, new_n49878_,
    new_n49879_, new_n49880_, new_n49881_, new_n49882_, new_n49883_,
    new_n49884_, new_n49885_, new_n49886_, new_n49887_, new_n49888_,
    new_n49889_, new_n49890_, new_n49891_, new_n49892_, new_n49893_,
    new_n49894_, new_n49895_, new_n49896_, new_n49897_, new_n49898_,
    new_n49899_, new_n49900_, new_n49901_, new_n49902_, new_n49903_,
    new_n49904_, new_n49905_, new_n49906_, new_n49907_, new_n49908_,
    new_n49909_, new_n49910_, new_n49911_, new_n49912_, new_n49913_,
    new_n49914_, new_n49915_, new_n49916_, new_n49917_, new_n49918_,
    new_n49919_, new_n49920_, new_n49921_, new_n49922_, new_n49923_,
    new_n49924_, new_n49925_, new_n49926_, new_n49927_, new_n49928_,
    new_n49929_, new_n49930_, new_n49931_, new_n49932_, new_n49933_,
    new_n49934_, new_n49935_, new_n49936_, new_n49937_, new_n49938_,
    new_n49939_, new_n49940_, new_n49941_, new_n49942_, new_n49943_,
    new_n49944_, new_n49945_, new_n49946_, new_n49947_, new_n49948_,
    new_n49949_, new_n49950_, new_n49951_, new_n49952_, new_n49953_,
    new_n49954_, new_n49955_, new_n49956_, new_n49957_, new_n49958_,
    new_n49959_, new_n49960_, new_n49961_, new_n49962_, new_n49963_,
    new_n49964_, new_n49965_, new_n49966_, new_n49967_, new_n49968_,
    new_n49969_, new_n49970_, new_n49971_, new_n49972_, new_n49973_,
    new_n49974_, new_n49975_, new_n49976_, new_n49977_, new_n49978_,
    new_n49979_, new_n49980_, new_n49981_, new_n49982_, new_n49983_,
    new_n49984_, new_n49985_, new_n49986_, new_n49987_, new_n49988_,
    new_n49989_, new_n49990_, new_n49991_, new_n49992_, new_n49993_,
    new_n49994_, new_n49995_, new_n49996_, new_n49997_, new_n49998_,
    new_n49999_, new_n50000_, new_n50001_, new_n50002_, new_n50003_,
    new_n50004_, new_n50005_, new_n50006_, new_n50007_, new_n50008_,
    new_n50009_, new_n50010_, new_n50011_, new_n50012_, new_n50013_,
    new_n50014_, new_n50015_, new_n50016_, new_n50017_, new_n50018_,
    new_n50019_, new_n50020_, new_n50021_, new_n50022_, new_n50023_,
    new_n50024_, new_n50025_, new_n50026_, new_n50027_, new_n50028_,
    new_n50029_, new_n50030_, new_n50031_, new_n50032_, new_n50033_,
    new_n50034_, new_n50035_, new_n50036_, new_n50037_, new_n50038_,
    new_n50039_, new_n50040_, new_n50041_, new_n50042_, new_n50043_,
    new_n50044_, new_n50045_, new_n50046_, new_n50047_, new_n50048_,
    new_n50049_, new_n50050_, new_n50051_, new_n50052_, new_n50053_,
    new_n50054_, new_n50055_, new_n50056_, new_n50057_, new_n50058_,
    new_n50059_, new_n50060_, new_n50061_, new_n50062_, new_n50063_,
    new_n50064_, new_n50065_, new_n50066_, new_n50067_, new_n50068_,
    new_n50069_, new_n50070_, new_n50071_, new_n50072_, new_n50073_,
    new_n50074_, new_n50075_, new_n50076_, new_n50077_, new_n50078_,
    new_n50079_, new_n50080_, new_n50081_, new_n50082_, new_n50083_,
    new_n50084_, new_n50085_, new_n50086_, new_n50087_, new_n50088_,
    new_n50089_, new_n50090_, new_n50091_, new_n50092_, new_n50093_,
    new_n50094_, new_n50095_, new_n50096_, new_n50097_, new_n50098_,
    new_n50099_, new_n50100_, new_n50101_, new_n50102_, new_n50103_,
    new_n50104_, new_n50105_, new_n50106_, new_n50107_, new_n50108_,
    new_n50109_, new_n50110_, new_n50111_, new_n50112_, new_n50113_,
    new_n50114_, new_n50115_, new_n50116_, new_n50117_, new_n50118_,
    new_n50119_, new_n50120_, new_n50121_, new_n50122_, new_n50123_,
    new_n50124_, new_n50125_, new_n50126_, new_n50127_, new_n50128_,
    new_n50129_, new_n50130_, new_n50131_, new_n50132_, new_n50133_,
    new_n50134_, new_n50135_, new_n50136_, new_n50137_, new_n50138_,
    new_n50139_, new_n50140_, new_n50141_, new_n50142_, new_n50143_,
    new_n50144_, new_n50145_, new_n50146_, new_n50147_, new_n50148_,
    new_n50149_, new_n50150_, new_n50151_, new_n50152_, new_n50153_,
    new_n50154_, new_n50155_, new_n50156_, new_n50157_, new_n50158_,
    new_n50159_, new_n50160_, new_n50161_, new_n50162_, new_n50163_,
    new_n50164_, new_n50165_, new_n50166_, new_n50167_, new_n50168_,
    new_n50169_, new_n50170_, new_n50171_, new_n50172_, new_n50173_,
    new_n50174_, new_n50175_, new_n50176_, new_n50177_, new_n50178_,
    new_n50179_, new_n50180_, new_n50181_, new_n50182_, new_n50183_,
    new_n50184_, new_n50185_, new_n50186_, new_n50187_, new_n50188_,
    new_n50189_, new_n50190_, new_n50191_, new_n50192_, new_n50193_,
    new_n50194_, new_n50195_, new_n50196_, new_n50197_, new_n50198_,
    new_n50199_, new_n50200_, new_n50201_, new_n50202_, new_n50203_,
    new_n50204_, new_n50205_, new_n50206_, new_n50207_, new_n50208_,
    new_n50209_, new_n50210_, new_n50211_, new_n50212_, new_n50213_,
    new_n50214_, new_n50215_, new_n50216_, new_n50217_, new_n50218_,
    new_n50219_, new_n50220_, new_n50221_, new_n50222_, new_n50223_,
    new_n50224_, new_n50225_, new_n50226_, new_n50227_, new_n50228_,
    new_n50229_, new_n50230_, new_n50231_, new_n50232_, new_n50233_,
    new_n50234_, new_n50235_, new_n50236_, new_n50237_, new_n50238_,
    new_n50239_, new_n50240_, new_n50241_, new_n50242_, new_n50243_,
    new_n50244_, new_n50245_, new_n50246_, new_n50247_, new_n50248_,
    new_n50249_, new_n50250_, new_n50251_, new_n50252_, new_n50253_,
    new_n50254_, new_n50255_, new_n50256_, new_n50257_, new_n50258_,
    new_n50259_, new_n50260_, new_n50261_, new_n50262_, new_n50263_,
    new_n50264_, new_n50265_, new_n50266_, new_n50267_, new_n50268_,
    new_n50269_, new_n50270_, new_n50271_, new_n50272_, new_n50273_,
    new_n50274_, new_n50275_, new_n50276_, new_n50277_, new_n50278_,
    new_n50279_, new_n50280_, new_n50281_, new_n50282_, new_n50283_,
    new_n50284_, new_n50285_, new_n50286_, new_n50287_, new_n50288_,
    new_n50289_, new_n50290_, new_n50291_, new_n50292_, new_n50293_,
    new_n50294_, new_n50295_, new_n50296_, new_n50297_, new_n50298_,
    new_n50299_, new_n50300_, new_n50301_, new_n50302_, new_n50303_,
    new_n50304_, new_n50305_, new_n50306_, new_n50307_, new_n50308_,
    new_n50309_, new_n50310_, new_n50311_, new_n50312_, new_n50313_,
    new_n50314_, new_n50315_, new_n50316_, new_n50317_, new_n50318_,
    new_n50319_, new_n50320_, new_n50321_, new_n50322_, new_n50323_,
    new_n50324_, new_n50325_, new_n50326_, new_n50327_, new_n50328_,
    new_n50329_, new_n50330_, new_n50331_, new_n50332_, new_n50333_,
    new_n50334_, new_n50335_, new_n50336_, new_n50337_, new_n50338_,
    new_n50339_, new_n50340_, new_n50341_, new_n50342_, new_n50343_,
    new_n50344_, new_n50345_, new_n50346_, new_n50347_, new_n50348_,
    new_n50349_, new_n50350_, new_n50351_, new_n50352_, new_n50353_,
    new_n50354_, new_n50355_, new_n50356_, new_n50357_, new_n50358_,
    new_n50359_, new_n50360_, new_n50361_, new_n50362_, new_n50363_,
    new_n50364_, new_n50365_, new_n50366_, new_n50367_, new_n50368_,
    new_n50369_, new_n50370_, new_n50371_, new_n50372_, new_n50373_,
    new_n50374_, new_n50375_, new_n50376_, new_n50377_, new_n50378_,
    new_n50379_, new_n50380_, new_n50381_, new_n50382_, new_n50383_,
    new_n50384_, new_n50385_, new_n50386_, new_n50387_, new_n50388_,
    new_n50389_, new_n50390_, new_n50391_, new_n50392_, new_n50393_,
    new_n50394_, new_n50395_, new_n50396_, new_n50397_, new_n50398_,
    new_n50399_, new_n50400_, new_n50401_, new_n50402_, new_n50403_,
    new_n50404_, new_n50405_, new_n50406_, new_n50407_, new_n50408_,
    new_n50409_, new_n50410_, new_n50411_, new_n50412_, new_n50413_,
    new_n50414_, new_n50415_, new_n50416_, new_n50417_, new_n50418_,
    new_n50419_, new_n50420_, new_n50421_, new_n50422_, new_n50423_,
    new_n50424_, new_n50425_, new_n50426_, new_n50427_, new_n50428_,
    new_n50429_, new_n50430_, new_n50431_, new_n50432_, new_n50433_,
    new_n50434_, new_n50435_, new_n50436_, new_n50437_, new_n50438_,
    new_n50439_, new_n50440_, new_n50441_, new_n50442_, new_n50443_,
    new_n50444_, new_n50445_, new_n50446_, new_n50447_, new_n50448_,
    new_n50449_, new_n50450_, new_n50451_, new_n50452_, new_n50453_,
    new_n50454_, new_n50455_, new_n50456_, new_n50457_, new_n50458_,
    new_n50459_, new_n50460_, new_n50461_, new_n50462_, new_n50463_,
    new_n50464_, new_n50465_, new_n50466_, new_n50467_, new_n50468_,
    new_n50469_, new_n50470_, new_n50471_, new_n50472_, new_n50473_,
    new_n50474_, new_n50475_, new_n50476_, new_n50477_, new_n50478_,
    new_n50479_, new_n50480_, new_n50481_, new_n50482_, new_n50483_,
    new_n50484_, new_n50485_, new_n50486_, new_n50487_, new_n50488_,
    new_n50489_, new_n50490_, new_n50491_, new_n50492_, new_n50493_,
    new_n50494_, new_n50495_, new_n50496_, new_n50497_, new_n50498_,
    new_n50499_, new_n50500_, new_n50501_, new_n50502_, new_n50503_,
    new_n50504_, new_n50505_, new_n50506_, new_n50507_, new_n50508_,
    new_n50509_, new_n50510_, new_n50511_, new_n50512_, new_n50513_,
    new_n50514_, new_n50515_, new_n50516_, new_n50517_, new_n50518_,
    new_n50519_, new_n50520_, new_n50521_, new_n50522_, new_n50523_,
    new_n50524_, new_n50525_, new_n50526_, new_n50527_, new_n50528_,
    new_n50529_, new_n50530_, new_n50531_, new_n50532_, new_n50533_,
    new_n50534_, new_n50535_, new_n50536_, new_n50537_, new_n50538_,
    new_n50539_, new_n50540_, new_n50541_, new_n50542_, new_n50543_,
    new_n50544_, new_n50545_, new_n50546_, new_n50547_, new_n50548_,
    new_n50549_, new_n50550_, new_n50551_, new_n50552_, new_n50553_,
    new_n50554_, new_n50555_, new_n50556_, new_n50557_, new_n50558_,
    new_n50559_, new_n50560_, new_n50561_, new_n50562_, new_n50563_,
    new_n50564_, new_n50565_, new_n50566_, new_n50567_, new_n50568_,
    new_n50569_, new_n50570_, new_n50571_, new_n50572_, new_n50573_,
    new_n50574_, new_n50575_, new_n50576_, new_n50577_, new_n50578_,
    new_n50579_, new_n50580_, new_n50581_, new_n50582_, new_n50583_,
    new_n50584_, new_n50585_, new_n50586_, new_n50587_, new_n50588_,
    new_n50589_, new_n50590_, new_n50591_, new_n50592_, new_n50593_,
    new_n50594_, new_n50595_, new_n50596_, new_n50597_, new_n50598_,
    new_n50599_, new_n50600_, new_n50601_, new_n50602_, new_n50603_,
    new_n50604_, new_n50605_, new_n50606_, new_n50607_, new_n50608_,
    new_n50609_, new_n50610_, new_n50611_, new_n50612_, new_n50613_,
    new_n50614_, new_n50615_, new_n50616_, new_n50617_, new_n50618_,
    new_n50619_, new_n50620_, new_n50621_, new_n50622_, new_n50623_,
    new_n50624_, new_n50625_, new_n50626_, new_n50627_, new_n50628_,
    new_n50629_, new_n50630_, new_n50631_, new_n50632_, new_n50633_,
    new_n50634_, new_n50635_, new_n50636_, new_n50637_, new_n50638_,
    new_n50639_, new_n50640_, new_n50641_, new_n50642_, new_n50643_,
    new_n50644_, new_n50645_, new_n50646_, new_n50647_, new_n50648_,
    new_n50649_, new_n50650_, new_n50651_, new_n50652_, new_n50653_,
    new_n50654_, new_n50655_, new_n50656_, new_n50657_, new_n50658_,
    new_n50659_, new_n50660_, new_n50661_, new_n50662_, new_n50663_,
    new_n50664_, new_n50665_, new_n50666_, new_n50667_, new_n50668_,
    new_n50669_, new_n50670_, new_n50671_, new_n50672_, new_n50673_,
    new_n50674_, new_n50675_, new_n50676_, new_n50677_, new_n50678_,
    new_n50679_, new_n50680_, new_n50681_, new_n50682_, new_n50683_,
    new_n50684_, new_n50685_, new_n50686_, new_n50687_, new_n50688_,
    new_n50689_, new_n50690_, new_n50691_, new_n50692_, new_n50693_,
    new_n50694_, new_n50695_, new_n50696_, new_n50697_, new_n50698_,
    new_n50699_, new_n50700_, new_n50701_, new_n50702_, new_n50703_,
    new_n50704_, new_n50705_, new_n50706_, new_n50707_, new_n50708_,
    new_n50709_, new_n50710_, new_n50711_, new_n50712_, new_n50713_,
    new_n50714_, new_n50715_, new_n50716_, new_n50717_, new_n50718_,
    new_n50719_, new_n50720_, new_n50721_, new_n50722_, new_n50723_,
    new_n50724_, new_n50725_, new_n50726_, new_n50727_, new_n50728_,
    new_n50729_, new_n50730_, new_n50731_, new_n50732_, new_n50733_,
    new_n50734_, new_n50735_, new_n50736_, new_n50737_, new_n50738_,
    new_n50739_, new_n50740_, new_n50741_, new_n50742_, new_n50743_,
    new_n50744_, new_n50745_, new_n50746_, new_n50747_, new_n50748_,
    new_n50749_, new_n50750_, new_n50751_, new_n50752_, new_n50753_,
    new_n50754_, new_n50755_, new_n50756_, new_n50757_, new_n50758_,
    new_n50759_, new_n50760_, new_n50761_, new_n50762_, new_n50763_,
    new_n50764_, new_n50765_, new_n50766_, new_n50767_, new_n50768_,
    new_n50769_, new_n50770_, new_n50771_, new_n50772_, new_n50773_,
    new_n50774_, new_n50775_, new_n50776_, new_n50777_, new_n50778_,
    new_n50779_, new_n50780_, new_n50781_, new_n50782_, new_n50783_,
    new_n50784_, new_n50785_, new_n50786_, new_n50787_, new_n50788_,
    new_n50789_, new_n50790_, new_n50791_, new_n50792_, new_n50793_,
    new_n50794_, new_n50795_, new_n50796_, new_n50797_, new_n50798_,
    new_n50799_, new_n50800_, new_n50801_, new_n50802_, new_n50803_,
    new_n50804_, new_n50805_, new_n50806_, new_n50807_, new_n50808_,
    new_n50809_, new_n50810_, new_n50811_, new_n50812_, new_n50813_,
    new_n50814_, new_n50815_, new_n50816_, new_n50817_, new_n50818_,
    new_n50819_, new_n50820_, new_n50821_, new_n50822_, new_n50823_,
    new_n50824_, new_n50825_, new_n50826_, new_n50827_, new_n50828_,
    new_n50829_, new_n50830_, new_n50831_, new_n50832_, new_n50833_,
    new_n50834_, new_n50835_, new_n50836_, new_n50837_, new_n50838_,
    new_n50839_, new_n50840_, new_n50841_, new_n50842_, new_n50843_,
    new_n50844_, new_n50845_, new_n50846_, new_n50847_, new_n50848_,
    new_n50849_, new_n50850_, new_n50851_, new_n50852_, new_n50853_,
    new_n50854_, new_n50855_, new_n50856_, new_n50857_, new_n50858_,
    new_n50859_, new_n50860_, new_n50861_, new_n50862_, new_n50863_,
    new_n50864_, new_n50865_, new_n50866_, new_n50867_, new_n50868_,
    new_n50869_, new_n50870_, new_n50871_, new_n50872_, new_n50873_,
    new_n50874_, new_n50875_, new_n50876_, new_n50877_, new_n50878_,
    new_n50879_, new_n50880_, new_n50881_, new_n50882_, new_n50883_,
    new_n50884_, new_n50885_, new_n50886_, new_n50887_, new_n50888_,
    new_n50889_, new_n50890_, new_n50891_, new_n50892_, new_n50893_,
    new_n50894_, new_n50895_, new_n50896_, new_n50897_, new_n50898_,
    new_n50899_, new_n50900_, new_n50901_, new_n50902_, new_n50903_,
    new_n50904_, new_n50905_, new_n50906_, new_n50907_, new_n50908_,
    new_n50909_, new_n50910_, new_n50911_, new_n50912_, new_n50913_,
    new_n50914_, new_n50915_, new_n50916_, new_n50917_, new_n50918_,
    new_n50919_, new_n50920_, new_n50921_, new_n50922_, new_n50923_,
    new_n50924_, new_n50925_, new_n50926_, new_n50927_, new_n50928_,
    new_n50929_, new_n50930_, new_n50931_, new_n50932_, new_n50933_,
    new_n50934_, new_n50935_, new_n50936_, new_n50937_, new_n50938_,
    new_n50939_, new_n50940_, new_n50941_, new_n50942_, new_n50943_,
    new_n50944_, new_n50945_, new_n50946_, new_n50947_, new_n50948_,
    new_n50949_, new_n50950_, new_n50951_, new_n50952_, new_n50953_,
    new_n50954_, new_n50955_, new_n50956_, new_n50957_, new_n50958_,
    new_n50959_, new_n50960_, new_n50961_, new_n50962_, new_n50963_,
    new_n50964_, new_n50965_, new_n50966_, new_n50967_, new_n50968_,
    new_n50969_, new_n50970_, new_n50971_, new_n50972_, new_n50973_,
    new_n50974_, new_n50975_, new_n50976_, new_n50977_, new_n50978_,
    new_n50979_, new_n50980_, new_n50981_, new_n50982_, new_n50983_,
    new_n50984_, new_n50985_, new_n50986_, new_n50987_, new_n50988_,
    new_n50989_, new_n50990_, new_n50991_, new_n50992_, new_n50993_,
    new_n50994_, new_n50995_, new_n50996_, new_n50997_, new_n50998_,
    new_n50999_, new_n51000_, new_n51001_, new_n51002_, new_n51003_,
    new_n51004_, new_n51005_, new_n51006_, new_n51007_, new_n51008_,
    new_n51009_, new_n51010_, new_n51011_, new_n51012_, new_n51013_,
    new_n51014_, new_n51015_, new_n51016_, new_n51017_, new_n51018_,
    new_n51019_, new_n51020_, new_n51021_, new_n51022_, new_n51023_,
    new_n51024_, new_n51025_, new_n51026_, new_n51027_, new_n51028_,
    new_n51029_, new_n51030_, new_n51031_, new_n51032_, new_n51033_,
    new_n51034_, new_n51035_, new_n51036_, new_n51037_, new_n51038_,
    new_n51039_, new_n51040_, new_n51041_, new_n51042_, new_n51043_,
    new_n51044_, new_n51045_, new_n51046_, new_n51047_, new_n51048_,
    new_n51049_, new_n51050_, new_n51051_, new_n51052_, new_n51053_,
    new_n51054_, new_n51055_, new_n51056_, new_n51057_, new_n51058_,
    new_n51059_, new_n51060_, new_n51061_, new_n51062_, new_n51063_,
    new_n51064_, new_n51065_, new_n51066_, new_n51067_, new_n51068_,
    new_n51069_, new_n51070_, new_n51071_, new_n51072_, new_n51073_,
    new_n51074_, new_n51075_, new_n51076_, new_n51077_, new_n51078_,
    new_n51079_, new_n51080_, new_n51081_, new_n51082_, new_n51083_,
    new_n51084_, new_n51085_, new_n51086_, new_n51087_, new_n51088_,
    new_n51089_, new_n51090_, new_n51091_, new_n51092_, new_n51093_,
    new_n51094_, new_n51095_, new_n51096_, new_n51097_, new_n51098_,
    new_n51099_, new_n51100_, new_n51101_, new_n51102_, new_n51103_,
    new_n51104_, new_n51105_, new_n51106_, new_n51107_, new_n51108_,
    new_n51109_, new_n51110_, new_n51111_, new_n51112_, new_n51113_,
    new_n51114_, new_n51115_, new_n51116_, new_n51117_, new_n51118_,
    new_n51119_, new_n51120_, new_n51121_, new_n51122_, new_n51123_,
    new_n51124_, new_n51125_, new_n51126_, new_n51127_, new_n51128_,
    new_n51129_, new_n51130_, new_n51131_, new_n51132_, new_n51133_,
    new_n51134_, new_n51135_, new_n51136_, new_n51137_, new_n51138_,
    new_n51139_, new_n51140_, new_n51141_, new_n51142_, new_n51143_,
    new_n51144_, new_n51145_, new_n51146_, new_n51147_, new_n51148_,
    new_n51149_, new_n51150_, new_n51151_, new_n51152_, new_n51153_,
    new_n51154_, new_n51155_, new_n51156_, new_n51157_, new_n51158_,
    new_n51159_, new_n51160_, new_n51161_, new_n51162_, new_n51163_,
    new_n51164_, new_n51165_, new_n51166_, new_n51167_, new_n51168_,
    new_n51169_, new_n51170_, new_n51171_, new_n51172_, new_n51173_,
    new_n51174_, new_n51175_, new_n51176_, new_n51177_, new_n51178_,
    new_n51179_, new_n51180_, new_n51181_, new_n51182_, new_n51183_,
    new_n51184_, new_n51185_, new_n51186_, new_n51187_, new_n51188_,
    new_n51189_, new_n51190_, new_n51191_, new_n51192_, new_n51193_,
    new_n51194_, new_n51195_, new_n51196_, new_n51197_, new_n51198_,
    new_n51199_, new_n51200_, new_n51201_, new_n51202_, new_n51203_,
    new_n51204_, new_n51205_, new_n51206_, new_n51207_, new_n51208_,
    new_n51209_, new_n51210_, new_n51211_, new_n51212_, new_n51213_,
    new_n51214_, new_n51215_, new_n51216_, new_n51217_, new_n51218_,
    new_n51219_, new_n51220_, new_n51221_, new_n51222_, new_n51223_,
    new_n51224_, new_n51225_, new_n51226_, new_n51227_, new_n51228_,
    new_n51229_, new_n51230_, new_n51231_, new_n51232_, new_n51233_,
    new_n51234_, new_n51235_, new_n51236_, new_n51237_, new_n51238_,
    new_n51239_, new_n51240_, new_n51241_, new_n51242_, new_n51243_,
    new_n51244_, new_n51245_, new_n51246_, new_n51247_, new_n51248_,
    new_n51249_, new_n51250_, new_n51251_, new_n51252_, new_n51253_,
    new_n51254_, new_n51255_, new_n51256_, new_n51257_, new_n51258_,
    new_n51259_, new_n51260_, new_n51261_, new_n51262_, new_n51263_,
    new_n51264_, new_n51265_, new_n51266_, new_n51267_, new_n51268_,
    new_n51269_, new_n51270_, new_n51271_, new_n51272_, new_n51273_,
    new_n51274_, new_n51275_, new_n51276_, new_n51277_, new_n51278_,
    new_n51279_, new_n51280_, new_n51281_, new_n51282_, new_n51283_,
    new_n51284_, new_n51285_, new_n51286_, new_n51287_, new_n51288_,
    new_n51289_, new_n51290_, new_n51291_, new_n51292_, new_n51293_,
    new_n51294_, new_n51295_, new_n51296_, new_n51297_, new_n51298_,
    new_n51299_, new_n51300_, new_n51301_, new_n51302_, new_n51303_,
    new_n51304_, new_n51305_, new_n51306_, new_n51307_, new_n51308_,
    new_n51309_, new_n51310_, new_n51311_, new_n51312_, new_n51313_,
    new_n51314_, new_n51315_, new_n51316_, new_n51317_, new_n51318_,
    new_n51319_, new_n51320_, new_n51321_, new_n51322_, new_n51323_,
    new_n51324_, new_n51325_, new_n51326_, new_n51327_, new_n51328_,
    new_n51329_, new_n51330_, new_n51331_, new_n51332_, new_n51333_,
    new_n51334_, new_n51335_, new_n51336_, new_n51337_, new_n51338_,
    new_n51339_, new_n51340_, new_n51341_, new_n51342_, new_n51343_,
    new_n51344_, new_n51345_, new_n51346_, new_n51347_, new_n51348_,
    new_n51349_, new_n51350_, new_n51351_, new_n51352_, new_n51353_,
    new_n51354_, new_n51355_, new_n51356_, new_n51357_, new_n51358_,
    new_n51359_, new_n51360_, new_n51361_, new_n51362_, new_n51363_,
    new_n51364_, new_n51365_, new_n51366_, new_n51367_, new_n51368_,
    new_n51369_, new_n51370_, new_n51371_, new_n51372_, new_n51373_,
    new_n51374_, new_n51375_, new_n51376_, new_n51377_, new_n51378_,
    new_n51379_, new_n51380_, new_n51381_, new_n51382_, new_n51383_,
    new_n51384_, new_n51385_, new_n51386_, new_n51387_, new_n51388_,
    new_n51389_, new_n51390_, new_n51391_, new_n51392_, new_n51393_,
    new_n51394_, new_n51395_, new_n51396_, new_n51397_, new_n51398_,
    new_n51399_, new_n51400_, new_n51401_, new_n51402_, new_n51403_,
    new_n51404_, new_n51405_, new_n51406_, new_n51407_, new_n51408_,
    new_n51409_, new_n51410_, new_n51411_, new_n51412_, new_n51413_,
    new_n51414_, new_n51415_, new_n51416_, new_n51417_, new_n51418_,
    new_n51419_, new_n51420_, new_n51421_, new_n51422_, new_n51423_,
    new_n51424_, new_n51425_, new_n51426_, new_n51427_, new_n51428_,
    new_n51429_, new_n51430_, new_n51431_, new_n51432_, new_n51433_,
    new_n51434_, new_n51435_, new_n51436_, new_n51437_, new_n51438_,
    new_n51439_, new_n51440_, new_n51441_, new_n51442_, new_n51443_,
    new_n51444_, new_n51445_, new_n51446_, new_n51447_, new_n51448_,
    new_n51449_, new_n51450_, new_n51451_, new_n51452_, new_n51453_,
    new_n51454_, new_n51455_, new_n51456_, new_n51457_, new_n51458_,
    new_n51459_, new_n51460_, new_n51461_, new_n51462_, new_n51463_,
    new_n51464_, new_n51465_, new_n51466_, new_n51467_, new_n51468_,
    new_n51469_, new_n51470_, new_n51471_, new_n51472_, new_n51473_,
    new_n51474_, new_n51475_, new_n51476_, new_n51477_, new_n51478_,
    new_n51479_, new_n51480_, new_n51481_, new_n51482_, new_n51483_,
    new_n51484_, new_n51485_, new_n51486_, new_n51487_, new_n51488_,
    new_n51489_, new_n51490_, new_n51491_, new_n51492_, new_n51493_,
    new_n51494_, new_n51495_, new_n51496_, new_n51497_, new_n51498_,
    new_n51499_, new_n51500_, new_n51501_, new_n51502_, new_n51503_,
    new_n51504_, new_n51505_, new_n51506_, new_n51507_, new_n51508_,
    new_n51509_, new_n51510_, new_n51511_, new_n51512_, new_n51513_,
    new_n51514_, new_n51515_, new_n51516_, new_n51517_, new_n51518_,
    new_n51519_, new_n51520_, new_n51521_, new_n51522_, new_n51523_,
    new_n51524_, new_n51525_, new_n51526_, new_n51527_, new_n51528_,
    new_n51529_, new_n51530_, new_n51531_, new_n51532_, new_n51533_,
    new_n51534_, new_n51535_, new_n51536_, new_n51537_, new_n51538_,
    new_n51539_, new_n51540_, new_n51541_, new_n51542_, new_n51543_,
    new_n51544_, new_n51545_, new_n51546_, new_n51547_, new_n51548_,
    new_n51549_, new_n51550_, new_n51551_, new_n51552_, new_n51553_,
    new_n51554_, new_n51555_, new_n51556_, new_n51557_, new_n51558_,
    new_n51559_, new_n51560_, new_n51561_, new_n51562_, new_n51563_,
    new_n51564_, new_n51565_, new_n51566_, new_n51567_, new_n51568_,
    new_n51569_, new_n51570_, new_n51571_, new_n51572_, new_n51573_,
    new_n51574_, new_n51575_, new_n51576_, new_n51577_, new_n51578_,
    new_n51579_, new_n51580_, new_n51581_, new_n51582_, new_n51583_,
    new_n51584_, new_n51585_, new_n51586_, new_n51587_, new_n51588_,
    new_n51589_, new_n51590_, new_n51591_, new_n51592_, new_n51593_,
    new_n51594_, new_n51595_, new_n51596_, new_n51597_, new_n51598_,
    new_n51599_, new_n51600_, new_n51601_, new_n51602_, new_n51603_,
    new_n51604_, new_n51605_, new_n51606_, new_n51607_, new_n51608_,
    new_n51609_, new_n51610_, new_n51611_, new_n51612_, new_n51613_,
    new_n51614_, new_n51615_, new_n51616_, new_n51617_, new_n51618_,
    new_n51619_, new_n51620_, new_n51621_, new_n51622_, new_n51623_,
    new_n51624_, new_n51625_, new_n51626_, new_n51627_, new_n51628_,
    new_n51629_, new_n51630_, new_n51631_, new_n51632_, new_n51633_,
    new_n51634_, new_n51635_, new_n51636_, new_n51637_, new_n51638_,
    new_n51639_, new_n51640_, new_n51641_, new_n51642_, new_n51643_,
    new_n51644_, new_n51645_, new_n51646_, new_n51647_, new_n51648_,
    new_n51649_, new_n51650_, new_n51651_, new_n51652_, new_n51653_,
    new_n51654_, new_n51655_, new_n51656_, new_n51657_, new_n51658_,
    new_n51659_, new_n51660_, new_n51661_, new_n51662_, new_n51663_,
    new_n51664_, new_n51665_, new_n51666_, new_n51667_, new_n51668_,
    new_n51669_, new_n51670_, new_n51671_, new_n51672_, new_n51673_,
    new_n51674_, new_n51675_, new_n51676_, new_n51677_, new_n51678_,
    new_n51679_, new_n51680_, new_n51681_, new_n51682_, new_n51683_,
    new_n51684_, new_n51685_, new_n51686_, new_n51687_, new_n51688_,
    new_n51689_, new_n51690_, new_n51691_, new_n51692_, new_n51693_,
    new_n51694_, new_n51695_, new_n51696_, new_n51697_, new_n51698_,
    new_n51699_, new_n51700_, new_n51701_, new_n51702_, new_n51703_,
    new_n51704_, new_n51705_, new_n51706_, new_n51707_, new_n51708_,
    new_n51709_, new_n51710_, new_n51711_, new_n51712_, new_n51713_,
    new_n51714_, new_n51715_, new_n51716_, new_n51717_, new_n51718_,
    new_n51719_, new_n51720_, new_n51721_, new_n51722_, new_n51723_,
    new_n51724_, new_n51725_, new_n51726_, new_n51727_, new_n51728_,
    new_n51729_, new_n51730_, new_n51731_, new_n51732_, new_n51733_,
    new_n51734_, new_n51735_, new_n51736_, new_n51737_, new_n51738_,
    new_n51739_, new_n51740_, new_n51741_, new_n51742_, new_n51743_,
    new_n51744_, new_n51745_, new_n51746_, new_n51747_, new_n51748_,
    new_n51749_, new_n51750_, new_n51751_, new_n51752_, new_n51753_,
    new_n51754_, new_n51755_, new_n51756_, new_n51757_, new_n51758_,
    new_n51759_, new_n51760_, new_n51761_, new_n51762_, new_n51763_,
    new_n51764_, new_n51765_, new_n51766_, new_n51767_, new_n51768_,
    new_n51769_, new_n51770_, new_n51771_, new_n51772_, new_n51773_,
    new_n51774_, new_n51775_, new_n51776_, new_n51777_, new_n51778_,
    new_n51779_, new_n51780_, new_n51781_, new_n51782_, new_n51783_,
    new_n51784_, new_n51785_, new_n51786_, new_n51787_, new_n51788_,
    new_n51789_, new_n51790_, new_n51791_, new_n51792_, new_n51793_,
    new_n51794_, new_n51795_, new_n51796_, new_n51797_, new_n51798_,
    new_n51799_, new_n51800_, new_n51801_, new_n51802_, new_n51803_,
    new_n51804_, new_n51805_, new_n51806_, new_n51807_, new_n51808_,
    new_n51809_, new_n51810_, new_n51811_, new_n51812_, new_n51813_,
    new_n51814_, new_n51815_, new_n51816_, new_n51817_, new_n51818_,
    new_n51819_, new_n51820_, new_n51821_, new_n51822_, new_n51823_,
    new_n51824_, new_n51825_, new_n51826_, new_n51827_, new_n51828_,
    new_n51829_, new_n51830_, new_n51831_, new_n51832_, new_n51833_,
    new_n51834_, new_n51835_, new_n51836_, new_n51837_, new_n51838_,
    new_n51839_, new_n51840_, new_n51841_, new_n51842_, new_n51843_,
    new_n51844_, new_n51845_, new_n51846_, new_n51847_, new_n51848_,
    new_n51849_, new_n51850_, new_n51851_, new_n51852_, new_n51853_,
    new_n51854_, new_n51855_, new_n51856_, new_n51857_, new_n51858_,
    new_n51859_, new_n51860_, new_n51861_, new_n51862_, new_n51863_,
    new_n51864_, new_n51865_, new_n51866_, new_n51867_, new_n51868_,
    new_n51869_, new_n51870_, new_n51871_, new_n51872_, new_n51873_,
    new_n51874_, new_n51875_, new_n51876_, new_n51877_, new_n51878_,
    new_n51879_, new_n51880_, new_n51881_, new_n51882_, new_n51883_,
    new_n51884_, new_n51885_, new_n51886_, new_n51887_, new_n51888_,
    new_n51889_, new_n51890_, new_n51891_, new_n51892_, new_n51893_,
    new_n51894_, new_n51895_, new_n51896_, new_n51897_, new_n51898_,
    new_n51899_, new_n51900_, new_n51901_, new_n51902_, new_n51903_,
    new_n51904_, new_n51905_, new_n51906_, new_n51907_, new_n51908_,
    new_n51909_, new_n51910_, new_n51911_, new_n51912_, new_n51913_,
    new_n51914_, new_n51915_, new_n51916_, new_n51917_, new_n51918_,
    new_n51919_, new_n51920_, new_n51921_, new_n51922_, new_n51923_,
    new_n51924_, new_n51925_, new_n51926_, new_n51927_, new_n51928_,
    new_n51929_, new_n51930_, new_n51931_, new_n51932_, new_n51933_,
    new_n51934_, new_n51935_, new_n51936_, new_n51937_, new_n51938_,
    new_n51939_, new_n51940_, new_n51941_, new_n51942_, new_n51943_,
    new_n51944_, new_n51945_, new_n51946_, new_n51947_, new_n51948_,
    new_n51949_, new_n51950_, new_n51951_, new_n51952_, new_n51953_,
    new_n51954_, new_n51955_, new_n51956_, new_n51957_, new_n51958_,
    new_n51959_, new_n51960_, new_n51961_, new_n51962_, new_n51963_,
    new_n51964_, new_n51965_, new_n51966_, new_n51967_, new_n51968_,
    new_n51969_, new_n51970_, new_n51971_, new_n51972_, new_n51973_,
    new_n51974_, new_n51975_, new_n51976_, new_n51977_, new_n51978_,
    new_n51979_, new_n51980_, new_n51981_, new_n51982_, new_n51983_,
    new_n51984_, new_n51985_, new_n51986_, new_n51987_, new_n51988_,
    new_n51989_, new_n51990_, new_n51991_, new_n51992_, new_n51993_,
    new_n51994_, new_n51995_, new_n51996_, new_n51997_, new_n51998_,
    new_n51999_, new_n52000_, new_n52001_, new_n52002_, new_n52003_,
    new_n52004_, new_n52005_, new_n52006_, new_n52007_, new_n52008_,
    new_n52009_, new_n52010_, new_n52011_, new_n52012_, new_n52013_,
    new_n52014_, new_n52015_, new_n52016_, new_n52017_, new_n52018_,
    new_n52019_, new_n52020_, new_n52021_, new_n52022_, new_n52023_,
    new_n52024_, new_n52025_, new_n52026_, new_n52027_, new_n52028_,
    new_n52029_, new_n52030_, new_n52031_, new_n52032_, new_n52033_,
    new_n52034_, new_n52035_, new_n52036_, new_n52037_, new_n52038_,
    new_n52039_, new_n52040_, new_n52041_, new_n52042_, new_n52043_,
    new_n52044_, new_n52045_, new_n52046_, new_n52047_, new_n52048_,
    new_n52049_, new_n52050_, new_n52051_, new_n52052_, new_n52053_,
    new_n52054_, new_n52055_, new_n52056_, new_n52057_, new_n52058_,
    new_n52059_, new_n52060_, new_n52061_, new_n52062_, new_n52063_,
    new_n52064_, new_n52065_, new_n52066_, new_n52067_, new_n52068_,
    new_n52069_, new_n52070_, new_n52071_, new_n52072_, new_n52073_,
    new_n52074_, new_n52075_, new_n52076_, new_n52077_, new_n52078_,
    new_n52079_, new_n52080_, new_n52081_, new_n52082_, new_n52083_,
    new_n52084_, new_n52085_, new_n52086_, new_n52087_, new_n52088_,
    new_n52089_, new_n52090_, new_n52091_, new_n52092_, new_n52093_,
    new_n52094_, new_n52095_, new_n52096_, new_n52097_, new_n52098_,
    new_n52099_, new_n52100_, new_n52101_, new_n52102_, new_n52103_,
    new_n52104_, new_n52105_, new_n52106_, new_n52107_, new_n52108_,
    new_n52109_, new_n52110_, new_n52111_, new_n52112_, new_n52113_,
    new_n52114_, new_n52115_, new_n52116_, new_n52117_, new_n52118_,
    new_n52119_, new_n52120_, new_n52121_, new_n52122_, new_n52123_,
    new_n52124_, new_n52125_, new_n52126_, new_n52127_, new_n52128_,
    new_n52129_, new_n52130_, new_n52131_, new_n52132_, new_n52133_,
    new_n52134_, new_n52135_, new_n52136_, new_n52137_, new_n52138_,
    new_n52139_, new_n52140_, new_n52141_, new_n52142_, new_n52143_,
    new_n52144_, new_n52145_, new_n52146_, new_n52147_, new_n52148_,
    new_n52149_, new_n52150_, new_n52151_, new_n52152_, new_n52153_,
    new_n52154_, new_n52155_, new_n52156_, new_n52157_, new_n52158_,
    new_n52159_, new_n52160_, new_n52161_, new_n52162_, new_n52163_,
    new_n52164_, new_n52165_, new_n52166_, new_n52167_, new_n52168_,
    new_n52169_, new_n52170_, new_n52171_, new_n52172_, new_n52173_,
    new_n52174_, new_n52175_, new_n52176_, new_n52177_, new_n52178_,
    new_n52179_, new_n52180_, new_n52181_, new_n52182_, new_n52183_,
    new_n52184_, new_n52185_, new_n52186_, new_n52187_, new_n52188_,
    new_n52189_, new_n52190_, new_n52191_, new_n52192_, new_n52193_,
    new_n52194_, new_n52195_, new_n52196_, new_n52197_, new_n52198_,
    new_n52199_, new_n52200_, new_n52201_, new_n52202_, new_n52203_,
    new_n52204_, new_n52205_, new_n52206_, new_n52207_, new_n52208_,
    new_n52209_, new_n52210_, new_n52211_, new_n52212_, new_n52213_,
    new_n52214_, new_n52215_, new_n52216_, new_n52217_, new_n52218_,
    new_n52219_, new_n52220_, new_n52221_, new_n52222_, new_n52223_,
    new_n52224_, new_n52225_, new_n52226_, new_n52227_, new_n52228_,
    new_n52229_, new_n52230_, new_n52231_, new_n52232_, new_n52233_,
    new_n52234_, new_n52235_, new_n52236_, new_n52237_, new_n52238_,
    new_n52239_, new_n52240_, new_n52241_, new_n52242_, new_n52243_,
    new_n52244_, new_n52245_, new_n52246_, new_n52247_, new_n52248_,
    new_n52249_, new_n52250_, new_n52251_, new_n52252_, new_n52253_,
    new_n52254_, new_n52255_, new_n52256_, new_n52257_, new_n52258_,
    new_n52259_, new_n52260_, new_n52261_, new_n52262_, new_n52263_,
    new_n52264_, new_n52265_, new_n52266_, new_n52267_, new_n52268_,
    new_n52269_, new_n52270_, new_n52271_, new_n52272_, new_n52273_,
    new_n52274_, new_n52275_, new_n52276_, new_n52277_, new_n52278_,
    new_n52279_, new_n52280_, new_n52281_, new_n52282_, new_n52283_,
    new_n52284_, new_n52285_, new_n52286_, new_n52287_, new_n52288_,
    new_n52289_, new_n52290_, new_n52291_, new_n52292_, new_n52293_,
    new_n52294_, new_n52295_, new_n52296_, new_n52297_, new_n52298_,
    new_n52299_, new_n52300_, new_n52301_, new_n52302_, new_n52303_,
    new_n52304_, new_n52305_, new_n52306_, new_n52307_, new_n52308_,
    new_n52309_, new_n52310_, new_n52311_, new_n52312_, new_n52313_,
    new_n52314_, new_n52315_, new_n52316_, new_n52317_, new_n52318_,
    new_n52319_, new_n52320_, new_n52321_, new_n52322_, new_n52323_,
    new_n52324_, new_n52325_, new_n52326_, new_n52327_, new_n52328_,
    new_n52329_, new_n52330_, new_n52331_, new_n52332_, new_n52333_,
    new_n52334_, new_n52335_, new_n52336_, new_n52337_, new_n52338_,
    new_n52339_, new_n52340_, new_n52341_, new_n52342_, new_n52343_,
    new_n52344_, new_n52345_, new_n52346_, new_n52347_, new_n52348_,
    new_n52349_, new_n52350_, new_n52351_, new_n52352_, new_n52353_,
    new_n52354_, new_n52355_, new_n52356_, new_n52357_, new_n52358_,
    new_n52359_, new_n52360_, new_n52361_, new_n52362_, new_n52363_,
    new_n52364_, new_n52365_, new_n52366_, new_n52367_, new_n52368_,
    new_n52369_, new_n52370_, new_n52371_, new_n52372_, new_n52373_,
    new_n52374_, new_n52375_, new_n52376_, new_n52377_, new_n52378_,
    new_n52379_, new_n52380_, new_n52381_, new_n52382_, new_n52383_,
    new_n52384_, new_n52385_, new_n52386_, new_n52387_, new_n52388_,
    new_n52389_, new_n52390_, new_n52391_, new_n52392_, new_n52393_,
    new_n52394_, new_n52395_, new_n52396_, new_n52397_, new_n52398_,
    new_n52399_, new_n52400_, new_n52401_, new_n52402_, new_n52403_,
    new_n52404_, new_n52405_, new_n52406_, new_n52407_, new_n52408_,
    new_n52409_, new_n52410_, new_n52411_, new_n52412_, new_n52413_,
    new_n52414_, new_n52415_, new_n52416_, new_n52417_, new_n52418_,
    new_n52419_, new_n52420_, new_n52421_, new_n52422_, new_n52423_,
    new_n52424_, new_n52425_, new_n52426_, new_n52427_, new_n52428_,
    new_n52429_, new_n52430_, new_n52431_, new_n52432_, new_n52433_,
    new_n52434_, new_n52435_, new_n52436_, new_n52437_, new_n52438_,
    new_n52439_, new_n52440_, new_n52441_, new_n52442_, new_n52443_,
    new_n52444_, new_n52445_, new_n52446_, new_n52447_, new_n52448_,
    new_n52449_, new_n52450_, new_n52451_, new_n52452_, new_n52453_,
    new_n52454_, new_n52455_, new_n52456_, new_n52457_, new_n52458_,
    new_n52459_, new_n52460_, new_n52461_, new_n52462_, new_n52463_,
    new_n52464_, new_n52465_, new_n52466_, new_n52467_, new_n52468_,
    new_n52469_, new_n52470_, new_n52471_, new_n52472_, new_n52473_,
    new_n52474_, new_n52475_, new_n52476_, new_n52477_, new_n52478_,
    new_n52479_, new_n52480_, new_n52481_, new_n52482_, new_n52483_,
    new_n52484_, new_n52485_, new_n52486_, new_n52487_, new_n52488_,
    new_n52489_, new_n52490_, new_n52491_, new_n52492_, new_n52493_,
    new_n52494_, new_n52495_, new_n52496_, new_n52497_, new_n52498_,
    new_n52499_, new_n52500_, new_n52501_, new_n52502_, new_n52503_,
    new_n52504_, new_n52505_, new_n52506_, new_n52507_, new_n52508_,
    new_n52509_, new_n52510_, new_n52511_, new_n52512_, new_n52513_,
    new_n52514_, new_n52515_, new_n52516_, new_n52517_, new_n52518_,
    new_n52519_, new_n52520_, new_n52521_, new_n52522_, new_n52523_,
    new_n52524_, new_n52525_, new_n52526_, new_n52527_, new_n52528_,
    new_n52529_, new_n52530_, new_n52531_, new_n52532_, new_n52533_,
    new_n52534_, new_n52535_, new_n52536_, new_n52537_, new_n52538_,
    new_n52539_, new_n52540_, new_n52541_, new_n52542_, new_n52543_,
    new_n52544_, new_n52545_, new_n52546_, new_n52547_, new_n52548_,
    new_n52549_, new_n52550_, new_n52551_, new_n52552_, new_n52553_,
    new_n52554_, new_n52555_, new_n52556_, new_n52557_, new_n52558_,
    new_n52559_, new_n52560_, new_n52561_, new_n52562_, new_n52563_,
    new_n52564_, new_n52565_, new_n52566_, new_n52567_, new_n52568_,
    new_n52569_, new_n52570_, new_n52571_, new_n52572_, new_n52573_,
    new_n52574_, new_n52575_, new_n52576_, new_n52577_, new_n52578_,
    new_n52579_, new_n52580_, new_n52581_, new_n52582_, new_n52583_,
    new_n52584_, new_n52585_, new_n52586_, new_n52587_, new_n52588_,
    new_n52589_, new_n52590_, new_n52591_, new_n52592_, new_n52593_,
    new_n52594_, new_n52595_, new_n52596_, new_n52597_, new_n52598_,
    new_n52599_, new_n52600_, new_n52601_, new_n52602_, new_n52603_,
    new_n52604_, new_n52605_, new_n52606_, new_n52607_, new_n52608_,
    new_n52609_, new_n52610_, new_n52611_, new_n52612_, new_n52613_,
    new_n52614_, new_n52615_, new_n52616_, new_n52617_, new_n52618_,
    new_n52619_, new_n52620_, new_n52621_, new_n52622_, new_n52623_,
    new_n52624_, new_n52625_, new_n52626_, new_n52627_, new_n52628_,
    new_n52629_, new_n52630_, new_n52631_, new_n52632_, new_n52633_,
    new_n52634_, new_n52635_, new_n52636_, new_n52637_, new_n52638_,
    new_n52639_, new_n52640_, new_n52641_, new_n52642_, new_n52643_,
    new_n52644_, new_n52645_, new_n52646_, new_n52647_, new_n52648_,
    new_n52649_, new_n52650_, new_n52651_, new_n52652_, new_n52653_,
    new_n52654_, new_n52655_, new_n52656_, new_n52657_, new_n52658_,
    new_n52659_, new_n52660_, new_n52661_, new_n52662_, new_n52663_,
    new_n52664_, new_n52665_, new_n52666_, new_n52667_, new_n52668_,
    new_n52669_, new_n52670_, new_n52671_, new_n52672_, new_n52673_,
    new_n52674_, new_n52675_, new_n52676_, new_n52677_, new_n52678_,
    new_n52679_, new_n52680_, new_n52681_, new_n52682_, new_n52683_,
    new_n52684_, new_n52685_, new_n52686_, new_n52687_, new_n52688_,
    new_n52689_, new_n52690_, new_n52691_, new_n52692_, new_n52693_,
    new_n52694_, new_n52695_, new_n52696_, new_n52697_, new_n52698_,
    new_n52699_, new_n52700_, new_n52701_, new_n52702_, new_n52703_,
    new_n52704_, new_n52705_, new_n52706_, new_n52707_, new_n52708_,
    new_n52709_, new_n52710_, new_n52711_, new_n52712_, new_n52713_,
    new_n52714_, new_n52715_, new_n52716_, new_n52717_, new_n52718_,
    new_n52719_, new_n52720_, new_n52721_, new_n52722_, new_n52723_,
    new_n52724_, new_n52725_, new_n52726_, new_n52727_, new_n52728_,
    new_n52729_, new_n52730_, new_n52731_, new_n52732_, new_n52733_,
    new_n52734_, new_n52735_, new_n52736_, new_n52737_, new_n52738_,
    new_n52739_, new_n52740_, new_n52741_, new_n52742_, new_n52743_,
    new_n52744_, new_n52745_, new_n52746_, new_n52747_, new_n52748_,
    new_n52749_, new_n52750_, new_n52751_, new_n52752_, new_n52753_,
    new_n52754_, new_n52755_, new_n52756_, new_n52757_, new_n52758_,
    new_n52759_, new_n52760_, new_n52761_, new_n52762_, new_n52763_,
    new_n52764_, new_n52765_, new_n52766_, new_n52767_, new_n52768_,
    new_n52769_, new_n52770_, new_n52771_, new_n52772_, new_n52773_,
    new_n52774_, new_n52775_, new_n52776_, new_n52777_, new_n52778_,
    new_n52779_, new_n52780_, new_n52781_, new_n52782_, new_n52783_,
    new_n52784_, new_n52785_, new_n52786_, new_n52787_, new_n52788_,
    new_n52789_, new_n52790_, new_n52791_, new_n52792_, new_n52793_,
    new_n52794_, new_n52795_, new_n52796_, new_n52797_, new_n52798_,
    new_n52799_, new_n52800_, new_n52801_, new_n52802_, new_n52803_,
    new_n52804_, new_n52805_, new_n52806_, new_n52807_, new_n52808_,
    new_n52809_, new_n52810_, new_n52811_, new_n52812_, new_n52813_,
    new_n52814_, new_n52815_, new_n52816_, new_n52817_, new_n52818_,
    new_n52819_, new_n52820_, new_n52821_, new_n52822_, new_n52823_,
    new_n52824_, new_n52825_, new_n52826_, new_n52827_, new_n52828_,
    new_n52829_, new_n52830_, new_n52831_, new_n52832_, new_n52833_,
    new_n52834_, new_n52835_, new_n52836_, new_n52837_, new_n52838_,
    new_n52839_, new_n52840_, new_n52841_, new_n52842_, new_n52843_,
    new_n52844_, new_n52845_, new_n52846_, new_n52847_, new_n52848_,
    new_n52849_, new_n52850_, new_n52851_, new_n52852_, new_n52853_,
    new_n52854_, new_n52855_, new_n52856_, new_n52857_, new_n52858_,
    new_n52859_, new_n52860_, new_n52861_, new_n52862_, new_n52863_,
    new_n52864_, new_n52865_, new_n52866_, new_n52867_, new_n52868_,
    new_n52869_, new_n52870_, new_n52871_, new_n52872_, new_n52873_,
    new_n52874_, new_n52875_, new_n52876_, new_n52877_, new_n52878_,
    new_n52879_, new_n52880_, new_n52881_, new_n52882_, new_n52883_,
    new_n52884_, new_n52885_, new_n52886_, new_n52887_, new_n52888_,
    new_n52889_, new_n52890_, new_n52891_, new_n52892_, new_n52893_,
    new_n52894_, new_n52895_, new_n52896_, new_n52897_, new_n52898_,
    new_n52899_, new_n52900_, new_n52901_, new_n52902_, new_n52903_,
    new_n52904_, new_n52905_, new_n52906_, new_n52907_, new_n52908_,
    new_n52909_, new_n52910_, new_n52911_, new_n52912_, new_n52913_,
    new_n52914_, new_n52915_, new_n52916_, new_n52917_, new_n52918_,
    new_n52919_, new_n52920_, new_n52921_, new_n52922_, new_n52923_,
    new_n52924_, new_n52925_, new_n52926_, new_n52927_, new_n52928_,
    new_n52929_, new_n52930_, new_n52931_, new_n52932_, new_n52933_,
    new_n52934_, new_n52935_, new_n52936_, new_n52937_, new_n52938_,
    new_n52939_, new_n52940_, new_n52941_, new_n52942_, new_n52943_,
    new_n52944_, new_n52945_, new_n52946_, new_n52947_, new_n52948_,
    new_n52949_, new_n52950_, new_n52951_, new_n52952_, new_n52953_,
    new_n52954_, new_n52955_, new_n52956_, new_n52957_, new_n52958_,
    new_n52959_, new_n52960_, new_n52961_, new_n52962_, new_n52963_,
    new_n52964_, new_n52965_, new_n52966_, new_n52967_, new_n52968_,
    new_n52969_, new_n52970_, new_n52971_, new_n52972_, new_n52973_,
    new_n52974_, new_n52975_, new_n52976_, new_n52977_, new_n52978_,
    new_n52979_, new_n52980_, new_n52981_, new_n52982_, new_n52983_,
    new_n52984_, new_n52985_, new_n52986_, new_n52987_, new_n52988_,
    new_n52989_, new_n52990_, new_n52991_, new_n52992_, new_n52993_,
    new_n52994_, new_n52995_, new_n52996_, new_n52997_, new_n52998_,
    new_n52999_, new_n53000_, new_n53001_, new_n53002_, new_n53003_,
    new_n53004_, new_n53005_, new_n53006_, new_n53007_, new_n53008_,
    new_n53009_, new_n53010_, new_n53011_, new_n53012_, new_n53013_,
    new_n53014_, new_n53015_, new_n53016_, new_n53017_, new_n53018_,
    new_n53019_, new_n53020_, new_n53021_, new_n53022_, new_n53023_,
    new_n53024_, new_n53025_, new_n53026_, new_n53027_, new_n53028_,
    new_n53029_, new_n53030_, new_n53031_, new_n53032_, new_n53033_,
    new_n53034_, new_n53035_, new_n53036_, new_n53037_, new_n53038_,
    new_n53039_, new_n53040_, new_n53041_, new_n53042_, new_n53043_,
    new_n53044_, new_n53045_, new_n53046_, new_n53047_, new_n53048_,
    new_n53049_, new_n53050_, new_n53051_, new_n53052_, new_n53053_,
    new_n53054_, new_n53055_, new_n53056_, new_n53057_, new_n53058_,
    new_n53059_, new_n53060_, new_n53061_, new_n53062_, new_n53063_,
    new_n53064_, new_n53065_, new_n53066_, new_n53067_, new_n53068_,
    new_n53069_, new_n53070_, new_n53071_, new_n53072_, new_n53073_,
    new_n53074_, new_n53075_, new_n53076_, new_n53077_, new_n53078_,
    new_n53079_, new_n53080_, new_n53081_, new_n53082_, new_n53083_,
    new_n53084_, new_n53085_, new_n53086_, new_n53087_, new_n53088_,
    new_n53089_, new_n53090_, new_n53091_, new_n53092_, new_n53093_,
    new_n53094_, new_n53095_, new_n53096_, new_n53097_, new_n53098_,
    new_n53099_, new_n53100_, new_n53101_, new_n53102_, new_n53103_,
    new_n53104_, new_n53105_, new_n53106_, new_n53107_, new_n53108_,
    new_n53109_, new_n53110_, new_n53111_, new_n53112_, new_n53113_,
    new_n53114_, new_n53115_, new_n53116_, new_n53117_, new_n53118_,
    new_n53119_, new_n53120_, new_n53121_, new_n53122_, new_n53123_,
    new_n53124_, new_n53125_, new_n53126_, new_n53127_, new_n53128_,
    new_n53129_, new_n53130_, new_n53131_, new_n53132_, new_n53133_,
    new_n53134_, new_n53135_, new_n53136_, new_n53137_, new_n53138_,
    new_n53139_, new_n53140_, new_n53141_, new_n53142_, new_n53143_,
    new_n53144_, new_n53145_, new_n53146_, new_n53147_, new_n53148_,
    new_n53149_, new_n53150_, new_n53151_, new_n53152_, new_n53153_,
    new_n53154_, new_n53155_, new_n53156_, new_n53157_, new_n53158_,
    new_n53159_, new_n53160_, new_n53161_, new_n53162_, new_n53163_,
    new_n53164_, new_n53165_, new_n53166_, new_n53167_, new_n53168_,
    new_n53169_, new_n53170_, new_n53171_, new_n53172_, new_n53173_,
    new_n53174_, new_n53175_, new_n53176_, new_n53177_, new_n53178_,
    new_n53179_, new_n53180_, new_n53181_, new_n53182_, new_n53183_,
    new_n53184_, new_n53185_, new_n53186_, new_n53187_, new_n53188_,
    new_n53189_, new_n53190_, new_n53191_, new_n53192_, new_n53193_,
    new_n53194_, new_n53195_, new_n53196_, new_n53197_, new_n53198_,
    new_n53199_, new_n53200_, new_n53201_, new_n53202_, new_n53203_,
    new_n53204_, new_n53205_, new_n53206_, new_n53207_, new_n53208_,
    new_n53209_, new_n53210_, new_n53211_, new_n53212_, new_n53213_,
    new_n53214_, new_n53215_, new_n53216_, new_n53217_, new_n53218_,
    new_n53219_, new_n53220_, new_n53221_, new_n53222_, new_n53223_,
    new_n53224_, new_n53225_, new_n53226_, new_n53227_, new_n53228_,
    new_n53229_, new_n53230_, new_n53231_, new_n53232_, new_n53233_,
    new_n53234_, new_n53235_, new_n53236_, new_n53237_, new_n53238_,
    new_n53239_, new_n53240_, new_n53241_, new_n53242_, new_n53243_,
    new_n53244_, new_n53245_, new_n53246_, new_n53247_, new_n53248_,
    new_n53249_, new_n53250_, new_n53251_, new_n53252_, new_n53253_,
    new_n53254_, new_n53255_, new_n53256_, new_n53257_, new_n53258_,
    new_n53259_, new_n53260_, new_n53261_, new_n53262_, new_n53263_,
    new_n53264_, new_n53265_, new_n53266_, new_n53267_, new_n53268_,
    new_n53269_, new_n53270_, new_n53271_, new_n53272_, new_n53273_,
    new_n53274_, new_n53275_, new_n53276_, new_n53277_, new_n53278_,
    new_n53279_, new_n53280_, new_n53281_, new_n53282_, new_n53283_,
    new_n53284_, new_n53285_, new_n53286_, new_n53287_, new_n53288_,
    new_n53289_, new_n53290_, new_n53291_, new_n53292_, new_n53293_,
    new_n53294_, new_n53295_, new_n53296_, new_n53297_, new_n53298_,
    new_n53299_, new_n53300_, new_n53301_, new_n53302_, new_n53303_,
    new_n53304_, new_n53305_, new_n53306_, new_n53307_, new_n53308_,
    new_n53309_, new_n53310_, new_n53311_, new_n53312_, new_n53313_,
    new_n53314_, new_n53315_, new_n53316_, new_n53317_, new_n53318_,
    new_n53319_, new_n53320_, new_n53321_, new_n53322_, new_n53323_,
    new_n53324_, new_n53325_, new_n53326_, new_n53327_, new_n53328_,
    new_n53329_, new_n53330_, new_n53331_, new_n53332_, new_n53333_,
    new_n53334_, new_n53335_, new_n53336_, new_n53337_, new_n53338_,
    new_n53339_, new_n53340_, new_n53341_, new_n53342_, new_n53343_,
    new_n53344_, new_n53345_, new_n53346_, new_n53347_, new_n53348_,
    new_n53349_, new_n53350_, new_n53351_, new_n53352_, new_n53353_,
    new_n53354_, new_n53355_, new_n53356_, new_n53357_, new_n53358_,
    new_n53359_, new_n53360_, new_n53361_, new_n53362_, new_n53363_,
    new_n53364_, new_n53365_, new_n53366_, new_n53367_, new_n53368_,
    new_n53369_, new_n53370_, new_n53371_, new_n53372_, new_n53373_,
    new_n53374_, new_n53375_, new_n53376_, new_n53377_, new_n53378_,
    new_n53379_, new_n53380_, new_n53381_, new_n53382_, new_n53383_,
    new_n53384_, new_n53385_, new_n53386_, new_n53387_, new_n53388_,
    new_n53389_, new_n53390_, new_n53391_, new_n53392_, new_n53393_,
    new_n53394_, new_n53395_, new_n53396_, new_n53397_, new_n53398_,
    new_n53399_, new_n53400_, new_n53401_, new_n53402_, new_n53403_,
    new_n53404_, new_n53405_, new_n53406_, new_n53407_, new_n53408_,
    new_n53409_, new_n53410_, new_n53411_, new_n53412_, new_n53413_,
    new_n53414_, new_n53415_, new_n53416_, new_n53417_, new_n53418_,
    new_n53419_, new_n53420_, new_n53421_, new_n53422_, new_n53423_,
    new_n53424_, new_n53425_, new_n53426_, new_n53427_, new_n53428_,
    new_n53429_, new_n53430_, new_n53431_, new_n53432_, new_n53433_,
    new_n53434_, new_n53435_, new_n53436_, new_n53437_, new_n53438_,
    new_n53439_, new_n53440_, new_n53441_, new_n53442_, new_n53443_,
    new_n53444_, new_n53445_, new_n53446_, new_n53447_, new_n53448_,
    new_n53449_, new_n53450_, new_n53451_, new_n53452_, new_n53453_,
    new_n53454_, new_n53455_, new_n53456_, new_n53457_, new_n53458_,
    new_n53459_, new_n53460_, new_n53461_, new_n53462_, new_n53463_,
    new_n53464_, new_n53465_, new_n53466_, new_n53467_, new_n53468_,
    new_n53469_, new_n53470_, new_n53471_, new_n53472_, new_n53473_,
    new_n53474_, new_n53475_, new_n53476_, new_n53477_, new_n53478_,
    new_n53479_, new_n53480_, new_n53481_, new_n53482_, new_n53483_,
    new_n53484_, new_n53485_, new_n53486_, new_n53487_, new_n53488_,
    new_n53489_, new_n53490_, new_n53491_, new_n53492_, new_n53493_,
    new_n53494_, new_n53495_, new_n53496_, new_n53497_, new_n53498_,
    new_n53499_, new_n53500_, new_n53501_, new_n53502_, new_n53503_,
    new_n53504_, new_n53505_, new_n53506_, new_n53507_, new_n53508_,
    new_n53509_, new_n53510_, new_n53511_, new_n53512_, new_n53513_,
    new_n53514_, new_n53515_, new_n53516_, new_n53517_, new_n53518_,
    new_n53519_, new_n53520_, new_n53521_, new_n53522_, new_n53523_,
    new_n53524_, new_n53525_, new_n53526_, new_n53527_, new_n53528_,
    new_n53529_, new_n53530_, new_n53531_, new_n53532_, new_n53533_,
    new_n53534_, new_n53535_, new_n53536_, new_n53537_, new_n53538_,
    new_n53539_, new_n53540_, new_n53541_, new_n53542_, new_n53543_,
    new_n53544_, new_n53545_, new_n53546_, new_n53547_, new_n53548_,
    new_n53549_, new_n53550_, new_n53551_, new_n53552_, new_n53553_,
    new_n53554_, new_n53555_, new_n53556_, new_n53557_, new_n53558_,
    new_n53559_, new_n53560_, new_n53561_, new_n53562_, new_n53563_,
    new_n53564_, new_n53565_, new_n53566_, new_n53567_, new_n53568_,
    new_n53569_, new_n53570_, new_n53571_, new_n53572_, new_n53573_,
    new_n53574_, new_n53575_, new_n53576_, new_n53577_, new_n53578_,
    new_n53579_, new_n53580_, new_n53581_, new_n53582_, new_n53583_,
    new_n53584_, new_n53585_, new_n53586_, new_n53587_, new_n53588_,
    new_n53589_, new_n53590_, new_n53591_, new_n53592_, new_n53593_,
    new_n53594_, new_n53595_, new_n53596_, new_n53597_, new_n53598_,
    new_n53599_, new_n53600_, new_n53601_, new_n53602_, new_n53603_,
    new_n53604_, new_n53605_, new_n53606_, new_n53607_, new_n53608_,
    new_n53609_, new_n53610_, new_n53611_, new_n53612_, new_n53613_,
    new_n53614_, new_n53615_, new_n53616_, new_n53617_, new_n53618_,
    new_n53619_, new_n53620_, new_n53621_, new_n53622_, new_n53623_,
    new_n53624_, new_n53625_, new_n53626_, new_n53627_, new_n53628_,
    new_n53629_, new_n53630_, new_n53631_, new_n53632_, new_n53633_,
    new_n53634_, new_n53635_, new_n53636_, new_n53637_, new_n53638_,
    new_n53639_, new_n53640_, new_n53641_, new_n53642_, new_n53643_,
    new_n53644_, new_n53645_, new_n53646_, new_n53647_, new_n53648_,
    new_n53649_, new_n53650_, new_n53651_, new_n53652_, new_n53653_,
    new_n53654_, new_n53655_, new_n53656_, new_n53657_, new_n53658_,
    new_n53659_, new_n53660_, new_n53661_, new_n53662_, new_n53663_,
    new_n53664_, new_n53665_, new_n53666_, new_n53667_, new_n53668_,
    new_n53669_, new_n53670_, new_n53671_, new_n53672_, new_n53673_,
    new_n53674_, new_n53675_, new_n53676_, new_n53677_, new_n53678_,
    new_n53679_, new_n53680_, new_n53681_, new_n53682_, new_n53683_,
    new_n53684_, new_n53685_, new_n53686_, new_n53687_, new_n53688_,
    new_n53689_, new_n53690_, new_n53691_, new_n53692_, new_n53693_,
    new_n53694_, new_n53695_, new_n53696_, new_n53697_, new_n53698_,
    new_n53699_, new_n53700_, new_n53701_, new_n53702_, new_n53703_,
    new_n53704_, new_n53705_, new_n53706_, new_n53707_, new_n53708_,
    new_n53709_, new_n53710_, new_n53711_, new_n53712_, new_n53713_,
    new_n53714_, new_n53715_, new_n53716_, new_n53717_, new_n53718_,
    new_n53719_, new_n53720_, new_n53721_, new_n53722_, new_n53723_,
    new_n53724_, new_n53725_, new_n53726_, new_n53727_, new_n53728_,
    new_n53729_, new_n53730_, new_n53731_, new_n53732_, new_n53733_,
    new_n53734_, new_n53735_, new_n53736_, new_n53737_, new_n53738_,
    new_n53739_, new_n53740_, new_n53741_, new_n53742_, new_n53743_,
    new_n53744_, new_n53745_, new_n53746_, new_n53747_, new_n53748_,
    new_n53749_, new_n53750_, new_n53751_, new_n53752_, new_n53753_,
    new_n53754_, new_n53755_, new_n53756_, new_n53757_, new_n53758_,
    new_n53759_, new_n53760_, new_n53761_, new_n53762_, new_n53763_,
    new_n53764_, new_n53765_, new_n53766_, new_n53767_, new_n53768_,
    new_n53769_, new_n53770_, new_n53771_, new_n53772_, new_n53773_,
    new_n53774_, new_n53775_, new_n53776_, new_n53777_, new_n53778_,
    new_n53779_, new_n53780_, new_n53781_, new_n53782_, new_n53783_,
    new_n53784_, new_n53785_, new_n53786_, new_n53787_, new_n53788_,
    new_n53789_, new_n53790_, new_n53791_, new_n53792_, new_n53793_,
    new_n53794_, new_n53795_, new_n53796_, new_n53797_, new_n53798_,
    new_n53799_, new_n53800_, new_n53801_, new_n53802_, new_n53803_,
    new_n53804_, new_n53805_, new_n53806_, new_n53807_, new_n53808_,
    new_n53809_, new_n53810_, new_n53811_, new_n53812_, new_n53813_,
    new_n53814_, new_n53815_, new_n53816_, new_n53817_, new_n53818_,
    new_n53819_, new_n53820_, new_n53821_, new_n53822_, new_n53823_,
    new_n53824_, new_n53825_, new_n53826_, new_n53827_, new_n53828_,
    new_n53829_, new_n53830_, new_n53831_, new_n53832_, new_n53833_,
    new_n53834_, new_n53835_, new_n53836_, new_n53837_, new_n53838_,
    new_n53839_, new_n53840_, new_n53841_, new_n53842_, new_n53843_,
    new_n53844_, new_n53845_, new_n53846_, new_n53847_, new_n53848_,
    new_n53849_, new_n53850_, new_n53851_, new_n53852_, new_n53853_,
    new_n53854_, new_n53855_, new_n53856_, new_n53857_, new_n53858_,
    new_n53859_, new_n53860_, new_n53861_, new_n53862_, new_n53863_,
    new_n53864_, new_n53865_, new_n53866_, new_n53867_, new_n53868_,
    new_n53869_, new_n53870_, new_n53871_, new_n53872_, new_n53873_,
    new_n53874_, new_n53875_, new_n53876_, new_n53877_, new_n53878_,
    new_n53879_, new_n53880_, new_n53881_, new_n53882_, new_n53883_,
    new_n53884_, new_n53885_, new_n53886_, new_n53887_, new_n53888_,
    new_n53889_, new_n53890_, new_n53891_, new_n53892_, new_n53893_,
    new_n53894_, new_n53895_, new_n53896_, new_n53897_, new_n53898_,
    new_n53899_, new_n53900_, new_n53901_, new_n53902_, new_n53903_,
    new_n53904_, new_n53905_, new_n53906_, new_n53907_, new_n53908_,
    new_n53909_, new_n53910_, new_n53911_, new_n53912_, new_n53913_,
    new_n53914_, new_n53915_, new_n53916_, new_n53917_, new_n53918_,
    new_n53919_, new_n53920_, new_n53921_, new_n53922_, new_n53923_,
    new_n53924_, new_n53925_, new_n53926_, new_n53927_, new_n53928_,
    new_n53929_, new_n53930_, new_n53931_, new_n53932_, new_n53933_,
    new_n53934_, new_n53935_, new_n53936_, new_n53937_, new_n53938_,
    new_n53939_, new_n53940_, new_n53941_, new_n53942_, new_n53943_,
    new_n53944_, new_n53945_, new_n53946_, new_n53947_, new_n53948_,
    new_n53949_, new_n53950_, new_n53951_, new_n53952_, new_n53953_,
    new_n53954_, new_n53955_, new_n53956_, new_n53957_, new_n53958_,
    new_n53959_, new_n53960_, new_n53961_, new_n53962_, new_n53963_,
    new_n53964_, new_n53965_, new_n53966_, new_n53967_, new_n53968_,
    new_n53969_, new_n53970_, new_n53971_, new_n53972_, new_n53973_,
    new_n53974_, new_n53975_, new_n53976_, new_n53977_, new_n53978_,
    new_n53979_, new_n53980_, new_n53981_, new_n53982_, new_n53983_,
    new_n53984_, new_n53985_, new_n53986_, new_n53987_, new_n53988_,
    new_n53989_, new_n53990_, new_n53991_, new_n53992_, new_n53993_,
    new_n53994_, new_n53995_, new_n53996_, new_n53997_, new_n53998_,
    new_n53999_, new_n54000_, new_n54001_, new_n54002_, new_n54003_,
    new_n54004_, new_n54005_, new_n54006_, new_n54007_, new_n54008_,
    new_n54009_, new_n54010_, new_n54011_, new_n54012_, new_n54013_,
    new_n54014_, new_n54015_, new_n54016_, new_n54017_, new_n54018_,
    new_n54019_, new_n54020_, new_n54021_, new_n54022_, new_n54023_,
    new_n54024_, new_n54025_, new_n54026_, new_n54027_, new_n54028_,
    new_n54029_, new_n54030_, new_n54031_, new_n54032_, new_n54033_,
    new_n54034_, new_n54035_, new_n54036_, new_n54037_, new_n54038_,
    new_n54039_, new_n54040_, new_n54041_, new_n54042_, new_n54043_,
    new_n54044_, new_n54045_, new_n54046_, new_n54047_, new_n54048_,
    new_n54049_, new_n54050_, new_n54051_, new_n54052_, new_n54053_,
    new_n54054_, new_n54055_, new_n54056_, new_n54057_, new_n54058_,
    new_n54059_, new_n54060_, new_n54061_, new_n54062_, new_n54063_,
    new_n54064_, new_n54065_, new_n54066_, new_n54067_, new_n54068_,
    new_n54069_, new_n54070_, new_n54071_, new_n54072_, new_n54073_,
    new_n54074_, new_n54075_, new_n54076_, new_n54077_, new_n54078_,
    new_n54079_, new_n54080_, new_n54081_, new_n54082_, new_n54083_,
    new_n54084_, new_n54085_, new_n54086_, new_n54087_, new_n54088_,
    new_n54089_, new_n54090_, new_n54091_, new_n54092_, new_n54093_,
    new_n54094_, new_n54095_, new_n54096_, new_n54097_, new_n54098_,
    new_n54099_, new_n54100_, new_n54101_, new_n54102_, new_n54103_,
    new_n54104_, new_n54105_, new_n54106_, new_n54107_, new_n54108_,
    new_n54109_, new_n54110_, new_n54111_, new_n54112_, new_n54113_,
    new_n54114_, new_n54115_, new_n54116_, new_n54117_, new_n54118_,
    new_n54119_, new_n54120_, new_n54121_, new_n54122_, new_n54123_,
    new_n54124_, new_n54125_, new_n54126_, new_n54127_, new_n54128_,
    new_n54129_, new_n54130_, new_n54131_, new_n54132_, new_n54133_,
    new_n54134_, new_n54135_, new_n54136_, new_n54137_, new_n54138_,
    new_n54139_, new_n54140_, new_n54141_, new_n54142_, new_n54143_,
    new_n54144_, new_n54145_, new_n54146_, new_n54147_, new_n54148_,
    new_n54149_, new_n54150_, new_n54151_, new_n54152_, new_n54153_,
    new_n54154_, new_n54155_, new_n54156_, new_n54157_, new_n54158_,
    new_n54159_, new_n54160_, new_n54161_, new_n54162_, new_n54163_,
    new_n54164_, new_n54165_, new_n54166_, new_n54167_, new_n54168_,
    new_n54169_, new_n54170_, new_n54171_, new_n54172_, new_n54173_,
    new_n54174_, new_n54175_, new_n54176_, new_n54177_, new_n54178_,
    new_n54179_, new_n54180_, new_n54181_, new_n54182_, new_n54183_,
    new_n54184_, new_n54185_, new_n54186_, new_n54187_, new_n54188_,
    new_n54189_, new_n54190_, new_n54191_, new_n54192_, new_n54193_,
    new_n54194_, new_n54195_, new_n54196_, new_n54197_, new_n54198_,
    new_n54199_, new_n54200_, new_n54201_, new_n54202_, new_n54203_,
    new_n54204_, new_n54205_, new_n54206_, new_n54207_, new_n54208_,
    new_n54209_, new_n54210_, new_n54211_, new_n54212_, new_n54213_,
    new_n54214_, new_n54215_, new_n54216_, new_n54217_, new_n54218_,
    new_n54219_, new_n54220_, new_n54221_, new_n54222_, new_n54223_,
    new_n54224_, new_n54225_, new_n54226_, new_n54227_, new_n54228_,
    new_n54229_, new_n54230_, new_n54231_, new_n54232_, new_n54233_,
    new_n54234_, new_n54235_, new_n54236_, new_n54237_, new_n54238_,
    new_n54239_, new_n54240_, new_n54241_, new_n54242_, new_n54243_,
    new_n54244_, new_n54245_, new_n54246_, new_n54247_, new_n54248_,
    new_n54249_, new_n54250_, new_n54251_, new_n54252_, new_n54253_,
    new_n54254_, new_n54255_, new_n54256_, new_n54257_, new_n54258_,
    new_n54259_, new_n54260_, new_n54261_, new_n54262_, new_n54263_,
    new_n54264_, new_n54265_, new_n54266_, new_n54267_, new_n54268_,
    new_n54269_, new_n54270_, new_n54271_, new_n54272_, new_n54273_,
    new_n54274_, new_n54275_, new_n54276_, new_n54277_, new_n54278_,
    new_n54279_, new_n54280_, new_n54281_, new_n54282_, new_n54283_,
    new_n54284_, new_n54285_, new_n54286_, new_n54287_, new_n54288_,
    new_n54289_, new_n54290_, new_n54291_, new_n54292_, new_n54293_,
    new_n54294_, new_n54295_, new_n54296_, new_n54297_, new_n54298_,
    new_n54299_, new_n54300_, new_n54301_, new_n54302_, new_n54303_,
    new_n54304_, new_n54305_, new_n54306_, new_n54307_, new_n54308_,
    new_n54309_, new_n54310_, new_n54311_, new_n54312_, new_n54313_,
    new_n54314_, new_n54315_, new_n54316_, new_n54317_, new_n54318_,
    new_n54319_, new_n54320_, new_n54321_, new_n54322_, new_n54323_,
    new_n54324_, new_n54325_, new_n54326_, new_n54327_, new_n54328_,
    new_n54329_, new_n54330_, new_n54331_, new_n54332_, new_n54333_,
    new_n54334_, new_n54335_, new_n54336_, new_n54337_, new_n54338_,
    new_n54339_, new_n54340_, new_n54341_, new_n54342_, new_n54343_,
    new_n54344_, new_n54345_, new_n54346_, new_n54347_, new_n54348_,
    new_n54349_, new_n54350_, new_n54351_, new_n54352_, new_n54353_,
    new_n54354_, new_n54355_, new_n54356_, new_n54357_, new_n54358_,
    new_n54359_, new_n54360_, new_n54361_, new_n54362_, new_n54363_,
    new_n54364_, new_n54365_, new_n54366_, new_n54367_, new_n54368_,
    new_n54369_, new_n54370_, new_n54371_, new_n54372_, new_n54373_,
    new_n54374_, new_n54375_, new_n54376_, new_n54377_, new_n54378_,
    new_n54379_, new_n54380_, new_n54381_, new_n54382_, new_n54383_,
    new_n54384_, new_n54385_, new_n54386_, new_n54387_, new_n54388_,
    new_n54389_, new_n54390_, new_n54391_, new_n54392_, new_n54393_,
    new_n54394_, new_n54395_, new_n54396_, new_n54397_, new_n54398_,
    new_n54399_, new_n54400_, new_n54401_, new_n54402_, new_n54403_,
    new_n54404_, new_n54405_, new_n54406_, new_n54407_, new_n54408_,
    new_n54409_, new_n54410_, new_n54411_, new_n54412_, new_n54413_,
    new_n54414_, new_n54415_, new_n54416_, new_n54417_, new_n54418_,
    new_n54419_, new_n54420_, new_n54421_, new_n54422_, new_n54423_,
    new_n54424_, new_n54425_, new_n54426_, new_n54427_, new_n54428_,
    new_n54429_, new_n54430_, new_n54431_, new_n54432_, new_n54433_,
    new_n54434_, new_n54435_, new_n54436_, new_n54437_, new_n54438_,
    new_n54439_, new_n54440_, new_n54441_, new_n54442_, new_n54443_,
    new_n54444_, new_n54445_, new_n54446_, new_n54447_, new_n54448_,
    new_n54449_, new_n54450_, new_n54451_, new_n54452_, new_n54453_,
    new_n54454_, new_n54455_, new_n54456_, new_n54457_, new_n54458_,
    new_n54459_, new_n54460_, new_n54461_, new_n54462_, new_n54463_,
    new_n54464_, new_n54465_, new_n54466_, new_n54467_, new_n54468_,
    new_n54469_, new_n54470_, new_n54471_, new_n54472_, new_n54473_,
    new_n54474_, new_n54475_, new_n54476_, new_n54477_, new_n54478_,
    new_n54479_, new_n54480_, new_n54481_, new_n54482_, new_n54483_,
    new_n54484_, new_n54485_, new_n54486_, new_n54487_, new_n54488_,
    new_n54489_, new_n54490_, new_n54491_, new_n54492_, new_n54493_,
    new_n54494_, new_n54495_, new_n54496_, new_n54497_, new_n54498_,
    new_n54499_, new_n54500_, new_n54501_, new_n54502_, new_n54503_,
    new_n54504_, new_n54505_, new_n54506_, new_n54507_, new_n54508_,
    new_n54509_, new_n54510_, new_n54511_, new_n54512_, new_n54513_,
    new_n54514_, new_n54515_, new_n54516_, new_n54517_, new_n54518_,
    new_n54519_, new_n54520_, new_n54521_, new_n54522_, new_n54523_,
    new_n54524_, new_n54525_, new_n54526_, new_n54527_, new_n54528_,
    new_n54529_, new_n54530_, new_n54531_, new_n54532_, new_n54533_,
    new_n54534_, new_n54535_, new_n54536_, new_n54537_, new_n54538_,
    new_n54539_, new_n54540_, new_n54541_, new_n54542_, new_n54543_,
    new_n54544_, new_n54545_, new_n54546_, new_n54547_, new_n54548_,
    new_n54549_, new_n54550_, new_n54551_, new_n54552_, new_n54553_,
    new_n54554_, new_n54555_, new_n54556_, new_n54557_, new_n54558_,
    new_n54559_, new_n54560_, new_n54561_, new_n54562_, new_n54563_,
    new_n54564_, new_n54565_, new_n54566_, new_n54567_, new_n54568_,
    new_n54569_, new_n54570_, new_n54571_, new_n54572_, new_n54573_,
    new_n54574_, new_n54575_, new_n54576_, new_n54577_, new_n54578_,
    new_n54579_, new_n54580_, new_n54581_, new_n54582_, new_n54583_,
    new_n54584_, new_n54585_, new_n54586_, new_n54587_, new_n54588_,
    new_n54589_, new_n54590_, new_n54591_, new_n54592_, new_n54593_,
    new_n54594_, new_n54595_, new_n54596_, new_n54597_, new_n54598_,
    new_n54599_, new_n54600_, new_n54601_, new_n54602_, new_n54603_,
    new_n54604_, new_n54605_, new_n54606_, new_n54607_, new_n54608_,
    new_n54609_, new_n54610_, new_n54611_, new_n54612_, new_n54613_,
    new_n54614_, new_n54615_, new_n54616_, new_n54617_, new_n54618_,
    new_n54619_, new_n54620_, new_n54621_, new_n54622_, new_n54623_,
    new_n54624_, new_n54625_, new_n54626_, new_n54627_, new_n54628_,
    new_n54629_, new_n54630_, new_n54631_, new_n54632_, new_n54633_,
    new_n54634_, new_n54635_, new_n54636_, new_n54637_, new_n54638_,
    new_n54639_, new_n54640_, new_n54641_, new_n54642_, new_n54643_,
    new_n54644_, new_n54645_, new_n54646_, new_n54647_, new_n54648_,
    new_n54649_, new_n54650_, new_n54651_, new_n54652_, new_n54653_,
    new_n54654_, new_n54655_, new_n54656_, new_n54657_, new_n54658_,
    new_n54659_, new_n54660_, new_n54661_, new_n54662_, new_n54663_,
    new_n54664_, new_n54665_, new_n54666_, new_n54667_, new_n54668_,
    new_n54669_, new_n54670_, new_n54671_, new_n54672_, new_n54673_,
    new_n54674_, new_n54675_, new_n54676_, new_n54677_, new_n54678_,
    new_n54679_, new_n54680_, new_n54681_, new_n54682_, new_n54683_,
    new_n54684_, new_n54685_, new_n54686_, new_n54687_, new_n54688_,
    new_n54689_, new_n54690_, new_n54691_, new_n54692_, new_n54693_,
    new_n54694_, new_n54695_, new_n54696_, new_n54697_, new_n54698_,
    new_n54699_, new_n54700_, new_n54701_, new_n54702_, new_n54703_,
    new_n54704_, new_n54705_, new_n54706_, new_n54707_, new_n54708_,
    new_n54709_, new_n54710_, new_n54711_, new_n54712_, new_n54713_,
    new_n54714_, new_n54715_, new_n54716_, new_n54717_, new_n54718_,
    new_n54719_, new_n54720_, new_n54721_, new_n54722_, new_n54723_,
    new_n54724_, new_n54725_, new_n54726_, new_n54727_, new_n54728_,
    new_n54729_, new_n54730_, new_n54731_, new_n54732_, new_n54733_,
    new_n54734_, new_n54735_, new_n54736_, new_n54737_, new_n54738_,
    new_n54739_, new_n54740_, new_n54741_, new_n54742_, new_n54743_,
    new_n54744_, new_n54745_, new_n54746_, new_n54747_, new_n54748_,
    new_n54749_, new_n54750_, new_n54751_, new_n54752_, new_n54753_,
    new_n54754_, new_n54755_, new_n54756_, new_n54757_, new_n54758_,
    new_n54759_, new_n54760_, new_n54761_, new_n54762_, new_n54763_,
    new_n54764_, new_n54765_, new_n54766_, new_n54767_, new_n54768_,
    new_n54769_, new_n54770_, new_n54771_, new_n54772_, new_n54773_,
    new_n54774_, new_n54775_, new_n54776_, new_n54777_, new_n54778_,
    new_n54779_, new_n54780_, new_n54781_, new_n54782_, new_n54783_,
    new_n54784_, new_n54785_, new_n54786_, new_n54787_, new_n54788_,
    new_n54789_, new_n54790_, new_n54791_, new_n54792_, new_n54793_,
    new_n54794_, new_n54795_, new_n54796_, new_n54797_, new_n54798_,
    new_n54799_, new_n54800_, new_n54801_, new_n54802_, new_n54803_,
    new_n54804_, new_n54805_, new_n54806_, new_n54807_, new_n54808_,
    new_n54809_, new_n54810_, new_n54811_, new_n54812_, new_n54813_,
    new_n54814_, new_n54815_, new_n54816_, new_n54817_, new_n54818_,
    new_n54819_, new_n54820_, new_n54821_, new_n54822_, new_n54823_,
    new_n54824_, new_n54825_, new_n54826_, new_n54827_, new_n54828_,
    new_n54829_, new_n54830_, new_n54831_, new_n54832_, new_n54833_,
    new_n54834_, new_n54835_, new_n54836_, new_n54837_, new_n54838_,
    new_n54839_, new_n54840_, new_n54841_, new_n54842_, new_n54843_,
    new_n54844_, new_n54845_, new_n54846_, new_n54847_, new_n54848_,
    new_n54849_, new_n54850_, new_n54851_, new_n54852_, new_n54853_,
    new_n54854_, new_n54855_, new_n54856_, new_n54857_, new_n54858_,
    new_n54859_, new_n54860_, new_n54861_, new_n54862_, new_n54863_,
    new_n54864_, new_n54865_, new_n54866_, new_n54867_, new_n54868_,
    new_n54869_, new_n54870_, new_n54871_, new_n54872_, new_n54873_,
    new_n54874_, new_n54875_, new_n54876_, new_n54877_, new_n54878_,
    new_n54879_, new_n54880_, new_n54881_, new_n54882_, new_n54883_,
    new_n54884_, new_n54885_, new_n54886_, new_n54887_, new_n54888_,
    new_n54889_, new_n54890_, new_n54891_, new_n54892_, new_n54893_,
    new_n54894_, new_n54895_, new_n54896_, new_n54897_, new_n54898_,
    new_n54899_, new_n54900_, new_n54901_, new_n54902_, new_n54903_,
    new_n54904_, new_n54905_, new_n54906_, new_n54907_, new_n54908_,
    new_n54909_, new_n54910_, new_n54911_, new_n54912_, new_n54913_,
    new_n54914_, new_n54915_, new_n54916_, new_n54917_, new_n54918_,
    new_n54919_, new_n54920_, new_n54921_, new_n54922_, new_n54923_,
    new_n54924_, new_n54925_, new_n54926_, new_n54927_, new_n54928_,
    new_n54929_, new_n54930_, new_n54931_, new_n54932_, new_n54933_,
    new_n54934_, new_n54935_, new_n54936_, new_n54937_, new_n54938_,
    new_n54939_, new_n54940_, new_n54941_, new_n54942_, new_n54943_,
    new_n54944_, new_n54945_, new_n54946_, new_n54947_, new_n54948_,
    new_n54949_, new_n54950_, new_n54951_, new_n54952_, new_n54953_,
    new_n54954_, new_n54955_, new_n54956_, new_n54957_, new_n54958_,
    new_n54959_, new_n54960_, new_n54961_, new_n54962_, new_n54963_,
    new_n54964_, new_n54965_, new_n54966_, new_n54967_, new_n54968_,
    new_n54969_, new_n54970_, new_n54971_, new_n54972_, new_n54973_,
    new_n54974_, new_n54975_, new_n54976_, new_n54977_, new_n54978_,
    new_n54979_, new_n54980_, new_n54981_, new_n54982_, new_n54983_,
    new_n54984_, new_n54985_, new_n54986_, new_n54987_, new_n54988_,
    new_n54989_, new_n54990_, new_n54991_, new_n54992_, new_n54993_,
    new_n54994_, new_n54995_, new_n54996_, new_n54997_, new_n54998_,
    new_n54999_, new_n55000_, new_n55001_, new_n55002_, new_n55003_,
    new_n55004_, new_n55005_, new_n55006_, new_n55007_, new_n55008_,
    new_n55009_, new_n55010_, new_n55011_, new_n55012_, new_n55013_,
    new_n55014_, new_n55015_, new_n55016_, new_n55017_, new_n55018_,
    new_n55019_, new_n55020_, new_n55021_, new_n55022_, new_n55023_,
    new_n55024_, new_n55025_, new_n55026_, new_n55027_, new_n55028_,
    new_n55029_, new_n55030_, new_n55031_, new_n55032_, new_n55033_,
    new_n55034_, new_n55035_, new_n55036_, new_n55037_, new_n55038_,
    new_n55039_, new_n55040_, new_n55041_, new_n55042_, new_n55043_,
    new_n55044_, new_n55045_, new_n55046_, new_n55047_, new_n55048_,
    new_n55049_, new_n55050_, new_n55051_, new_n55052_, new_n55053_,
    new_n55054_, new_n55055_, new_n55056_, new_n55057_, new_n55058_,
    new_n55059_, new_n55060_, new_n55061_, new_n55062_, new_n55063_,
    new_n55064_, new_n55065_, new_n55066_, new_n55067_, new_n55068_,
    new_n55069_, new_n55070_, new_n55071_, new_n55072_, new_n55073_,
    new_n55074_, new_n55075_, new_n55076_, new_n55077_, new_n55078_,
    new_n55079_, new_n55080_, new_n55081_, new_n55082_, new_n55083_,
    new_n55084_, new_n55085_, new_n55086_, new_n55087_, new_n55088_,
    new_n55089_, new_n55090_, new_n55091_, new_n55092_, new_n55093_,
    new_n55094_, new_n55095_, new_n55096_, new_n55097_, new_n55098_,
    new_n55099_, new_n55100_, new_n55101_, new_n55102_, new_n55103_,
    new_n55104_, new_n55105_, new_n55106_, new_n55107_, new_n55108_,
    new_n55109_, new_n55110_, new_n55111_, new_n55112_, new_n55113_,
    new_n55114_, new_n55115_, new_n55116_, new_n55117_, new_n55118_,
    new_n55119_, new_n55120_, new_n55121_, new_n55122_, new_n55123_,
    new_n55124_, new_n55125_, new_n55126_, new_n55127_, new_n55128_,
    new_n55129_, new_n55130_, new_n55131_, new_n55132_, new_n55133_,
    new_n55134_, new_n55135_, new_n55136_, new_n55137_, new_n55138_,
    new_n55139_, new_n55140_, new_n55141_, new_n55142_, new_n55143_,
    new_n55144_, new_n55145_, new_n55146_, new_n55147_, new_n55148_,
    new_n55149_, new_n55150_, new_n55151_, new_n55152_, new_n55153_,
    new_n55154_, new_n55155_, new_n55156_, new_n55157_, new_n55158_,
    new_n55159_, new_n55160_, new_n55161_, new_n55162_, new_n55163_,
    new_n55164_, new_n55165_, new_n55166_, new_n55167_, new_n55168_,
    new_n55169_, new_n55170_, new_n55171_, new_n55172_, new_n55173_,
    new_n55174_, new_n55175_, new_n55176_, new_n55177_, new_n55178_,
    new_n55179_, new_n55180_, new_n55181_, new_n55182_, new_n55183_,
    new_n55184_, new_n55185_, new_n55186_, new_n55187_, new_n55188_,
    new_n55189_, new_n55190_, new_n55191_, new_n55192_, new_n55193_,
    new_n55194_, new_n55195_, new_n55196_, new_n55197_, new_n55198_,
    new_n55199_, new_n55200_, new_n55201_, new_n55202_, new_n55203_,
    new_n55204_, new_n55205_, new_n55206_, new_n55207_, new_n55208_,
    new_n55209_, new_n55210_, new_n55211_, new_n55212_, new_n55213_,
    new_n55214_, new_n55215_, new_n55216_, new_n55217_, new_n55218_,
    new_n55219_, new_n55220_, new_n55221_, new_n55222_, new_n55223_,
    new_n55224_, new_n55225_, new_n55226_, new_n55227_, new_n55228_,
    new_n55229_, new_n55230_, new_n55231_, new_n55232_, new_n55233_,
    new_n55234_, new_n55235_, new_n55236_, new_n55237_, new_n55238_,
    new_n55239_, new_n55240_, new_n55241_, new_n55242_, new_n55243_,
    new_n55244_, new_n55245_, new_n55246_, new_n55247_, new_n55248_,
    new_n55249_, new_n55250_, new_n55251_, new_n55252_, new_n55253_,
    new_n55254_, new_n55255_, new_n55256_, new_n55257_, new_n55258_,
    new_n55259_, new_n55260_, new_n55261_, new_n55262_, new_n55263_,
    new_n55264_, new_n55265_, new_n55266_, new_n55267_, new_n55268_,
    new_n55269_, new_n55270_, new_n55271_, new_n55272_, new_n55273_,
    new_n55274_, new_n55275_, new_n55276_, new_n55277_, new_n55278_,
    new_n55279_, new_n55280_, new_n55281_, new_n55282_, new_n55283_,
    new_n55284_, new_n55285_, new_n55286_, new_n55287_, new_n55288_,
    new_n55289_, new_n55290_, new_n55291_, new_n55292_, new_n55293_,
    new_n55294_, new_n55295_, new_n55296_, new_n55297_, new_n55298_,
    new_n55299_, new_n55300_, new_n55301_, new_n55302_, new_n55303_,
    new_n55304_, new_n55305_, new_n55306_, new_n55307_, new_n55308_,
    new_n55309_, new_n55310_, new_n55311_, new_n55312_, new_n55313_,
    new_n55314_, new_n55315_, new_n55316_, new_n55317_, new_n55318_,
    new_n55319_, new_n55320_, new_n55321_, new_n55322_, new_n55323_,
    new_n55324_, new_n55325_, new_n55326_, new_n55327_, new_n55328_,
    new_n55329_, new_n55330_, new_n55331_, new_n55332_, new_n55333_,
    new_n55334_, new_n55335_, new_n55336_, new_n55337_, new_n55338_,
    new_n55339_, new_n55340_, new_n55341_, new_n55342_, new_n55343_,
    new_n55344_, new_n55345_, new_n55346_, new_n55347_, new_n55348_,
    new_n55349_, new_n55350_, new_n55351_, new_n55352_, new_n55353_,
    new_n55354_, new_n55355_, new_n55356_, new_n55357_, new_n55358_,
    new_n55359_, new_n55360_, new_n55361_, new_n55362_, new_n55363_,
    new_n55364_, new_n55365_, new_n55366_, new_n55367_, new_n55368_,
    new_n55369_, new_n55370_, new_n55371_, new_n55372_, new_n55373_,
    new_n55374_, new_n55375_, new_n55376_, new_n55377_, new_n55378_,
    new_n55379_, new_n55380_, new_n55381_, new_n55382_, new_n55383_,
    new_n55384_, new_n55385_, new_n55386_, new_n55387_, new_n55388_,
    new_n55389_, new_n55390_, new_n55391_, new_n55392_, new_n55393_,
    new_n55394_, new_n55395_, new_n55396_, new_n55397_, new_n55398_,
    new_n55399_, new_n55400_, new_n55401_, new_n55402_, new_n55403_,
    new_n55404_, new_n55405_, new_n55406_, new_n55407_, new_n55408_,
    new_n55409_, new_n55410_, new_n55411_, new_n55412_, new_n55413_,
    new_n55414_, new_n55415_, new_n55416_, new_n55417_, new_n55418_,
    new_n55419_, new_n55420_, new_n55421_, new_n55422_, new_n55423_,
    new_n55424_, new_n55425_, new_n55426_, new_n55427_, new_n55428_,
    new_n55429_, new_n55430_, new_n55431_, new_n55432_, new_n55433_,
    new_n55434_, new_n55435_, new_n55436_, new_n55437_, new_n55438_,
    new_n55439_, new_n55440_, new_n55441_, new_n55442_, new_n55443_,
    new_n55444_, new_n55445_, new_n55446_, new_n55447_, new_n55448_,
    new_n55449_, new_n55450_, new_n55451_, new_n55452_, new_n55453_,
    new_n55454_, new_n55455_, new_n55456_, new_n55457_, new_n55458_,
    new_n55459_, new_n55460_, new_n55461_, new_n55462_, new_n55463_,
    new_n55464_, new_n55465_, new_n55466_, new_n55467_, new_n55468_,
    new_n55469_, new_n55470_, new_n55471_, new_n55472_, new_n55473_,
    new_n55474_, new_n55475_, new_n55476_, new_n55477_, new_n55478_,
    new_n55479_, new_n55480_, new_n55481_, new_n55482_, new_n55483_,
    new_n55484_, new_n55485_, new_n55486_, new_n55487_, new_n55488_,
    new_n55489_, new_n55490_, new_n55491_, new_n55492_, new_n55493_,
    new_n55494_, new_n55495_, new_n55496_, new_n55497_, new_n55498_,
    new_n55499_, new_n55500_, new_n55501_, new_n55502_, new_n55503_,
    new_n55504_, new_n55505_, new_n55506_, new_n55507_, new_n55508_,
    new_n55509_, new_n55510_, new_n55511_, new_n55512_, new_n55513_,
    new_n55514_, new_n55515_, new_n55516_, new_n55517_, new_n55518_,
    new_n55519_, new_n55520_, new_n55521_, new_n55522_, new_n55523_,
    new_n55524_, new_n55525_, new_n55526_, new_n55527_, new_n55528_,
    new_n55529_, new_n55530_, new_n55531_, new_n55532_, new_n55533_,
    new_n55534_, new_n55535_, new_n55536_, new_n55537_, new_n55538_,
    new_n55539_, new_n55540_, new_n55541_, new_n55542_, new_n55543_,
    new_n55544_, new_n55545_, new_n55546_, new_n55547_, new_n55548_,
    new_n55549_, new_n55550_, new_n55551_, new_n55552_, new_n55553_,
    new_n55554_, new_n55555_, new_n55556_, new_n55557_, new_n55558_,
    new_n55559_, new_n55560_, new_n55561_, new_n55562_, new_n55563_,
    new_n55564_, new_n55565_, new_n55566_, new_n55567_, new_n55568_,
    new_n55569_, new_n55570_, new_n55571_, new_n55572_, new_n55573_,
    new_n55574_, new_n55575_, new_n55576_, new_n55577_, new_n55578_,
    new_n55579_, new_n55580_, new_n55581_, new_n55582_, new_n55583_,
    new_n55584_, new_n55585_, new_n55586_, new_n55587_, new_n55588_,
    new_n55589_, new_n55590_, new_n55591_, new_n55592_, new_n55593_,
    new_n55594_, new_n55595_, new_n55596_, new_n55597_, new_n55598_,
    new_n55599_, new_n55600_, new_n55601_, new_n55602_, new_n55603_,
    new_n55604_, new_n55605_, new_n55606_, new_n55607_, new_n55608_,
    new_n55609_, new_n55610_, new_n55611_, new_n55612_, new_n55613_,
    new_n55614_, new_n55615_, new_n55616_, new_n55617_, new_n55618_,
    new_n55619_, new_n55620_, new_n55621_, new_n55622_, new_n55623_,
    new_n55624_, new_n55625_, new_n55626_, new_n55627_, new_n55628_,
    new_n55629_, new_n55630_, new_n55631_, new_n55632_, new_n55633_,
    new_n55634_, new_n55635_, new_n55636_, new_n55637_, new_n55638_,
    new_n55639_, new_n55640_, new_n55641_, new_n55642_, new_n55643_,
    new_n55644_, new_n55645_, new_n55646_, new_n55647_, new_n55648_,
    new_n55649_, new_n55650_, new_n55651_, new_n55652_, new_n55653_,
    new_n55654_, new_n55655_, new_n55656_, new_n55657_, new_n55658_,
    new_n55659_, new_n55660_, new_n55661_, new_n55662_, new_n55663_,
    new_n55664_, new_n55665_, new_n55666_, new_n55667_, new_n55668_,
    new_n55669_, new_n55670_, new_n55671_, new_n55672_, new_n55673_,
    new_n55674_, new_n55675_, new_n55676_, new_n55677_, new_n55678_,
    new_n55679_, new_n55680_, new_n55681_, new_n55682_, new_n55683_,
    new_n55684_, new_n55685_, new_n55686_, new_n55687_, new_n55688_,
    new_n55689_, new_n55690_, new_n55691_, new_n55692_, new_n55693_,
    new_n55694_, new_n55695_, new_n55696_, new_n55697_, new_n55698_,
    new_n55699_, new_n55700_, new_n55701_, new_n55702_, new_n55703_,
    new_n55704_, new_n55705_, new_n55706_, new_n55707_, new_n55708_,
    new_n55709_, new_n55710_, new_n55711_, new_n55712_, new_n55713_,
    new_n55714_, new_n55715_, new_n55716_, new_n55717_, new_n55718_,
    new_n55719_, new_n55720_, new_n55721_, new_n55722_, new_n55723_,
    new_n55724_, new_n55725_, new_n55726_, new_n55727_, new_n55728_,
    new_n55729_, new_n55730_, new_n55731_, new_n55732_, new_n55733_,
    new_n55734_, new_n55735_, new_n55736_, new_n55737_, new_n55738_,
    new_n55739_, new_n55740_, new_n55741_, new_n55742_, new_n55743_,
    new_n55744_, new_n55745_, new_n55746_, new_n55747_, new_n55748_,
    new_n55749_, new_n55750_, new_n55751_, new_n55752_, new_n55753_,
    new_n55754_, new_n55755_, new_n55756_, new_n55757_, new_n55758_,
    new_n55759_, new_n55760_, new_n55761_, new_n55762_, new_n55763_,
    new_n55764_, new_n55765_, new_n55766_, new_n55767_, new_n55768_,
    new_n55769_, new_n55770_, new_n55771_, new_n55772_, new_n55773_,
    new_n55774_, new_n55775_, new_n55776_, new_n55777_, new_n55778_,
    new_n55779_, new_n55780_, new_n55781_, new_n55782_, new_n55783_,
    new_n55784_, new_n55785_, new_n55786_, new_n55787_, new_n55788_,
    new_n55789_, new_n55790_, new_n55791_, new_n55792_, new_n55793_,
    new_n55794_, new_n55795_, new_n55796_, new_n55797_, new_n55798_,
    new_n55799_, new_n55800_, new_n55801_, new_n55802_, new_n55803_,
    new_n55804_, new_n55805_, new_n55806_, new_n55807_, new_n55808_,
    new_n55809_, new_n55810_, new_n55811_, new_n55812_, new_n55813_,
    new_n55814_, new_n55815_, new_n55816_, new_n55817_, new_n55818_,
    new_n55819_, new_n55820_, new_n55821_, new_n55822_, new_n55823_,
    new_n55824_, new_n55825_, new_n55826_, new_n55827_, new_n55828_,
    new_n55829_, new_n55830_, new_n55831_, new_n55832_, new_n55833_,
    new_n55834_, new_n55835_, new_n55836_, new_n55837_, new_n55838_,
    new_n55839_, new_n55840_, new_n55841_, new_n55842_, new_n55843_,
    new_n55844_, new_n55845_, new_n55846_, new_n55847_, new_n55848_,
    new_n55849_, new_n55850_, new_n55851_, new_n55852_, new_n55853_,
    new_n55854_, new_n55855_, new_n55856_, new_n55857_, new_n55858_,
    new_n55859_, new_n55860_, new_n55861_, new_n55862_, new_n55863_,
    new_n55864_, new_n55865_, new_n55866_, new_n55867_, new_n55868_,
    new_n55869_, new_n55870_, new_n55871_, new_n55872_, new_n55873_,
    new_n55874_, new_n55875_, new_n55876_, new_n55877_, new_n55878_,
    new_n55879_, new_n55880_, new_n55881_, new_n55882_, new_n55883_,
    new_n55884_, new_n55885_, new_n55886_, new_n55887_, new_n55888_,
    new_n55889_, new_n55890_, new_n55891_, new_n55892_, new_n55893_,
    new_n55894_, new_n55895_, new_n55896_, new_n55897_, new_n55898_,
    new_n55899_, new_n55900_, new_n55901_, new_n55902_, new_n55903_,
    new_n55904_, new_n55905_, new_n55906_, new_n55907_, new_n55908_,
    new_n55909_, new_n55910_, new_n55911_, new_n55912_, new_n55913_,
    new_n55914_, new_n55915_, new_n55916_, new_n55917_, new_n55918_,
    new_n55919_, new_n55920_, new_n55921_, new_n55922_, new_n55923_,
    new_n55924_, new_n55925_, new_n55926_, new_n55927_, new_n55928_,
    new_n55929_, new_n55930_, new_n55931_, new_n55932_, new_n55933_,
    new_n55934_, new_n55935_, new_n55936_, new_n55937_, new_n55938_,
    new_n55939_, new_n55940_, new_n55941_, new_n55942_, new_n55943_,
    new_n55944_, new_n55945_, new_n55946_, new_n55947_, new_n55948_,
    new_n55949_, new_n55950_, new_n55951_, new_n55952_, new_n55953_,
    new_n55954_, new_n55955_, new_n55956_, new_n55957_, new_n55958_,
    new_n55959_, new_n55960_, new_n55961_, new_n55962_, new_n55963_,
    new_n55964_, new_n55965_, new_n55966_, new_n55967_, new_n55968_,
    new_n55969_, new_n55970_, new_n55971_, new_n55972_, new_n55973_,
    new_n55974_, new_n55975_, new_n55976_, new_n55977_, new_n55978_,
    new_n55979_, new_n55980_, new_n55981_, new_n55982_, new_n55983_,
    new_n55984_, new_n55985_, new_n55986_, new_n55987_, new_n55988_,
    new_n55989_, new_n55990_, new_n55991_, new_n55992_, new_n55993_,
    new_n55994_, new_n55995_, new_n55996_, new_n55997_, new_n55998_,
    new_n55999_, new_n56000_, new_n56001_, new_n56002_, new_n56003_,
    new_n56004_, new_n56005_, new_n56006_, new_n56007_, new_n56008_,
    new_n56009_, new_n56010_, new_n56011_, new_n56012_, new_n56013_,
    new_n56014_, new_n56015_, new_n56016_, new_n56017_, new_n56018_,
    new_n56019_, new_n56020_, new_n56021_, new_n56022_, new_n56023_,
    new_n56024_, new_n56025_, new_n56026_, new_n56027_, new_n56028_,
    new_n56029_, new_n56030_, new_n56031_, new_n56032_, new_n56033_,
    new_n56034_, new_n56035_, new_n56036_, new_n56037_, new_n56038_,
    new_n56039_, new_n56040_, new_n56041_, new_n56042_, new_n56043_,
    new_n56044_, new_n56045_, new_n56046_, new_n56047_, new_n56048_,
    new_n56049_, new_n56050_, new_n56051_, new_n56052_, new_n56053_,
    new_n56054_, new_n56055_, new_n56056_, new_n56057_, new_n56058_,
    new_n56059_, new_n56060_, new_n56061_, new_n56062_, new_n56063_,
    new_n56064_, new_n56065_, new_n56066_, new_n56067_, new_n56068_,
    new_n56069_, new_n56070_, new_n56071_, new_n56072_, new_n56073_,
    new_n56074_, new_n56075_, new_n56076_, new_n56077_, new_n56078_,
    new_n56079_, new_n56080_, new_n56081_, new_n56082_, new_n56083_,
    new_n56084_, new_n56085_, new_n56086_, new_n56087_, new_n56088_,
    new_n56089_, new_n56090_, new_n56091_, new_n56092_, new_n56093_,
    new_n56094_, new_n56095_, new_n56096_, new_n56097_, new_n56098_,
    new_n56099_, new_n56100_, new_n56101_, new_n56102_, new_n56103_,
    new_n56104_, new_n56105_, new_n56106_, new_n56107_, new_n56108_,
    new_n56109_, new_n56110_, new_n56111_, new_n56112_, new_n56113_,
    new_n56114_, new_n56115_, new_n56116_, new_n56117_, new_n56118_,
    new_n56119_, new_n56120_, new_n56121_, new_n56122_, new_n56123_,
    new_n56124_, new_n56125_, new_n56126_, new_n56127_, new_n56128_,
    new_n56129_, new_n56130_, new_n56131_, new_n56132_, new_n56133_,
    new_n56134_, new_n56135_, new_n56136_, new_n56137_, new_n56138_,
    new_n56139_, new_n56140_, new_n56141_, new_n56142_, new_n56143_,
    new_n56144_, new_n56145_, new_n56146_, new_n56147_, new_n56148_,
    new_n56149_, new_n56150_, new_n56151_, new_n56152_, new_n56153_,
    new_n56154_, new_n56155_, new_n56156_, new_n56157_, new_n56158_,
    new_n56159_, new_n56160_, new_n56161_, new_n56162_, new_n56163_,
    new_n56164_, new_n56165_, new_n56166_, new_n56167_, new_n56168_,
    new_n56169_, new_n56170_, new_n56171_, new_n56172_, new_n56173_,
    new_n56174_, new_n56175_, new_n56176_, new_n56177_, new_n56178_,
    new_n56179_, new_n56180_, new_n56181_, new_n56182_, new_n56183_,
    new_n56184_, new_n56185_, new_n56186_, new_n56187_, new_n56188_,
    new_n56189_, new_n56190_, new_n56191_, new_n56192_, new_n56193_,
    new_n56194_, new_n56195_, new_n56196_, new_n56197_, new_n56198_,
    new_n56199_, new_n56200_, new_n56201_, new_n56202_, new_n56203_,
    new_n56204_, new_n56205_, new_n56206_, new_n56207_, new_n56208_,
    new_n56209_, new_n56210_, new_n56211_, new_n56212_, new_n56213_,
    new_n56214_, new_n56215_, new_n56216_, new_n56217_, new_n56218_,
    new_n56219_, new_n56220_, new_n56221_, new_n56222_, new_n56223_,
    new_n56224_, new_n56225_, new_n56226_, new_n56227_, new_n56228_,
    new_n56229_, new_n56230_, new_n56231_, new_n56232_, new_n56233_,
    new_n56234_, new_n56235_, new_n56236_, new_n56237_, new_n56238_,
    new_n56239_, new_n56240_, new_n56241_, new_n56242_, new_n56243_,
    new_n56244_, new_n56245_, new_n56246_, new_n56247_, new_n56248_,
    new_n56249_, new_n56250_, new_n56251_, new_n56252_, new_n56253_,
    new_n56254_, new_n56255_, new_n56256_, new_n56257_, new_n56258_,
    new_n56259_, new_n56260_, new_n56261_, new_n56262_, new_n56263_,
    new_n56264_, new_n56265_, new_n56266_, new_n56267_, new_n56268_,
    new_n56269_, new_n56270_, new_n56271_, new_n56272_, new_n56273_,
    new_n56274_, new_n56275_, new_n56276_, new_n56277_, new_n56278_,
    new_n56279_, new_n56280_, new_n56281_, new_n56282_, new_n56283_,
    new_n56284_, new_n56285_, new_n56286_, new_n56287_, new_n56288_,
    new_n56289_, new_n56290_, new_n56291_, new_n56292_, new_n56293_,
    new_n56294_, new_n56295_, new_n56296_, new_n56297_, new_n56298_,
    new_n56299_, new_n56300_, new_n56301_, new_n56302_, new_n56303_,
    new_n56304_, new_n56305_, new_n56306_, new_n56307_, new_n56308_,
    new_n56309_, new_n56310_, new_n56311_, new_n56312_, new_n56313_,
    new_n56314_, new_n56315_, new_n56316_, new_n56317_, new_n56318_,
    new_n56319_, new_n56320_, new_n56321_, new_n56322_, new_n56323_,
    new_n56324_, new_n56325_, new_n56326_, new_n56327_, new_n56328_,
    new_n56329_, new_n56330_, new_n56331_, new_n56332_, new_n56333_,
    new_n56334_, new_n56335_, new_n56336_, new_n56337_, new_n56338_,
    new_n56339_, new_n56340_, new_n56341_, new_n56342_, new_n56343_,
    new_n56344_, new_n56345_, new_n56346_, new_n56347_, new_n56348_,
    new_n56349_, new_n56350_, new_n56351_, new_n56352_, new_n56353_,
    new_n56354_, new_n56355_, new_n56356_, new_n56357_, new_n56358_,
    new_n56359_, new_n56360_, new_n56361_, new_n56362_, new_n56363_,
    new_n56364_, new_n56365_, new_n56366_, new_n56367_, new_n56368_,
    new_n56369_, new_n56370_, new_n56371_, new_n56372_, new_n56373_,
    new_n56374_, new_n56375_, new_n56376_, new_n56377_, new_n56378_,
    new_n56379_, new_n56380_, new_n56381_, new_n56382_, new_n56383_,
    new_n56384_, new_n56385_, new_n56386_, new_n56387_, new_n56388_,
    new_n56389_, new_n56390_, new_n56391_, new_n56392_, new_n56393_,
    new_n56394_, new_n56395_, new_n56396_, new_n56397_, new_n56398_,
    new_n56399_, new_n56400_, new_n56401_, new_n56402_, new_n56403_,
    new_n56404_, new_n56405_, new_n56406_, new_n56407_, new_n56408_,
    new_n56409_, new_n56410_, new_n56411_, new_n56412_, new_n56413_,
    new_n56414_, new_n56415_, new_n56416_, new_n56417_, new_n56418_,
    new_n56419_, new_n56420_, new_n56421_, new_n56422_, new_n56423_,
    new_n56424_, new_n56425_, new_n56426_, new_n56427_, new_n56428_,
    new_n56429_, new_n56430_, new_n56431_, new_n56432_, new_n56433_,
    new_n56434_, new_n56435_, new_n56436_, new_n56437_, new_n56438_,
    new_n56439_, new_n56440_, new_n56441_, new_n56442_, new_n56443_,
    new_n56444_, new_n56445_, new_n56446_, new_n56447_, new_n56448_,
    new_n56449_, new_n56450_, new_n56451_, new_n56452_, new_n56453_,
    new_n56454_, new_n56455_, new_n56456_, new_n56457_, new_n56458_,
    new_n56459_, new_n56460_, new_n56461_, new_n56462_, new_n56463_,
    new_n56464_, new_n56465_, new_n56466_, new_n56467_, new_n56468_,
    new_n56469_, new_n56470_, new_n56471_, new_n56472_, new_n56473_,
    new_n56474_, new_n56475_, new_n56476_, new_n56477_, new_n56478_,
    new_n56479_, new_n56480_, new_n56481_, new_n56482_, new_n56483_,
    new_n56484_, new_n56485_, new_n56486_, new_n56487_, new_n56488_,
    new_n56489_, new_n56490_, new_n56491_, new_n56492_, new_n56493_,
    new_n56494_, new_n56495_, new_n56496_, new_n56497_, new_n56498_,
    new_n56499_, new_n56500_, new_n56501_, new_n56502_, new_n56503_,
    new_n56504_, new_n56505_, new_n56506_, new_n56507_, new_n56508_,
    new_n56509_, new_n56510_, new_n56511_, new_n56512_, new_n56513_,
    new_n56514_, new_n56515_, new_n56516_, new_n56517_, new_n56518_,
    new_n56519_, new_n56520_, new_n56521_, new_n56522_, new_n56523_,
    new_n56524_, new_n56525_, new_n56526_, new_n56527_, new_n56528_,
    new_n56529_, new_n56530_, new_n56531_, new_n56532_, new_n56533_,
    new_n56534_, new_n56535_, new_n56536_, new_n56537_, new_n56538_,
    new_n56539_, new_n56540_, new_n56541_, new_n56542_, new_n56543_,
    new_n56544_, new_n56545_, new_n56546_, new_n56547_, new_n56548_,
    new_n56549_, new_n56550_, new_n56551_, new_n56552_, new_n56553_,
    new_n56554_, new_n56555_, new_n56556_, new_n56557_, new_n56558_,
    new_n56559_, new_n56560_, new_n56561_, new_n56562_, new_n56563_,
    new_n56564_, new_n56565_, new_n56566_, new_n56567_, new_n56568_,
    new_n56569_, new_n56570_, new_n56571_, new_n56572_, new_n56573_,
    new_n56574_, new_n56575_, new_n56576_, new_n56577_, new_n56578_,
    new_n56579_, new_n56580_, new_n56581_, new_n56582_, new_n56583_,
    new_n56584_, new_n56585_, new_n56586_, new_n56587_, new_n56588_,
    new_n56589_, new_n56590_, new_n56591_, new_n56592_, new_n56593_,
    new_n56594_, new_n56595_, new_n56596_, new_n56597_, new_n56598_,
    new_n56599_, new_n56600_, new_n56601_, new_n56602_, new_n56603_,
    new_n56604_, new_n56605_, new_n56606_, new_n56607_, new_n56608_,
    new_n56609_, new_n56610_, new_n56611_, new_n56612_, new_n56613_,
    new_n56614_, new_n56615_, new_n56616_, new_n56617_, new_n56618_,
    new_n56619_, new_n56620_, new_n56621_, new_n56622_, new_n56623_,
    new_n56624_, new_n56625_, new_n56626_, new_n56627_, new_n56628_,
    new_n56629_, new_n56630_, new_n56631_, new_n56632_, new_n56633_,
    new_n56634_, new_n56635_, new_n56636_, new_n56637_, new_n56638_,
    new_n56639_, new_n56640_, new_n56641_, new_n56642_, new_n56643_,
    new_n56644_, new_n56645_, new_n56646_, new_n56647_, new_n56648_,
    new_n56649_, new_n56650_, new_n56651_, new_n56652_, new_n56653_,
    new_n56654_, new_n56655_, new_n56656_, new_n56657_, new_n56658_,
    new_n56659_, new_n56660_, new_n56661_, new_n56662_, new_n56663_,
    new_n56664_, new_n56665_, new_n56666_, new_n56667_, new_n56668_,
    new_n56669_, new_n56670_, new_n56671_, new_n56672_, new_n56673_,
    new_n56674_, new_n56675_, new_n56676_, new_n56677_, new_n56678_,
    new_n56679_, new_n56680_, new_n56681_, new_n56682_, new_n56683_,
    new_n56684_, new_n56685_, new_n56686_, new_n56687_, new_n56688_,
    new_n56689_, new_n56690_, new_n56691_, new_n56692_, new_n56693_,
    new_n56694_, new_n56695_, new_n56696_, new_n56697_, new_n56698_,
    new_n56699_, new_n56700_, new_n56701_, new_n56702_, new_n56703_,
    new_n56704_, new_n56705_, new_n56706_, new_n56707_, new_n56708_,
    new_n56709_, new_n56710_, new_n56711_, new_n56712_, new_n56713_,
    new_n56714_, new_n56715_, new_n56716_, new_n56717_, new_n56718_,
    new_n56719_, new_n56720_, new_n56721_, new_n56722_, new_n56723_,
    new_n56724_, new_n56725_, new_n56726_, new_n56727_, new_n56728_,
    new_n56729_, new_n56730_, new_n56731_, new_n56732_, new_n56733_,
    new_n56734_, new_n56735_, new_n56736_, new_n56737_, new_n56738_,
    new_n56739_, new_n56740_, new_n56741_, new_n56742_, new_n56743_,
    new_n56744_, new_n56745_, new_n56746_, new_n56747_, new_n56748_,
    new_n56749_, new_n56750_, new_n56751_, new_n56752_, new_n56753_,
    new_n56754_, new_n56755_, new_n56756_, new_n56757_, new_n56758_,
    new_n56759_, new_n56760_, new_n56761_, new_n56762_, new_n56763_,
    new_n56764_, new_n56765_, new_n56766_, new_n56767_, new_n56768_,
    new_n56769_, new_n56770_, new_n56771_, new_n56772_, new_n56773_,
    new_n56774_, new_n56775_, new_n56776_, new_n56777_, new_n56778_,
    new_n56779_, new_n56780_, new_n56781_, new_n56782_, new_n56783_,
    new_n56784_, new_n56785_, new_n56786_, new_n56787_, new_n56788_,
    new_n56789_, new_n56790_, new_n56791_, new_n56792_, new_n56793_,
    new_n56794_, new_n56795_, new_n56796_, new_n56797_, new_n56798_,
    new_n56799_, new_n56800_, new_n56801_, new_n56802_, new_n56803_,
    new_n56804_, new_n56805_, new_n56806_, new_n56807_, new_n56808_,
    new_n56809_, new_n56810_, new_n56811_, new_n56812_, new_n56813_,
    new_n56814_, new_n56815_, new_n56816_, new_n56817_, new_n56818_,
    new_n56819_, new_n56820_, new_n56821_, new_n56822_, new_n56823_,
    new_n56824_, new_n56825_, new_n56826_, new_n56827_, new_n56828_,
    new_n56829_, new_n56830_, new_n56831_, new_n56832_, new_n56833_,
    new_n56834_, new_n56835_, new_n56836_, new_n56837_, new_n56838_,
    new_n56839_, new_n56840_, new_n56841_, new_n56842_, new_n56843_,
    new_n56844_, new_n56845_, new_n56846_, new_n56847_, new_n56848_,
    new_n56849_, new_n56850_, new_n56851_, new_n56852_, new_n56853_,
    new_n56854_, new_n56855_, new_n56856_, new_n56857_, new_n56858_,
    new_n56859_, new_n56860_, new_n56861_, new_n56862_, new_n56863_,
    new_n56864_, new_n56865_, new_n56866_, new_n56867_, new_n56868_,
    new_n56869_, new_n56870_, new_n56871_, new_n56872_, new_n56873_,
    new_n56874_, new_n56875_, new_n56876_, new_n56877_, new_n56878_,
    new_n56879_, new_n56880_, new_n56881_, new_n56882_, new_n56883_,
    new_n56884_, new_n56885_, new_n56886_, new_n56887_, new_n56888_,
    new_n56889_, new_n56890_, new_n56891_, new_n56892_, new_n56893_,
    new_n56894_, new_n56895_, new_n56896_, new_n56897_, new_n56898_,
    new_n56899_, new_n56900_, new_n56901_, new_n56902_, new_n56903_,
    new_n56904_, new_n56905_, new_n56906_, new_n56907_, new_n56908_,
    new_n56909_, new_n56910_, new_n56911_, new_n56912_, new_n56913_,
    new_n56914_, new_n56915_, new_n56916_, new_n56917_, new_n56918_,
    new_n56919_, new_n56920_, new_n56921_, new_n56922_, new_n56923_,
    new_n56924_, new_n56925_, new_n56926_, new_n56927_, new_n56928_,
    new_n56929_, new_n56930_, new_n56931_, new_n56932_, new_n56933_,
    new_n56934_, new_n56935_, new_n56936_, new_n56937_, new_n56938_,
    new_n56939_, new_n56940_, new_n56941_, new_n56942_, new_n56943_,
    new_n56944_, new_n56945_, new_n56946_, new_n56947_, new_n56948_,
    new_n56949_, new_n56950_, new_n56951_, new_n56952_, new_n56953_,
    new_n56954_, new_n56955_, new_n56956_, new_n56957_, new_n56958_,
    new_n56959_, new_n56960_, new_n56961_, new_n56962_, new_n56963_,
    new_n56964_, new_n56965_, new_n56966_, new_n56967_, new_n56968_,
    new_n56969_, new_n56970_, new_n56971_, new_n56972_, new_n56973_,
    new_n56974_, new_n56975_, new_n56976_, new_n56977_, new_n56978_,
    new_n56979_, new_n56980_, new_n56981_, new_n56982_, new_n56983_,
    new_n56984_, new_n56985_, new_n56986_, new_n56987_, new_n56988_,
    new_n56989_, new_n56990_, new_n56991_, new_n56992_, new_n56993_,
    new_n56994_, new_n56995_, new_n56996_, new_n56997_, new_n56998_,
    new_n56999_, new_n57001_, new_n57002_, new_n57003_, new_n57004_,
    new_n57005_, new_n57006_, new_n57008_, new_n57009_, new_n57010_,
    new_n57011_, new_n57012_, new_n57013_, new_n57014_, new_n57016_,
    new_n57017_, new_n57018_, new_n57019_, new_n57020_, new_n57021_,
    new_n57022_, new_n57024_, new_n57025_, new_n57026_, new_n57027_,
    new_n57028_, new_n57029_, new_n57030_, new_n57032_, new_n57033_,
    new_n57034_, new_n57035_, new_n57036_, new_n57037_, new_n57038_,
    new_n57040_, new_n57041_, new_n57042_, new_n57043_, new_n57044_,
    new_n57045_, new_n57046_, new_n57048_, new_n57049_, new_n57050_,
    new_n57051_, new_n57052_, new_n57053_, new_n57054_, new_n57056_,
    new_n57057_, new_n57058_, new_n57059_, new_n57060_, new_n57061_,
    new_n57062_, new_n57064_, new_n57065_, new_n57066_, new_n57067_,
    new_n57068_, new_n57069_, new_n57070_, new_n57072_, new_n57073_,
    new_n57074_, new_n57075_, new_n57076_, new_n57077_, new_n57078_,
    new_n57080_, new_n57081_, new_n57082_, new_n57083_, new_n57084_,
    new_n57085_, new_n57086_, new_n57088_, new_n57089_, new_n57090_,
    new_n57091_, new_n57092_, new_n57093_, new_n57094_, new_n57096_,
    new_n57097_, new_n57098_, new_n57099_, new_n57100_, new_n57101_,
    new_n57102_, new_n57104_, new_n57105_, new_n57106_, new_n57107_,
    new_n57108_, new_n57109_, new_n57110_, new_n57112_, new_n57113_,
    new_n57114_, new_n57115_, new_n57116_, new_n57117_, new_n57118_,
    new_n57120_, new_n57121_, new_n57122_, new_n57123_, new_n57124_,
    new_n57125_, new_n57126_, new_n57128_, new_n57129_, new_n57130_,
    new_n57131_, new_n57132_, new_n57133_, new_n57134_, new_n57136_,
    new_n57137_, new_n57138_, new_n57139_, new_n57140_, new_n57141_,
    new_n57142_, new_n57144_, new_n57145_, new_n57146_, new_n57147_,
    new_n57148_, new_n57149_, new_n57150_, new_n57152_, new_n57153_,
    new_n57154_, new_n57155_, new_n57156_, new_n57157_, new_n57158_,
    new_n57160_, new_n57161_, new_n57162_, new_n57163_, new_n57164_,
    new_n57165_, new_n57166_, new_n57168_, new_n57169_, new_n57170_,
    new_n57171_, new_n57172_, new_n57173_, new_n57174_, new_n57176_,
    new_n57177_, new_n57178_, new_n57179_, new_n57180_, new_n57181_,
    new_n57182_, new_n57184_, new_n57185_, new_n57186_, new_n57187_,
    new_n57188_, new_n57189_, new_n57190_, new_n57192_, new_n57193_,
    new_n57194_, new_n57195_, new_n57196_, new_n57197_, new_n57198_,
    new_n57200_, new_n57201_, new_n57202_, new_n57203_, new_n57204_,
    new_n57205_, new_n57206_, new_n57208_, new_n57209_, new_n57210_,
    new_n57211_, new_n57212_, new_n57213_, new_n57214_, new_n57216_,
    new_n57217_, new_n57218_, new_n57219_, new_n57220_, new_n57221_,
    new_n57222_, new_n57224_, new_n57225_, new_n57226_, new_n57227_,
    new_n57228_, new_n57229_, new_n57230_, new_n57232_, new_n57233_,
    new_n57234_, new_n57235_, new_n57236_, new_n57237_, new_n57238_,
    new_n57240_, new_n57241_, new_n57242_, new_n57243_, new_n57244_,
    new_n57245_, new_n57246_, new_n57248_, new_n57249_, new_n57250_,
    new_n57251_, new_n57252_, new_n57253_, new_n57254_, new_n57256_,
    new_n57257_, new_n57258_, new_n57259_, new_n57260_, new_n57261_,
    new_n57262_, new_n57264_, new_n57265_, new_n57266_, new_n57267_,
    new_n57268_, new_n57269_, new_n57270_, new_n57272_, new_n57273_,
    new_n57274_, new_n57275_, new_n57276_, new_n57277_, new_n57278_,
    new_n57280_, new_n57281_, new_n57282_, new_n57283_, new_n57284_,
    new_n57285_, new_n57286_, new_n57288_, new_n57289_, new_n57290_,
    new_n57291_, new_n57292_, new_n57293_, new_n57294_, new_n57296_,
    new_n57297_, new_n57298_, new_n57299_, new_n57300_, new_n57301_,
    new_n57302_, new_n57304_, new_n57305_, new_n57306_, new_n57307_,
    new_n57308_, new_n57309_, new_n57310_, new_n57312_, new_n57313_,
    new_n57314_, new_n57315_, new_n57316_, new_n57317_, new_n57318_,
    new_n57320_, new_n57321_, new_n57322_, new_n57323_, new_n57324_,
    new_n57325_, new_n57326_, new_n57328_, new_n57329_, new_n57330_,
    new_n57331_, new_n57332_, new_n57333_, new_n57334_, new_n57336_,
    new_n57337_, new_n57338_, new_n57339_, new_n57340_, new_n57341_,
    new_n57342_, new_n57344_, new_n57345_, new_n57346_, new_n57347_,
    new_n57348_, new_n57349_, new_n57350_, new_n57352_, new_n57353_,
    new_n57354_, new_n57355_, new_n57356_, new_n57357_, new_n57358_,
    new_n57360_, new_n57361_, new_n57362_, new_n57363_, new_n57364_,
    new_n57365_, new_n57366_, new_n57368_, new_n57369_, new_n57370_,
    new_n57371_, new_n57372_, new_n57373_, new_n57374_, new_n57376_,
    new_n57377_, new_n57378_, new_n57379_, new_n57380_, new_n57381_,
    new_n57382_, new_n57384_, new_n57385_, new_n57386_, new_n57387_,
    new_n57388_, new_n57389_, new_n57390_, new_n57392_, new_n57393_,
    new_n57394_, new_n57395_, new_n57396_, new_n57397_, new_n57398_,
    new_n57400_, new_n57401_, new_n57402_, new_n57403_, new_n57404_,
    new_n57405_, new_n57406_, new_n57408_, new_n57409_, new_n57410_,
    new_n57411_, new_n57412_, new_n57413_, new_n57414_, new_n57416_,
    new_n57417_, new_n57418_, new_n57419_, new_n57420_, new_n57421_,
    new_n57422_, new_n57424_, new_n57425_, new_n57426_, new_n57427_,
    new_n57428_, new_n57429_, new_n57430_, new_n57432_, new_n57433_,
    new_n57434_, new_n57435_, new_n57436_, new_n57437_, new_n57438_,
    new_n57440_, new_n57441_, new_n57442_, new_n57443_, new_n57444_,
    new_n57445_, new_n57446_, new_n57448_, new_n57449_, new_n57450_,
    new_n57451_, new_n57452_, new_n57453_, new_n57454_, new_n57456_,
    new_n57457_, new_n57458_, new_n57459_, new_n57460_, new_n57461_,
    new_n57462_, new_n57464_, new_n57465_, new_n57466_, new_n57467_,
    new_n57468_, new_n57469_, new_n57470_, new_n57472_, new_n57473_,
    new_n57474_, new_n57475_, new_n57476_, new_n57477_, new_n57478_,
    new_n57480_, new_n57481_, new_n57482_, new_n57483_, new_n57484_,
    new_n57485_, new_n57486_, new_n57488_, new_n57489_, new_n57490_,
    new_n57491_, new_n57492_, new_n57493_, new_n57494_, new_n57496_,
    new_n57497_, new_n57498_, new_n57499_, new_n57500_, new_n57501_,
    new_n57502_;
  assign new_n257_ = ~\a[63]  & \b[0] ;
  assign new_n258_ = \b[0]  & ~\b[1] ;
  assign new_n259_ = ~\b[2]  & ~\b[3] ;
  assign new_n260_ = new_n258_ & new_n259_;
  assign new_n261_ = ~new_n257_ & new_n260_;
  assign new_n262_ = ~\b[8]  & ~\b[9] ;
  assign new_n263_ = ~\b[10]  & ~\b[11] ;
  assign new_n264_ = new_n262_ & new_n263_;
  assign new_n265_ = ~\b[4]  & ~\b[5] ;
  assign new_n266_ = ~\b[6]  & ~\b[7] ;
  assign new_n267_ = new_n265_ & new_n266_;
  assign new_n268_ = new_n264_ & new_n267_;
  assign new_n269_ = ~\b[16]  & ~\b[17] ;
  assign new_n270_ = ~\b[18]  & ~\b[19] ;
  assign new_n271_ = new_n269_ & new_n270_;
  assign new_n272_ = ~\b[12]  & ~\b[13] ;
  assign new_n273_ = ~\b[14]  & ~\b[15] ;
  assign new_n274_ = new_n272_ & new_n273_;
  assign new_n275_ = new_n271_ & new_n274_;
  assign new_n276_ = new_n268_ & new_n275_;
  assign new_n277_ = new_n261_ & new_n276_;
  assign new_n278_ = ~\b[60]  & ~\b[61] ;
  assign new_n279_ = ~\b[62]  & ~\b[63] ;
  assign new_n280_ = new_n278_ & new_n279_;
  assign new_n281_ = ~\b[56]  & ~\b[57] ;
  assign new_n282_ = ~\b[58]  & ~\b[59] ;
  assign new_n283_ = new_n281_ & new_n282_;
  assign new_n284_ = ~\b[52]  & ~\b[53] ;
  assign new_n285_ = ~\b[54]  & ~\b[55] ;
  assign new_n286_ = new_n284_ & new_n285_;
  assign new_n287_ = new_n283_ & new_n286_;
  assign new_n288_ = new_n280_ & new_n287_;
  assign new_n289_ = ~\b[40]  & ~\b[41] ;
  assign new_n290_ = ~\b[42]  & ~\b[43] ;
  assign new_n291_ = new_n289_ & new_n290_;
  assign new_n292_ = ~\b[36]  & ~\b[37] ;
  assign new_n293_ = ~\b[38]  & ~\b[39] ;
  assign new_n294_ = new_n292_ & new_n293_;
  assign new_n295_ = new_n291_ & new_n294_;
  assign new_n296_ = ~\b[48]  & ~\b[49] ;
  assign new_n297_ = ~\b[50]  & ~\b[51] ;
  assign new_n298_ = new_n296_ & new_n297_;
  assign new_n299_ = ~\b[44]  & ~\b[45] ;
  assign new_n300_ = ~\b[46]  & ~\b[47] ;
  assign new_n301_ = new_n299_ & new_n300_;
  assign new_n302_ = new_n298_ & new_n301_;
  assign new_n303_ = new_n295_ & new_n302_;
  assign new_n304_ = ~\b[24]  & ~\b[25] ;
  assign new_n305_ = ~\b[26]  & ~\b[27] ;
  assign new_n306_ = new_n304_ & new_n305_;
  assign new_n307_ = ~\b[20]  & ~\b[21] ;
  assign new_n308_ = ~\b[22]  & ~\b[23] ;
  assign new_n309_ = new_n307_ & new_n308_;
  assign new_n310_ = new_n306_ & new_n309_;
  assign new_n311_ = ~\b[32]  & ~\b[33] ;
  assign new_n312_ = ~\b[34]  & ~\b[35] ;
  assign new_n313_ = new_n311_ & new_n312_;
  assign new_n314_ = ~\b[28]  & ~\b[29] ;
  assign new_n315_ = ~\b[30]  & ~\b[31] ;
  assign new_n316_ = new_n314_ & new_n315_;
  assign new_n317_ = new_n313_ & new_n316_;
  assign new_n318_ = new_n310_ & new_n317_;
  assign new_n319_ = new_n303_ & new_n318_;
  assign new_n320_ = new_n288_ & new_n319_;
  assign new_n321_ = new_n277_ & new_n320_;
  assign new_n322_ = ~\a[62]  & \b[0] ;
  assign new_n323_ = \b[1]  & new_n322_;
  assign new_n324_ = \a[63]  & ~new_n323_;
  assign new_n325_ = ~new_n321_ & new_n324_;
  assign new_n326_ = ~\b[1]  & ~new_n322_;
  assign new_n327_ = ~new_n325_ & ~new_n326_;
  assign new_n328_ = \a[63]  & ~new_n321_;
  assign new_n329_ = \b[1]  & ~new_n322_;
  assign new_n330_ = ~\b[1]  & new_n322_;
  assign new_n331_ = ~new_n329_ & ~new_n330_;
  assign new_n332_ = new_n259_ & new_n267_;
  assign new_n333_ = new_n264_ & new_n274_;
  assign new_n334_ = new_n332_ & new_n333_;
  assign new_n335_ = ~new_n331_ & new_n334_;
  assign new_n336_ = new_n286_ & new_n298_;
  assign new_n337_ = new_n280_ & new_n283_;
  assign new_n338_ = new_n336_ & new_n337_;
  assign new_n339_ = new_n294_ & new_n313_;
  assign new_n340_ = new_n291_ & new_n301_;
  assign new_n341_ = new_n339_ & new_n340_;
  assign new_n342_ = new_n271_ & new_n309_;
  assign new_n343_ = new_n306_ & new_n316_;
  assign new_n344_ = new_n342_ & new_n343_;
  assign new_n345_ = new_n341_ & new_n344_;
  assign new_n346_ = new_n338_ & new_n345_;
  assign new_n347_ = new_n335_ & new_n346_;
  assign new_n348_ = ~new_n328_ & new_n347_;
  assign new_n349_ = ~new_n327_ & new_n348_;
  assign new_n350_ = new_n333_ & new_n342_;
  assign new_n351_ = new_n332_ & new_n350_;
  assign new_n352_ = ~new_n323_ & ~new_n326_;
  assign new_n353_ = new_n337_ & new_n352_;
  assign new_n354_ = new_n336_ & new_n340_;
  assign new_n355_ = new_n339_ & new_n343_;
  assign new_n356_ = new_n354_ & new_n355_;
  assign new_n357_ = new_n353_ & new_n356_;
  assign new_n358_ = new_n351_ & new_n357_;
  assign new_n359_ = ~new_n327_ & new_n358_;
  assign new_n360_ = new_n328_ & ~new_n359_;
  assign new_n361_ = ~new_n349_ & ~new_n360_;
  assign new_n362_ = ~\a[61]  & \b[0] ;
  assign new_n363_ = \b[1]  & new_n362_;
  assign new_n364_ = ~\b[21]  & ~\b[22] ;
  assign new_n365_ = ~\b[23]  & ~\b[24] ;
  assign new_n366_ = new_n364_ & new_n365_;
  assign new_n367_ = ~\b[17]  & ~\b[18] ;
  assign new_n368_ = ~\b[19]  & ~\b[20] ;
  assign new_n369_ = new_n367_ & new_n368_;
  assign new_n370_ = new_n366_ & new_n369_;
  assign new_n371_ = ~\b[29]  & ~\b[30] ;
  assign new_n372_ = ~\b[31]  & ~\b[32] ;
  assign new_n373_ = new_n371_ & new_n372_;
  assign new_n374_ = ~\b[25]  & ~\b[26] ;
  assign new_n375_ = ~\b[27]  & ~\b[28] ;
  assign new_n376_ = new_n374_ & new_n375_;
  assign new_n377_ = new_n373_ & new_n376_;
  assign new_n378_ = new_n370_ & new_n377_;
  assign new_n379_ = ~\b[5]  & ~\b[6] ;
  assign new_n380_ = ~\b[7]  & ~\b[8] ;
  assign new_n381_ = new_n379_ & new_n380_;
  assign new_n382_ = \b[0]  & ~\b[2] ;
  assign new_n383_ = ~\b[3]  & ~\b[4] ;
  assign new_n384_ = new_n382_ & new_n383_;
  assign new_n385_ = new_n381_ & new_n384_;
  assign new_n386_ = ~\b[13]  & ~\b[14] ;
  assign new_n387_ = ~\b[15]  & ~\b[16] ;
  assign new_n388_ = new_n386_ & new_n387_;
  assign new_n389_ = ~\b[9]  & ~\b[10] ;
  assign new_n390_ = ~\b[11]  & ~\b[12] ;
  assign new_n391_ = new_n389_ & new_n390_;
  assign new_n392_ = new_n388_ & new_n391_;
  assign new_n393_ = new_n385_ & new_n392_;
  assign new_n394_ = new_n378_ & new_n393_;
  assign new_n395_ = ~\b[53]  & ~\b[54] ;
  assign new_n396_ = ~\b[55]  & ~\b[56] ;
  assign new_n397_ = new_n395_ & new_n396_;
  assign new_n398_ = ~\b[49]  & ~\b[50] ;
  assign new_n399_ = ~\b[51]  & ~\b[52] ;
  assign new_n400_ = new_n398_ & new_n399_;
  assign new_n401_ = new_n397_ & new_n400_;
  assign new_n402_ = ~\b[61]  & ~\b[62] ;
  assign new_n403_ = ~\b[63]  & new_n402_;
  assign new_n404_ = ~\b[57]  & ~\b[58] ;
  assign new_n405_ = ~\b[59]  & ~\b[60] ;
  assign new_n406_ = new_n404_ & new_n405_;
  assign new_n407_ = new_n403_ & new_n406_;
  assign new_n408_ = new_n401_ & new_n407_;
  assign new_n409_ = ~\b[37]  & ~\b[38] ;
  assign new_n410_ = ~\b[39]  & ~\b[40] ;
  assign new_n411_ = new_n409_ & new_n410_;
  assign new_n412_ = ~\b[33]  & ~\b[34] ;
  assign new_n413_ = ~\b[35]  & ~\b[36] ;
  assign new_n414_ = new_n412_ & new_n413_;
  assign new_n415_ = new_n411_ & new_n414_;
  assign new_n416_ = ~\b[45]  & ~\b[46] ;
  assign new_n417_ = ~\b[47]  & ~\b[48] ;
  assign new_n418_ = new_n416_ & new_n417_;
  assign new_n419_ = ~\b[41]  & ~\b[42] ;
  assign new_n420_ = ~\b[43]  & ~\b[44] ;
  assign new_n421_ = new_n419_ & new_n420_;
  assign new_n422_ = new_n418_ & new_n421_;
  assign new_n423_ = new_n415_ & new_n422_;
  assign new_n424_ = new_n408_ & new_n423_;
  assign new_n425_ = new_n394_ & new_n424_;
  assign new_n426_ = ~new_n327_ & new_n425_;
  assign new_n427_ = \a[62]  & ~new_n426_;
  assign new_n428_ = new_n259_ & new_n322_;
  assign new_n429_ = new_n267_ & new_n428_;
  assign new_n430_ = new_n333_ & new_n429_;
  assign new_n431_ = new_n344_ & new_n430_;
  assign new_n432_ = new_n338_ & new_n341_;
  assign new_n433_ = new_n431_ & new_n432_;
  assign new_n434_ = ~new_n327_ & new_n433_;
  assign new_n435_ = ~new_n427_ & ~new_n434_;
  assign new_n436_ = ~new_n363_ & ~new_n435_;
  assign new_n437_ = ~\b[1]  & ~new_n362_;
  assign new_n438_ = ~new_n436_ & ~new_n437_;
  assign new_n439_ = \b[2]  & ~new_n349_;
  assign new_n440_ = ~new_n360_ & new_n439_;
  assign new_n441_ = ~\b[2]  & ~new_n361_;
  assign new_n442_ = ~new_n440_ & ~new_n441_;
  assign new_n443_ = new_n438_ & ~new_n442_;
  assign new_n444_ = ~\b[2]  & ~new_n443_;
  assign new_n445_ = ~new_n438_ & ~new_n440_;
  assign new_n446_ = ~new_n441_ & ~new_n445_;
  assign new_n447_ = new_n381_ & new_n383_;
  assign new_n448_ = new_n392_ & new_n447_;
  assign new_n449_ = new_n378_ & new_n448_;
  assign new_n450_ = new_n424_ & new_n449_;
  assign \quotient[61]  = ~new_n446_ & new_n450_;
  assign new_n452_ = ~new_n444_ & \quotient[61] ;
  assign new_n453_ = ~new_n361_ & ~new_n452_;
  assign new_n454_ = ~new_n445_ & new_n450_;
  assign new_n455_ = ~new_n443_ & new_n454_;
  assign new_n456_ = ~new_n446_ & new_n455_;
  assign new_n457_ = \b[3]  & ~new_n456_;
  assign new_n458_ = ~new_n453_ & new_n457_;
  assign new_n459_ = new_n370_ & new_n392_;
  assign new_n460_ = new_n447_ & new_n459_;
  assign new_n461_ = ~new_n363_ & ~new_n437_;
  assign new_n462_ = new_n407_ & new_n461_;
  assign new_n463_ = new_n401_ & new_n422_;
  assign new_n464_ = new_n377_ & new_n415_;
  assign new_n465_ = new_n463_ & new_n464_;
  assign new_n466_ = new_n462_ & new_n465_;
  assign new_n467_ = new_n460_ & new_n466_;
  assign new_n468_ = ~new_n446_ & new_n467_;
  assign new_n469_ = ~new_n435_ & ~new_n468_;
  assign new_n470_ = \b[1]  & ~new_n362_;
  assign new_n471_ = ~\b[1]  & new_n362_;
  assign new_n472_ = ~new_n470_ & ~new_n471_;
  assign new_n473_ = new_n448_ & ~new_n472_;
  assign new_n474_ = new_n378_ & new_n423_;
  assign new_n475_ = new_n408_ & new_n474_;
  assign new_n476_ = new_n473_ & new_n475_;
  assign new_n477_ = ~new_n434_ & new_n476_;
  assign new_n478_ = ~new_n427_ & new_n477_;
  assign new_n479_ = ~new_n446_ & new_n478_;
  assign new_n480_ = ~new_n469_ & ~new_n479_;
  assign new_n481_ = ~\b[2]  & ~new_n480_;
  assign new_n482_ = \b[2]  & ~new_n479_;
  assign new_n483_ = ~new_n469_ & new_n482_;
  assign new_n484_ = \b[0]  & ~\b[3] ;
  assign new_n485_ = new_n267_ & new_n484_;
  assign new_n486_ = new_n333_ & new_n485_;
  assign new_n487_ = new_n344_ & new_n486_;
  assign new_n488_ = new_n432_ & new_n487_;
  assign new_n489_ = ~new_n446_ & new_n488_;
  assign new_n490_ = \a[61]  & ~new_n489_;
  assign new_n491_ = new_n362_ & new_n383_;
  assign new_n492_ = new_n381_ & new_n491_;
  assign new_n493_ = new_n392_ & new_n492_;
  assign new_n494_ = new_n378_ & new_n493_;
  assign new_n495_ = new_n424_ & new_n494_;
  assign new_n496_ = ~new_n446_ & new_n495_;
  assign new_n497_ = ~new_n490_ & ~new_n496_;
  assign new_n498_ = ~\a[60]  & \b[0] ;
  assign new_n499_ = \b[1]  & new_n498_;
  assign new_n500_ = ~new_n497_ & ~new_n499_;
  assign new_n501_ = ~\b[1]  & ~new_n498_;
  assign new_n502_ = ~new_n500_ & ~new_n501_;
  assign new_n503_ = ~new_n483_ & ~new_n502_;
  assign new_n504_ = ~new_n481_ & ~new_n503_;
  assign new_n505_ = ~new_n458_ & ~new_n504_;
  assign new_n506_ = ~new_n453_ & ~new_n456_;
  assign new_n507_ = ~\b[3]  & ~new_n506_;
  assign new_n508_ = ~new_n505_ & ~new_n507_;
  assign new_n509_ = ~new_n458_ & ~new_n507_;
  assign new_n510_ = ~new_n504_ & new_n509_;
  assign new_n511_ = new_n276_ & new_n318_;
  assign new_n512_ = new_n288_ & new_n303_;
  assign new_n513_ = new_n511_ & new_n512_;
  assign new_n514_ = new_n504_ & ~new_n509_;
  assign new_n515_ = new_n513_ & ~new_n514_;
  assign new_n516_ = ~new_n510_ & new_n515_;
  assign new_n517_ = ~new_n508_ & new_n516_;
  assign \quotient[60]  = ~new_n508_ & new_n513_;
  assign new_n519_ = ~new_n506_ & ~\quotient[60] ;
  assign new_n520_ = \b[4]  & ~new_n519_;
  assign new_n521_ = ~new_n517_ & new_n520_;
  assign new_n522_ = ~new_n481_ & ~new_n483_;
  assign new_n523_ = new_n502_ & ~new_n522_;
  assign new_n524_ = ~new_n503_ & new_n513_;
  assign new_n525_ = ~new_n523_ & new_n524_;
  assign new_n526_ = ~new_n508_ & new_n525_;
  assign new_n527_ = ~\b[2]  & ~new_n523_;
  assign new_n528_ = new_n513_ & ~new_n527_;
  assign new_n529_ = ~new_n508_ & new_n528_;
  assign new_n530_ = ~new_n480_ & ~new_n529_;
  assign new_n531_ = ~new_n526_ & ~new_n530_;
  assign new_n532_ = ~\b[3]  & ~new_n531_;
  assign new_n533_ = \b[3]  & ~new_n526_;
  assign new_n534_ = ~new_n530_ & new_n533_;
  assign new_n535_ = new_n275_ & new_n310_;
  assign new_n536_ = new_n268_ & new_n535_;
  assign new_n537_ = new_n280_ & ~new_n499_;
  assign new_n538_ = ~new_n501_ & new_n537_;
  assign new_n539_ = new_n287_ & new_n302_;
  assign new_n540_ = new_n295_ & new_n317_;
  assign new_n541_ = new_n539_ & new_n540_;
  assign new_n542_ = new_n538_ & new_n541_;
  assign new_n543_ = new_n536_ & new_n542_;
  assign new_n544_ = ~new_n508_ & new_n543_;
  assign new_n545_ = ~new_n497_ & ~new_n544_;
  assign new_n546_ = \b[1]  & ~new_n498_;
  assign new_n547_ = ~\b[1]  & new_n498_;
  assign new_n548_ = ~new_n546_ & ~new_n547_;
  assign new_n549_ = new_n276_ & ~new_n548_;
  assign new_n550_ = new_n320_ & new_n549_;
  assign new_n551_ = ~new_n496_ & new_n550_;
  assign new_n552_ = ~new_n490_ & new_n551_;
  assign new_n553_ = ~new_n508_ & new_n552_;
  assign new_n554_ = ~new_n545_ & ~new_n553_;
  assign new_n555_ = ~\b[2]  & ~new_n554_;
  assign new_n556_ = \b[2]  & ~new_n553_;
  assign new_n557_ = ~new_n545_ & new_n556_;
  assign new_n558_ = ~\a[59]  & \b[0] ;
  assign new_n559_ = \b[1]  & new_n558_;
  assign new_n560_ = \b[0]  & ~\b[4] ;
  assign new_n561_ = new_n381_ & new_n560_;
  assign new_n562_ = new_n392_ & new_n561_;
  assign new_n563_ = new_n378_ & new_n562_;
  assign new_n564_ = new_n424_ & new_n563_;
  assign new_n565_ = ~new_n508_ & new_n564_;
  assign new_n566_ = \a[60]  & ~new_n565_;
  assign new_n567_ = new_n267_ & new_n498_;
  assign new_n568_ = new_n333_ & new_n567_;
  assign new_n569_ = new_n344_ & new_n568_;
  assign new_n570_ = new_n432_ & new_n569_;
  assign new_n571_ = ~new_n508_ & new_n570_;
  assign new_n572_ = ~new_n566_ & ~new_n571_;
  assign new_n573_ = ~new_n559_ & ~new_n572_;
  assign new_n574_ = ~\b[1]  & ~new_n558_;
  assign new_n575_ = ~new_n573_ & ~new_n574_;
  assign new_n576_ = ~new_n557_ & ~new_n575_;
  assign new_n577_ = ~new_n555_ & ~new_n576_;
  assign new_n578_ = ~new_n534_ & ~new_n577_;
  assign new_n579_ = ~new_n532_ & ~new_n578_;
  assign new_n580_ = ~new_n521_ & ~new_n579_;
  assign new_n581_ = ~new_n517_ & ~new_n519_;
  assign new_n582_ = ~\b[4]  & ~new_n581_;
  assign new_n583_ = ~new_n580_ & ~new_n582_;
  assign new_n584_ = ~new_n532_ & ~new_n534_;
  assign new_n585_ = ~new_n555_ & ~new_n584_;
  assign new_n586_ = ~new_n576_ & new_n585_;
  assign new_n587_ = new_n366_ & new_n376_;
  assign new_n588_ = new_n373_ & new_n414_;
  assign new_n589_ = new_n587_ & new_n588_;
  assign new_n590_ = new_n381_ & new_n391_;
  assign new_n591_ = new_n369_ & new_n388_;
  assign new_n592_ = new_n590_ & new_n591_;
  assign new_n593_ = new_n589_ & new_n592_;
  assign new_n594_ = new_n397_ & new_n406_;
  assign new_n595_ = new_n403_ & new_n594_;
  assign new_n596_ = new_n411_ & new_n421_;
  assign new_n597_ = new_n400_ & new_n418_;
  assign new_n598_ = new_n596_ & new_n597_;
  assign new_n599_ = new_n595_ & new_n598_;
  assign new_n600_ = new_n593_ & new_n599_;
  assign new_n601_ = ~new_n586_ & new_n600_;
  assign new_n602_ = ~new_n578_ & new_n601_;
  assign new_n603_ = ~new_n583_ & new_n602_;
  assign new_n604_ = ~\b[3]  & ~new_n586_;
  assign new_n605_ = new_n600_ & ~new_n604_;
  assign new_n606_ = ~new_n583_ & new_n605_;
  assign new_n607_ = ~new_n531_ & ~new_n606_;
  assign new_n608_ = ~new_n603_ & ~new_n607_;
  assign new_n609_ = \b[4]  & ~new_n608_;
  assign new_n610_ = ~\b[4]  & ~new_n603_;
  assign new_n611_ = ~new_n607_ & new_n610_;
  assign new_n612_ = ~new_n609_ & ~new_n611_;
  assign new_n613_ = ~new_n555_ & ~new_n557_;
  assign new_n614_ = new_n575_ & ~new_n613_;
  assign new_n615_ = ~new_n576_ & new_n600_;
  assign new_n616_ = ~new_n614_ & new_n615_;
  assign new_n617_ = ~new_n583_ & new_n616_;
  assign new_n618_ = ~\b[2]  & ~new_n614_;
  assign new_n619_ = new_n600_ & ~new_n618_;
  assign new_n620_ = ~new_n583_ & new_n619_;
  assign new_n621_ = ~new_n554_ & ~new_n620_;
  assign new_n622_ = ~new_n617_ & ~new_n621_;
  assign new_n623_ = \b[3]  & ~new_n622_;
  assign new_n624_ = ~\b[3]  & ~new_n617_;
  assign new_n625_ = ~new_n621_ & new_n624_;
  assign new_n626_ = ~new_n623_ & ~new_n625_;
  assign new_n627_ = new_n587_ & new_n591_;
  assign new_n628_ = new_n590_ & new_n627_;
  assign new_n629_ = new_n403_ & ~new_n559_;
  assign new_n630_ = ~new_n574_ & new_n629_;
  assign new_n631_ = new_n594_ & new_n597_;
  assign new_n632_ = new_n588_ & new_n596_;
  assign new_n633_ = new_n631_ & new_n632_;
  assign new_n634_ = new_n630_ & new_n633_;
  assign new_n635_ = new_n628_ & new_n634_;
  assign new_n636_ = ~new_n583_ & new_n635_;
  assign new_n637_ = ~new_n572_ & ~new_n636_;
  assign new_n638_ = \b[1]  & ~new_n558_;
  assign new_n639_ = ~\b[1]  & new_n558_;
  assign new_n640_ = ~new_n638_ & ~new_n639_;
  assign new_n641_ = new_n592_ & ~new_n640_;
  assign new_n642_ = new_n589_ & new_n598_;
  assign new_n643_ = new_n595_ & new_n642_;
  assign new_n644_ = new_n641_ & new_n643_;
  assign new_n645_ = ~new_n571_ & new_n644_;
  assign new_n646_ = ~new_n566_ & new_n645_;
  assign new_n647_ = ~new_n583_ & new_n646_;
  assign new_n648_ = ~new_n637_ & ~new_n647_;
  assign new_n649_ = ~\b[2]  & ~new_n648_;
  assign new_n650_ = \b[0]  & ~\b[5] ;
  assign new_n651_ = new_n266_ & new_n650_;
  assign new_n652_ = new_n264_ & new_n651_;
  assign new_n653_ = new_n275_ & new_n652_;
  assign new_n654_ = new_n318_ & new_n653_;
  assign new_n655_ = new_n512_ & new_n654_;
  assign new_n656_ = ~new_n583_ & new_n655_;
  assign new_n657_ = \a[59]  & ~new_n656_;
  assign new_n658_ = new_n381_ & new_n558_;
  assign new_n659_ = new_n392_ & new_n658_;
  assign new_n660_ = new_n378_ & new_n659_;
  assign new_n661_ = new_n424_ & new_n660_;
  assign new_n662_ = ~new_n583_ & new_n661_;
  assign new_n663_ = ~new_n657_ & ~new_n662_;
  assign new_n664_ = \b[1]  & ~new_n663_;
  assign new_n665_ = ~\b[1]  & ~new_n662_;
  assign new_n666_ = ~new_n657_ & new_n665_;
  assign new_n667_ = ~new_n664_ & ~new_n666_;
  assign new_n668_ = ~\a[58]  & \b[0] ;
  assign new_n669_ = ~new_n667_ & ~new_n668_;
  assign new_n670_ = ~\b[1]  & ~new_n663_;
  assign new_n671_ = ~new_n669_ & ~new_n670_;
  assign new_n672_ = \b[2]  & ~new_n647_;
  assign new_n673_ = ~new_n637_ & new_n672_;
  assign new_n674_ = ~new_n649_ & ~new_n673_;
  assign new_n675_ = ~new_n671_ & new_n674_;
  assign new_n676_ = ~new_n649_ & ~new_n675_;
  assign new_n677_ = ~new_n626_ & ~new_n676_;
  assign new_n678_ = ~\b[3]  & ~new_n622_;
  assign new_n679_ = ~new_n677_ & ~new_n678_;
  assign new_n680_ = ~new_n612_ & ~new_n679_;
  assign new_n681_ = ~\b[4]  & ~new_n608_;
  assign new_n682_ = ~new_n680_ & ~new_n681_;
  assign new_n683_ = ~new_n521_ & ~new_n582_;
  assign new_n684_ = ~new_n532_ & ~new_n683_;
  assign new_n685_ = ~new_n578_ & new_n684_;
  assign new_n686_ = new_n600_ & ~new_n685_;
  assign new_n687_ = ~new_n580_ & new_n686_;
  assign new_n688_ = ~new_n583_ & new_n687_;
  assign new_n689_ = ~\b[4]  & ~new_n685_;
  assign new_n690_ = new_n600_ & ~new_n689_;
  assign new_n691_ = ~new_n583_ & new_n690_;
  assign new_n692_ = ~new_n581_ & ~new_n691_;
  assign new_n693_ = ~new_n688_ & ~new_n692_;
  assign new_n694_ = \b[5]  & ~new_n693_;
  assign new_n695_ = ~\b[5]  & ~new_n688_;
  assign new_n696_ = ~new_n692_ & new_n695_;
  assign new_n697_ = ~new_n694_ & ~new_n696_;
  assign new_n698_ = new_n264_ & new_n266_;
  assign new_n699_ = new_n275_ & new_n698_;
  assign new_n700_ = new_n318_ & new_n699_;
  assign new_n701_ = new_n512_ & new_n700_;
  assign new_n702_ = ~new_n697_ & new_n701_;
  assign new_n703_ = ~new_n682_ & new_n702_;
  assign new_n704_ = new_n600_ & ~new_n693_;
  assign \quotient[58]  = new_n703_ | new_n704_;
  assign new_n706_ = new_n612_ & ~new_n678_;
  assign new_n707_ = ~new_n677_ & new_n706_;
  assign new_n708_ = ~new_n680_ & ~new_n707_;
  assign new_n709_ = \quotient[58]  & new_n708_;
  assign new_n710_ = ~new_n608_ & ~new_n704_;
  assign new_n711_ = ~new_n703_ & new_n710_;
  assign new_n712_ = ~new_n709_ & ~new_n711_;
  assign new_n713_ = ~new_n682_ & ~new_n697_;
  assign new_n714_ = ~new_n681_ & new_n697_;
  assign new_n715_ = ~new_n680_ & new_n714_;
  assign new_n716_ = ~new_n713_ & ~new_n715_;
  assign new_n717_ = \quotient[58]  & new_n716_;
  assign new_n718_ = ~new_n693_ & ~new_n704_;
  assign new_n719_ = ~new_n703_ & new_n718_;
  assign new_n720_ = ~new_n717_ & ~new_n719_;
  assign new_n721_ = ~\b[6]  & ~new_n720_;
  assign new_n722_ = ~\b[5]  & ~new_n712_;
  assign new_n723_ = new_n626_ & ~new_n649_;
  assign new_n724_ = ~new_n675_ & new_n723_;
  assign new_n725_ = ~new_n677_ & ~new_n724_;
  assign new_n726_ = \quotient[58]  & new_n725_;
  assign new_n727_ = ~new_n622_ & ~new_n704_;
  assign new_n728_ = ~new_n703_ & new_n727_;
  assign new_n729_ = ~new_n726_ & ~new_n728_;
  assign new_n730_ = ~\b[4]  & ~new_n729_;
  assign new_n731_ = ~new_n670_ & new_n674_;
  assign new_n732_ = ~new_n669_ & new_n731_;
  assign new_n733_ = ~new_n671_ & ~new_n674_;
  assign new_n734_ = ~new_n732_ & ~new_n733_;
  assign new_n735_ = \quotient[58]  & ~new_n734_;
  assign new_n736_ = ~new_n648_ & ~new_n704_;
  assign new_n737_ = ~new_n703_ & new_n736_;
  assign new_n738_ = ~new_n735_ & ~new_n737_;
  assign new_n739_ = ~\b[3]  & ~new_n738_;
  assign new_n740_ = ~new_n666_ & new_n668_;
  assign new_n741_ = ~new_n664_ & new_n740_;
  assign new_n742_ = ~new_n669_ & ~new_n741_;
  assign new_n743_ = \quotient[58]  & new_n742_;
  assign new_n744_ = ~new_n663_ & ~new_n704_;
  assign new_n745_ = ~new_n703_ & new_n744_;
  assign new_n746_ = ~new_n743_ & ~new_n745_;
  assign new_n747_ = ~\b[2]  & ~new_n746_;
  assign new_n748_ = \b[0]  & \quotient[58] ;
  assign new_n749_ = \a[58]  & ~new_n748_;
  assign new_n750_ = new_n668_ & \quotient[58] ;
  assign new_n751_ = ~new_n749_ & ~new_n750_;
  assign new_n752_ = \b[1]  & ~new_n751_;
  assign new_n753_ = ~\b[1]  & ~new_n750_;
  assign new_n754_ = ~new_n749_ & new_n753_;
  assign new_n755_ = ~new_n752_ & ~new_n754_;
  assign new_n756_ = ~\a[57]  & \b[0] ;
  assign new_n757_ = ~new_n755_ & ~new_n756_;
  assign new_n758_ = ~\b[1]  & ~new_n751_;
  assign new_n759_ = ~new_n757_ & ~new_n758_;
  assign new_n760_ = \b[2]  & ~new_n745_;
  assign new_n761_ = ~new_n743_ & new_n760_;
  assign new_n762_ = ~new_n747_ & ~new_n761_;
  assign new_n763_ = ~new_n759_ & new_n762_;
  assign new_n764_ = ~new_n747_ & ~new_n763_;
  assign new_n765_ = \b[3]  & ~new_n737_;
  assign new_n766_ = ~new_n735_ & new_n765_;
  assign new_n767_ = ~new_n739_ & ~new_n766_;
  assign new_n768_ = ~new_n764_ & new_n767_;
  assign new_n769_ = ~new_n739_ & ~new_n768_;
  assign new_n770_ = \b[4]  & ~new_n728_;
  assign new_n771_ = ~new_n726_ & new_n770_;
  assign new_n772_ = ~new_n730_ & ~new_n771_;
  assign new_n773_ = ~new_n769_ & new_n772_;
  assign new_n774_ = ~new_n730_ & ~new_n773_;
  assign new_n775_ = \b[5]  & ~new_n711_;
  assign new_n776_ = ~new_n709_ & new_n775_;
  assign new_n777_ = ~new_n722_ & ~new_n776_;
  assign new_n778_ = ~new_n774_ & new_n777_;
  assign new_n779_ = ~new_n722_ & ~new_n778_;
  assign new_n780_ = \b[6]  & ~new_n719_;
  assign new_n781_ = ~new_n717_ & new_n780_;
  assign new_n782_ = ~new_n721_ & ~new_n781_;
  assign new_n783_ = ~new_n779_ & new_n782_;
  assign new_n784_ = ~new_n721_ & ~new_n783_;
  assign new_n785_ = new_n380_ & new_n391_;
  assign new_n786_ = new_n591_ & new_n785_;
  assign new_n787_ = new_n589_ & new_n786_;
  assign new_n788_ = new_n599_ & new_n787_;
  assign \quotient[57]  = ~new_n784_ & new_n788_;
  assign new_n790_ = ~new_n712_ & ~\quotient[57] ;
  assign new_n791_ = ~new_n730_ & new_n777_;
  assign new_n792_ = ~new_n773_ & new_n791_;
  assign new_n793_ = ~new_n774_ & ~new_n777_;
  assign new_n794_ = ~new_n792_ & ~new_n793_;
  assign new_n795_ = new_n788_ & ~new_n794_;
  assign new_n796_ = ~new_n784_ & new_n795_;
  assign new_n797_ = ~new_n790_ & ~new_n796_;
  assign new_n798_ = ~new_n720_ & ~\quotient[57] ;
  assign new_n799_ = ~new_n722_ & new_n782_;
  assign new_n800_ = ~new_n778_ & new_n799_;
  assign new_n801_ = ~new_n779_ & ~new_n782_;
  assign new_n802_ = ~new_n800_ & ~new_n801_;
  assign new_n803_ = \quotient[57]  & ~new_n802_;
  assign new_n804_ = ~new_n798_ & ~new_n803_;
  assign new_n805_ = ~\b[7]  & ~new_n804_;
  assign new_n806_ = ~\b[6]  & ~new_n797_;
  assign new_n807_ = ~new_n729_ & ~\quotient[57] ;
  assign new_n808_ = ~new_n739_ & new_n772_;
  assign new_n809_ = ~new_n768_ & new_n808_;
  assign new_n810_ = ~new_n769_ & ~new_n772_;
  assign new_n811_ = ~new_n809_ & ~new_n810_;
  assign new_n812_ = new_n788_ & ~new_n811_;
  assign new_n813_ = ~new_n784_ & new_n812_;
  assign new_n814_ = ~new_n807_ & ~new_n813_;
  assign new_n815_ = ~\b[5]  & ~new_n814_;
  assign new_n816_ = ~new_n738_ & ~\quotient[57] ;
  assign new_n817_ = ~new_n747_ & new_n767_;
  assign new_n818_ = ~new_n763_ & new_n817_;
  assign new_n819_ = ~new_n764_ & ~new_n767_;
  assign new_n820_ = ~new_n818_ & ~new_n819_;
  assign new_n821_ = new_n788_ & ~new_n820_;
  assign new_n822_ = ~new_n784_ & new_n821_;
  assign new_n823_ = ~new_n816_ & ~new_n822_;
  assign new_n824_ = ~\b[4]  & ~new_n823_;
  assign new_n825_ = ~new_n746_ & ~\quotient[57] ;
  assign new_n826_ = ~new_n758_ & new_n762_;
  assign new_n827_ = ~new_n757_ & new_n826_;
  assign new_n828_ = ~new_n759_ & ~new_n762_;
  assign new_n829_ = ~new_n827_ & ~new_n828_;
  assign new_n830_ = new_n788_ & ~new_n829_;
  assign new_n831_ = ~new_n784_ & new_n830_;
  assign new_n832_ = ~new_n825_ & ~new_n831_;
  assign new_n833_ = ~\b[3]  & ~new_n832_;
  assign new_n834_ = ~new_n751_ & ~\quotient[57] ;
  assign new_n835_ = ~new_n754_ & new_n756_;
  assign new_n836_ = ~new_n752_ & new_n835_;
  assign new_n837_ = new_n788_ & ~new_n836_;
  assign new_n838_ = ~new_n757_ & new_n837_;
  assign new_n839_ = ~new_n784_ & new_n838_;
  assign new_n840_ = ~new_n834_ & ~new_n839_;
  assign new_n841_ = ~\b[2]  & ~new_n840_;
  assign new_n842_ = \b[0]  & ~\b[7] ;
  assign new_n843_ = new_n264_ & new_n842_;
  assign new_n844_ = new_n275_ & new_n843_;
  assign new_n845_ = new_n318_ & new_n844_;
  assign new_n846_ = new_n512_ & new_n845_;
  assign new_n847_ = ~new_n784_ & new_n846_;
  assign new_n848_ = \a[57]  & ~new_n847_;
  assign new_n849_ = new_n380_ & new_n756_;
  assign new_n850_ = new_n391_ & new_n849_;
  assign new_n851_ = new_n591_ & new_n850_;
  assign new_n852_ = new_n589_ & new_n851_;
  assign new_n853_ = new_n599_ & new_n852_;
  assign new_n854_ = ~new_n784_ & new_n853_;
  assign new_n855_ = ~new_n848_ & ~new_n854_;
  assign new_n856_ = \b[1]  & ~new_n855_;
  assign new_n857_ = ~\b[1]  & ~new_n854_;
  assign new_n858_ = ~new_n848_ & new_n857_;
  assign new_n859_ = ~new_n856_ & ~new_n858_;
  assign new_n860_ = ~\a[56]  & \b[0] ;
  assign new_n861_ = ~new_n859_ & ~new_n860_;
  assign new_n862_ = ~\b[1]  & ~new_n855_;
  assign new_n863_ = ~new_n861_ & ~new_n862_;
  assign new_n864_ = \b[2]  & ~new_n839_;
  assign new_n865_ = ~new_n834_ & new_n864_;
  assign new_n866_ = ~new_n841_ & ~new_n865_;
  assign new_n867_ = ~new_n863_ & new_n866_;
  assign new_n868_ = ~new_n841_ & ~new_n867_;
  assign new_n869_ = \b[3]  & ~new_n831_;
  assign new_n870_ = ~new_n825_ & new_n869_;
  assign new_n871_ = ~new_n833_ & ~new_n870_;
  assign new_n872_ = ~new_n868_ & new_n871_;
  assign new_n873_ = ~new_n833_ & ~new_n872_;
  assign new_n874_ = \b[4]  & ~new_n822_;
  assign new_n875_ = ~new_n816_ & new_n874_;
  assign new_n876_ = ~new_n824_ & ~new_n875_;
  assign new_n877_ = ~new_n873_ & new_n876_;
  assign new_n878_ = ~new_n824_ & ~new_n877_;
  assign new_n879_ = \b[5]  & ~new_n813_;
  assign new_n880_ = ~new_n807_ & new_n879_;
  assign new_n881_ = ~new_n815_ & ~new_n880_;
  assign new_n882_ = ~new_n878_ & new_n881_;
  assign new_n883_ = ~new_n815_ & ~new_n882_;
  assign new_n884_ = \b[6]  & ~new_n796_;
  assign new_n885_ = ~new_n790_ & new_n884_;
  assign new_n886_ = ~new_n806_ & ~new_n885_;
  assign new_n887_ = ~new_n883_ & new_n886_;
  assign new_n888_ = ~new_n806_ & ~new_n887_;
  assign new_n889_ = \b[7]  & ~new_n798_;
  assign new_n890_ = ~new_n803_ & new_n889_;
  assign new_n891_ = ~new_n805_ & ~new_n890_;
  assign new_n892_ = ~new_n888_ & new_n891_;
  assign new_n893_ = ~new_n805_ & ~new_n892_;
  assign new_n894_ = new_n333_ & new_n344_;
  assign new_n895_ = new_n432_ & new_n894_;
  assign \quotient[56]  = ~new_n893_ & new_n895_;
  assign new_n897_ = ~new_n797_ & ~\quotient[56] ;
  assign new_n898_ = ~new_n815_ & new_n886_;
  assign new_n899_ = ~new_n882_ & new_n898_;
  assign new_n900_ = ~new_n883_ & ~new_n886_;
  assign new_n901_ = ~new_n899_ & ~new_n900_;
  assign new_n902_ = new_n895_ & ~new_n901_;
  assign new_n903_ = ~new_n893_ & new_n902_;
  assign new_n904_ = ~new_n897_ & ~new_n903_;
  assign new_n905_ = ~\b[7]  & ~new_n904_;
  assign new_n906_ = ~new_n814_ & ~\quotient[56] ;
  assign new_n907_ = ~new_n824_ & new_n881_;
  assign new_n908_ = ~new_n877_ & new_n907_;
  assign new_n909_ = ~new_n878_ & ~new_n881_;
  assign new_n910_ = ~new_n908_ & ~new_n909_;
  assign new_n911_ = new_n895_ & ~new_n910_;
  assign new_n912_ = ~new_n893_ & new_n911_;
  assign new_n913_ = ~new_n906_ & ~new_n912_;
  assign new_n914_ = ~\b[6]  & ~new_n913_;
  assign new_n915_ = ~new_n823_ & ~\quotient[56] ;
  assign new_n916_ = ~new_n833_ & new_n876_;
  assign new_n917_ = ~new_n872_ & new_n916_;
  assign new_n918_ = ~new_n873_ & ~new_n876_;
  assign new_n919_ = ~new_n917_ & ~new_n918_;
  assign new_n920_ = new_n895_ & ~new_n919_;
  assign new_n921_ = ~new_n893_ & new_n920_;
  assign new_n922_ = ~new_n915_ & ~new_n921_;
  assign new_n923_ = ~\b[5]  & ~new_n922_;
  assign new_n924_ = ~new_n832_ & ~\quotient[56] ;
  assign new_n925_ = ~new_n841_ & new_n871_;
  assign new_n926_ = ~new_n867_ & new_n925_;
  assign new_n927_ = ~new_n868_ & ~new_n871_;
  assign new_n928_ = ~new_n926_ & ~new_n927_;
  assign new_n929_ = new_n895_ & ~new_n928_;
  assign new_n930_ = ~new_n893_ & new_n929_;
  assign new_n931_ = ~new_n924_ & ~new_n930_;
  assign new_n932_ = ~\b[4]  & ~new_n931_;
  assign new_n933_ = ~new_n840_ & ~\quotient[56] ;
  assign new_n934_ = ~new_n862_ & new_n866_;
  assign new_n935_ = ~new_n861_ & new_n934_;
  assign new_n936_ = ~new_n863_ & ~new_n866_;
  assign new_n937_ = ~new_n935_ & ~new_n936_;
  assign new_n938_ = new_n895_ & ~new_n937_;
  assign new_n939_ = ~new_n893_ & new_n938_;
  assign new_n940_ = ~new_n933_ & ~new_n939_;
  assign new_n941_ = ~\b[3]  & ~new_n940_;
  assign new_n942_ = ~new_n855_ & ~\quotient[56] ;
  assign new_n943_ = ~new_n858_ & new_n860_;
  assign new_n944_ = ~new_n856_ & new_n943_;
  assign new_n945_ = new_n895_ & ~new_n944_;
  assign new_n946_ = ~new_n861_ & new_n945_;
  assign new_n947_ = ~new_n893_ & new_n946_;
  assign new_n948_ = ~new_n942_ & ~new_n947_;
  assign new_n949_ = ~\b[2]  & ~new_n948_;
  assign new_n950_ = \b[0]  & ~\b[8] ;
  assign new_n951_ = new_n391_ & new_n950_;
  assign new_n952_ = new_n591_ & new_n951_;
  assign new_n953_ = new_n589_ & new_n952_;
  assign new_n954_ = new_n599_ & new_n953_;
  assign new_n955_ = ~new_n893_ & new_n954_;
  assign new_n956_ = \a[56]  & ~new_n955_;
  assign new_n957_ = new_n264_ & new_n860_;
  assign new_n958_ = new_n275_ & new_n957_;
  assign new_n959_ = new_n318_ & new_n958_;
  assign new_n960_ = new_n512_ & new_n959_;
  assign new_n961_ = ~new_n893_ & new_n960_;
  assign new_n962_ = ~new_n956_ & ~new_n961_;
  assign new_n963_ = \b[1]  & ~new_n962_;
  assign new_n964_ = ~\b[1]  & ~new_n961_;
  assign new_n965_ = ~new_n956_ & new_n964_;
  assign new_n966_ = ~new_n963_ & ~new_n965_;
  assign new_n967_ = ~\a[55]  & \b[0] ;
  assign new_n968_ = ~new_n966_ & ~new_n967_;
  assign new_n969_ = ~\b[1]  & ~new_n962_;
  assign new_n970_ = ~new_n968_ & ~new_n969_;
  assign new_n971_ = \b[2]  & ~new_n947_;
  assign new_n972_ = ~new_n942_ & new_n971_;
  assign new_n973_ = ~new_n949_ & ~new_n972_;
  assign new_n974_ = ~new_n970_ & new_n973_;
  assign new_n975_ = ~new_n949_ & ~new_n974_;
  assign new_n976_ = \b[3]  & ~new_n939_;
  assign new_n977_ = ~new_n933_ & new_n976_;
  assign new_n978_ = ~new_n941_ & ~new_n977_;
  assign new_n979_ = ~new_n975_ & new_n978_;
  assign new_n980_ = ~new_n941_ & ~new_n979_;
  assign new_n981_ = \b[4]  & ~new_n930_;
  assign new_n982_ = ~new_n924_ & new_n981_;
  assign new_n983_ = ~new_n932_ & ~new_n982_;
  assign new_n984_ = ~new_n980_ & new_n983_;
  assign new_n985_ = ~new_n932_ & ~new_n984_;
  assign new_n986_ = \b[5]  & ~new_n921_;
  assign new_n987_ = ~new_n915_ & new_n986_;
  assign new_n988_ = ~new_n923_ & ~new_n987_;
  assign new_n989_ = ~new_n985_ & new_n988_;
  assign new_n990_ = ~new_n923_ & ~new_n989_;
  assign new_n991_ = \b[6]  & ~new_n912_;
  assign new_n992_ = ~new_n906_ & new_n991_;
  assign new_n993_ = ~new_n914_ & ~new_n992_;
  assign new_n994_ = ~new_n990_ & new_n993_;
  assign new_n995_ = ~new_n914_ & ~new_n994_;
  assign new_n996_ = \b[7]  & ~new_n903_;
  assign new_n997_ = ~new_n897_ & new_n996_;
  assign new_n998_ = ~new_n905_ & ~new_n997_;
  assign new_n999_ = ~new_n995_ & new_n998_;
  assign new_n1000_ = ~new_n905_ & ~new_n999_;
  assign new_n1001_ = ~new_n804_ & ~\quotient[56] ;
  assign new_n1002_ = ~new_n806_ & new_n891_;
  assign new_n1003_ = ~new_n887_ & new_n1002_;
  assign new_n1004_ = ~new_n888_ & ~new_n891_;
  assign new_n1005_ = ~new_n1003_ & ~new_n1004_;
  assign new_n1006_ = \quotient[56]  & ~new_n1005_;
  assign new_n1007_ = ~new_n1001_ & ~new_n1006_;
  assign new_n1008_ = ~\b[8]  & ~new_n1007_;
  assign new_n1009_ = \b[8]  & ~new_n1001_;
  assign new_n1010_ = ~new_n1006_ & new_n1009_;
  assign new_n1011_ = new_n378_ & new_n392_;
  assign new_n1012_ = new_n424_ & new_n1011_;
  assign new_n1013_ = ~new_n1010_ & new_n1012_;
  assign new_n1014_ = ~new_n1008_ & new_n1013_;
  assign new_n1015_ = ~new_n1000_ & new_n1014_;
  assign new_n1016_ = new_n895_ & ~new_n1007_;
  assign \quotient[55]  = new_n1015_ | new_n1016_;
  assign new_n1018_ = ~new_n914_ & new_n998_;
  assign new_n1019_ = ~new_n994_ & new_n1018_;
  assign new_n1020_ = ~new_n995_ & ~new_n998_;
  assign new_n1021_ = ~new_n1019_ & ~new_n1020_;
  assign new_n1022_ = \quotient[55]  & ~new_n1021_;
  assign new_n1023_ = ~new_n904_ & ~new_n1016_;
  assign new_n1024_ = ~new_n1015_ & new_n1023_;
  assign new_n1025_ = ~new_n1022_ & ~new_n1024_;
  assign new_n1026_ = ~new_n905_ & ~new_n1010_;
  assign new_n1027_ = ~new_n1008_ & new_n1026_;
  assign new_n1028_ = ~new_n999_ & new_n1027_;
  assign new_n1029_ = ~new_n1008_ & ~new_n1010_;
  assign new_n1030_ = ~new_n1000_ & ~new_n1029_;
  assign new_n1031_ = ~new_n1028_ & ~new_n1030_;
  assign new_n1032_ = \quotient[55]  & ~new_n1031_;
  assign new_n1033_ = ~new_n1007_ & ~new_n1016_;
  assign new_n1034_ = ~new_n1015_ & new_n1033_;
  assign new_n1035_ = ~new_n1032_ & ~new_n1034_;
  assign new_n1036_ = ~\b[9]  & ~new_n1035_;
  assign new_n1037_ = ~\b[8]  & ~new_n1025_;
  assign new_n1038_ = ~new_n923_ & new_n993_;
  assign new_n1039_ = ~new_n989_ & new_n1038_;
  assign new_n1040_ = ~new_n990_ & ~new_n993_;
  assign new_n1041_ = ~new_n1039_ & ~new_n1040_;
  assign new_n1042_ = \quotient[55]  & ~new_n1041_;
  assign new_n1043_ = ~new_n913_ & ~new_n1016_;
  assign new_n1044_ = ~new_n1015_ & new_n1043_;
  assign new_n1045_ = ~new_n1042_ & ~new_n1044_;
  assign new_n1046_ = ~\b[7]  & ~new_n1045_;
  assign new_n1047_ = ~new_n932_ & new_n988_;
  assign new_n1048_ = ~new_n984_ & new_n1047_;
  assign new_n1049_ = ~new_n985_ & ~new_n988_;
  assign new_n1050_ = ~new_n1048_ & ~new_n1049_;
  assign new_n1051_ = \quotient[55]  & ~new_n1050_;
  assign new_n1052_ = ~new_n922_ & ~new_n1016_;
  assign new_n1053_ = ~new_n1015_ & new_n1052_;
  assign new_n1054_ = ~new_n1051_ & ~new_n1053_;
  assign new_n1055_ = ~\b[6]  & ~new_n1054_;
  assign new_n1056_ = ~new_n941_ & new_n983_;
  assign new_n1057_ = ~new_n979_ & new_n1056_;
  assign new_n1058_ = ~new_n980_ & ~new_n983_;
  assign new_n1059_ = ~new_n1057_ & ~new_n1058_;
  assign new_n1060_ = \quotient[55]  & ~new_n1059_;
  assign new_n1061_ = ~new_n931_ & ~new_n1016_;
  assign new_n1062_ = ~new_n1015_ & new_n1061_;
  assign new_n1063_ = ~new_n1060_ & ~new_n1062_;
  assign new_n1064_ = ~\b[5]  & ~new_n1063_;
  assign new_n1065_ = ~new_n949_ & new_n978_;
  assign new_n1066_ = ~new_n974_ & new_n1065_;
  assign new_n1067_ = ~new_n975_ & ~new_n978_;
  assign new_n1068_ = ~new_n1066_ & ~new_n1067_;
  assign new_n1069_ = \quotient[55]  & ~new_n1068_;
  assign new_n1070_ = ~new_n940_ & ~new_n1016_;
  assign new_n1071_ = ~new_n1015_ & new_n1070_;
  assign new_n1072_ = ~new_n1069_ & ~new_n1071_;
  assign new_n1073_ = ~\b[4]  & ~new_n1072_;
  assign new_n1074_ = ~new_n969_ & new_n973_;
  assign new_n1075_ = ~new_n968_ & new_n1074_;
  assign new_n1076_ = ~new_n970_ & ~new_n973_;
  assign new_n1077_ = ~new_n1075_ & ~new_n1076_;
  assign new_n1078_ = \quotient[55]  & ~new_n1077_;
  assign new_n1079_ = ~new_n948_ & ~new_n1016_;
  assign new_n1080_ = ~new_n1015_ & new_n1079_;
  assign new_n1081_ = ~new_n1078_ & ~new_n1080_;
  assign new_n1082_ = ~\b[3]  & ~new_n1081_;
  assign new_n1083_ = ~new_n965_ & new_n967_;
  assign new_n1084_ = ~new_n963_ & new_n1083_;
  assign new_n1085_ = ~new_n968_ & ~new_n1084_;
  assign new_n1086_ = \quotient[55]  & new_n1085_;
  assign new_n1087_ = ~new_n962_ & ~new_n1016_;
  assign new_n1088_ = ~new_n1015_ & new_n1087_;
  assign new_n1089_ = ~new_n1086_ & ~new_n1088_;
  assign new_n1090_ = ~\b[2]  & ~new_n1089_;
  assign new_n1091_ = \b[0]  & \quotient[55] ;
  assign new_n1092_ = \a[55]  & ~new_n1091_;
  assign new_n1093_ = new_n967_ & \quotient[55] ;
  assign new_n1094_ = ~new_n1092_ & ~new_n1093_;
  assign new_n1095_ = \b[1]  & ~new_n1094_;
  assign new_n1096_ = ~\b[1]  & ~new_n1093_;
  assign new_n1097_ = ~new_n1092_ & new_n1096_;
  assign new_n1098_ = ~new_n1095_ & ~new_n1097_;
  assign new_n1099_ = ~\a[54]  & \b[0] ;
  assign new_n1100_ = ~new_n1098_ & ~new_n1099_;
  assign new_n1101_ = ~\b[1]  & ~new_n1094_;
  assign new_n1102_ = ~new_n1100_ & ~new_n1101_;
  assign new_n1103_ = \b[2]  & ~new_n1088_;
  assign new_n1104_ = ~new_n1086_ & new_n1103_;
  assign new_n1105_ = ~new_n1090_ & ~new_n1104_;
  assign new_n1106_ = ~new_n1102_ & new_n1105_;
  assign new_n1107_ = ~new_n1090_ & ~new_n1106_;
  assign new_n1108_ = \b[3]  & ~new_n1080_;
  assign new_n1109_ = ~new_n1078_ & new_n1108_;
  assign new_n1110_ = ~new_n1082_ & ~new_n1109_;
  assign new_n1111_ = ~new_n1107_ & new_n1110_;
  assign new_n1112_ = ~new_n1082_ & ~new_n1111_;
  assign new_n1113_ = \b[4]  & ~new_n1071_;
  assign new_n1114_ = ~new_n1069_ & new_n1113_;
  assign new_n1115_ = ~new_n1073_ & ~new_n1114_;
  assign new_n1116_ = ~new_n1112_ & new_n1115_;
  assign new_n1117_ = ~new_n1073_ & ~new_n1116_;
  assign new_n1118_ = \b[5]  & ~new_n1062_;
  assign new_n1119_ = ~new_n1060_ & new_n1118_;
  assign new_n1120_ = ~new_n1064_ & ~new_n1119_;
  assign new_n1121_ = ~new_n1117_ & new_n1120_;
  assign new_n1122_ = ~new_n1064_ & ~new_n1121_;
  assign new_n1123_ = \b[6]  & ~new_n1053_;
  assign new_n1124_ = ~new_n1051_ & new_n1123_;
  assign new_n1125_ = ~new_n1055_ & ~new_n1124_;
  assign new_n1126_ = ~new_n1122_ & new_n1125_;
  assign new_n1127_ = ~new_n1055_ & ~new_n1126_;
  assign new_n1128_ = \b[7]  & ~new_n1044_;
  assign new_n1129_ = ~new_n1042_ & new_n1128_;
  assign new_n1130_ = ~new_n1046_ & ~new_n1129_;
  assign new_n1131_ = ~new_n1127_ & new_n1130_;
  assign new_n1132_ = ~new_n1046_ & ~new_n1131_;
  assign new_n1133_ = \b[8]  & ~new_n1024_;
  assign new_n1134_ = ~new_n1022_ & new_n1133_;
  assign new_n1135_ = ~new_n1037_ & ~new_n1134_;
  assign new_n1136_ = ~new_n1132_ & new_n1135_;
  assign new_n1137_ = ~new_n1037_ & ~new_n1136_;
  assign new_n1138_ = \b[9]  & ~new_n1034_;
  assign new_n1139_ = ~new_n1032_ & new_n1138_;
  assign new_n1140_ = ~new_n1036_ & ~new_n1139_;
  assign new_n1141_ = ~new_n1137_ & new_n1140_;
  assign new_n1142_ = ~new_n1036_ & ~new_n1141_;
  assign new_n1143_ = new_n263_ & new_n274_;
  assign new_n1144_ = new_n344_ & new_n1143_;
  assign new_n1145_ = new_n432_ & new_n1144_;
  assign \quotient[54]  = ~new_n1142_ & new_n1145_;
  assign new_n1147_ = ~new_n1025_ & ~\quotient[54] ;
  assign new_n1148_ = ~new_n1046_ & new_n1135_;
  assign new_n1149_ = ~new_n1131_ & new_n1148_;
  assign new_n1150_ = ~new_n1132_ & ~new_n1135_;
  assign new_n1151_ = ~new_n1149_ & ~new_n1150_;
  assign new_n1152_ = new_n1145_ & ~new_n1151_;
  assign new_n1153_ = ~new_n1142_ & new_n1152_;
  assign new_n1154_ = ~new_n1147_ & ~new_n1153_;
  assign new_n1155_ = ~new_n1035_ & ~\quotient[54] ;
  assign new_n1156_ = ~new_n1037_ & new_n1140_;
  assign new_n1157_ = ~new_n1136_ & new_n1156_;
  assign new_n1158_ = ~new_n1137_ & ~new_n1140_;
  assign new_n1159_ = ~new_n1157_ & ~new_n1158_;
  assign new_n1160_ = \quotient[54]  & ~new_n1159_;
  assign new_n1161_ = ~new_n1155_ & ~new_n1160_;
  assign new_n1162_ = ~\b[10]  & ~new_n1161_;
  assign new_n1163_ = ~\b[9]  & ~new_n1154_;
  assign new_n1164_ = ~new_n1045_ & ~\quotient[54] ;
  assign new_n1165_ = ~new_n1055_ & new_n1130_;
  assign new_n1166_ = ~new_n1126_ & new_n1165_;
  assign new_n1167_ = ~new_n1127_ & ~new_n1130_;
  assign new_n1168_ = ~new_n1166_ & ~new_n1167_;
  assign new_n1169_ = new_n1145_ & ~new_n1168_;
  assign new_n1170_ = ~new_n1142_ & new_n1169_;
  assign new_n1171_ = ~new_n1164_ & ~new_n1170_;
  assign new_n1172_ = ~\b[8]  & ~new_n1171_;
  assign new_n1173_ = ~new_n1054_ & ~\quotient[54] ;
  assign new_n1174_ = ~new_n1064_ & new_n1125_;
  assign new_n1175_ = ~new_n1121_ & new_n1174_;
  assign new_n1176_ = ~new_n1122_ & ~new_n1125_;
  assign new_n1177_ = ~new_n1175_ & ~new_n1176_;
  assign new_n1178_ = new_n1145_ & ~new_n1177_;
  assign new_n1179_ = ~new_n1142_ & new_n1178_;
  assign new_n1180_ = ~new_n1173_ & ~new_n1179_;
  assign new_n1181_ = ~\b[7]  & ~new_n1180_;
  assign new_n1182_ = ~new_n1063_ & ~\quotient[54] ;
  assign new_n1183_ = ~new_n1073_ & new_n1120_;
  assign new_n1184_ = ~new_n1116_ & new_n1183_;
  assign new_n1185_ = ~new_n1117_ & ~new_n1120_;
  assign new_n1186_ = ~new_n1184_ & ~new_n1185_;
  assign new_n1187_ = new_n1145_ & ~new_n1186_;
  assign new_n1188_ = ~new_n1142_ & new_n1187_;
  assign new_n1189_ = ~new_n1182_ & ~new_n1188_;
  assign new_n1190_ = ~\b[6]  & ~new_n1189_;
  assign new_n1191_ = ~new_n1072_ & ~\quotient[54] ;
  assign new_n1192_ = ~new_n1082_ & new_n1115_;
  assign new_n1193_ = ~new_n1111_ & new_n1192_;
  assign new_n1194_ = ~new_n1112_ & ~new_n1115_;
  assign new_n1195_ = ~new_n1193_ & ~new_n1194_;
  assign new_n1196_ = new_n1145_ & ~new_n1195_;
  assign new_n1197_ = ~new_n1142_ & new_n1196_;
  assign new_n1198_ = ~new_n1191_ & ~new_n1197_;
  assign new_n1199_ = ~\b[5]  & ~new_n1198_;
  assign new_n1200_ = ~new_n1081_ & ~\quotient[54] ;
  assign new_n1201_ = ~new_n1090_ & new_n1110_;
  assign new_n1202_ = ~new_n1106_ & new_n1201_;
  assign new_n1203_ = ~new_n1107_ & ~new_n1110_;
  assign new_n1204_ = ~new_n1202_ & ~new_n1203_;
  assign new_n1205_ = new_n1145_ & ~new_n1204_;
  assign new_n1206_ = ~new_n1142_ & new_n1205_;
  assign new_n1207_ = ~new_n1200_ & ~new_n1206_;
  assign new_n1208_ = ~\b[4]  & ~new_n1207_;
  assign new_n1209_ = ~new_n1089_ & ~\quotient[54] ;
  assign new_n1210_ = ~new_n1101_ & new_n1105_;
  assign new_n1211_ = ~new_n1100_ & new_n1210_;
  assign new_n1212_ = ~new_n1102_ & ~new_n1105_;
  assign new_n1213_ = ~new_n1211_ & ~new_n1212_;
  assign new_n1214_ = new_n1145_ & ~new_n1213_;
  assign new_n1215_ = ~new_n1142_ & new_n1214_;
  assign new_n1216_ = ~new_n1209_ & ~new_n1215_;
  assign new_n1217_ = ~\b[3]  & ~new_n1216_;
  assign new_n1218_ = ~new_n1094_ & ~\quotient[54] ;
  assign new_n1219_ = ~new_n1097_ & new_n1099_;
  assign new_n1220_ = ~new_n1095_ & new_n1219_;
  assign new_n1221_ = new_n1145_ & ~new_n1220_;
  assign new_n1222_ = ~new_n1100_ & new_n1221_;
  assign new_n1223_ = ~new_n1142_ & new_n1222_;
  assign new_n1224_ = ~new_n1218_ & ~new_n1223_;
  assign new_n1225_ = ~\b[2]  & ~new_n1224_;
  assign new_n1226_ = \b[0]  & ~\b[10] ;
  assign new_n1227_ = new_n390_ & new_n1226_;
  assign new_n1228_ = new_n388_ & new_n1227_;
  assign new_n1229_ = new_n378_ & new_n1228_;
  assign new_n1230_ = new_n424_ & new_n1229_;
  assign new_n1231_ = ~new_n1142_ & new_n1230_;
  assign new_n1232_ = \a[54]  & ~new_n1231_;
  assign new_n1233_ = new_n263_ & new_n1099_;
  assign new_n1234_ = new_n274_ & new_n1233_;
  assign new_n1235_ = new_n344_ & new_n1234_;
  assign new_n1236_ = new_n432_ & new_n1235_;
  assign new_n1237_ = ~new_n1142_ & new_n1236_;
  assign new_n1238_ = ~new_n1232_ & ~new_n1237_;
  assign new_n1239_ = \b[1]  & ~new_n1238_;
  assign new_n1240_ = ~\b[1]  & ~new_n1237_;
  assign new_n1241_ = ~new_n1232_ & new_n1240_;
  assign new_n1242_ = ~new_n1239_ & ~new_n1241_;
  assign new_n1243_ = ~\a[53]  & \b[0] ;
  assign new_n1244_ = ~new_n1242_ & ~new_n1243_;
  assign new_n1245_ = ~\b[1]  & ~new_n1238_;
  assign new_n1246_ = ~new_n1244_ & ~new_n1245_;
  assign new_n1247_ = \b[2]  & ~new_n1223_;
  assign new_n1248_ = ~new_n1218_ & new_n1247_;
  assign new_n1249_ = ~new_n1225_ & ~new_n1248_;
  assign new_n1250_ = ~new_n1246_ & new_n1249_;
  assign new_n1251_ = ~new_n1225_ & ~new_n1250_;
  assign new_n1252_ = \b[3]  & ~new_n1215_;
  assign new_n1253_ = ~new_n1209_ & new_n1252_;
  assign new_n1254_ = ~new_n1217_ & ~new_n1253_;
  assign new_n1255_ = ~new_n1251_ & new_n1254_;
  assign new_n1256_ = ~new_n1217_ & ~new_n1255_;
  assign new_n1257_ = \b[4]  & ~new_n1206_;
  assign new_n1258_ = ~new_n1200_ & new_n1257_;
  assign new_n1259_ = ~new_n1208_ & ~new_n1258_;
  assign new_n1260_ = ~new_n1256_ & new_n1259_;
  assign new_n1261_ = ~new_n1208_ & ~new_n1260_;
  assign new_n1262_ = \b[5]  & ~new_n1197_;
  assign new_n1263_ = ~new_n1191_ & new_n1262_;
  assign new_n1264_ = ~new_n1199_ & ~new_n1263_;
  assign new_n1265_ = ~new_n1261_ & new_n1264_;
  assign new_n1266_ = ~new_n1199_ & ~new_n1265_;
  assign new_n1267_ = \b[6]  & ~new_n1188_;
  assign new_n1268_ = ~new_n1182_ & new_n1267_;
  assign new_n1269_ = ~new_n1190_ & ~new_n1268_;
  assign new_n1270_ = ~new_n1266_ & new_n1269_;
  assign new_n1271_ = ~new_n1190_ & ~new_n1270_;
  assign new_n1272_ = \b[7]  & ~new_n1179_;
  assign new_n1273_ = ~new_n1173_ & new_n1272_;
  assign new_n1274_ = ~new_n1181_ & ~new_n1273_;
  assign new_n1275_ = ~new_n1271_ & new_n1274_;
  assign new_n1276_ = ~new_n1181_ & ~new_n1275_;
  assign new_n1277_ = \b[8]  & ~new_n1170_;
  assign new_n1278_ = ~new_n1164_ & new_n1277_;
  assign new_n1279_ = ~new_n1172_ & ~new_n1278_;
  assign new_n1280_ = ~new_n1276_ & new_n1279_;
  assign new_n1281_ = ~new_n1172_ & ~new_n1280_;
  assign new_n1282_ = \b[9]  & ~new_n1153_;
  assign new_n1283_ = ~new_n1147_ & new_n1282_;
  assign new_n1284_ = ~new_n1163_ & ~new_n1283_;
  assign new_n1285_ = ~new_n1281_ & new_n1284_;
  assign new_n1286_ = ~new_n1163_ & ~new_n1285_;
  assign new_n1287_ = \b[10]  & ~new_n1155_;
  assign new_n1288_ = ~new_n1160_ & new_n1287_;
  assign new_n1289_ = ~new_n1162_ & ~new_n1288_;
  assign new_n1290_ = ~new_n1286_ & new_n1289_;
  assign new_n1291_ = ~new_n1162_ & ~new_n1290_;
  assign new_n1292_ = new_n388_ & new_n390_;
  assign new_n1293_ = new_n378_ & new_n1292_;
  assign new_n1294_ = new_n424_ & new_n1293_;
  assign \quotient[53]  = ~new_n1291_ & new_n1294_;
  assign new_n1296_ = ~new_n1154_ & ~\quotient[53] ;
  assign new_n1297_ = ~new_n1172_ & new_n1284_;
  assign new_n1298_ = ~new_n1280_ & new_n1297_;
  assign new_n1299_ = ~new_n1281_ & ~new_n1284_;
  assign new_n1300_ = ~new_n1298_ & ~new_n1299_;
  assign new_n1301_ = new_n1294_ & ~new_n1300_;
  assign new_n1302_ = ~new_n1291_ & new_n1301_;
  assign new_n1303_ = ~new_n1296_ & ~new_n1302_;
  assign new_n1304_ = ~\b[10]  & ~new_n1303_;
  assign new_n1305_ = ~new_n1171_ & ~\quotient[53] ;
  assign new_n1306_ = ~new_n1181_ & new_n1279_;
  assign new_n1307_ = ~new_n1275_ & new_n1306_;
  assign new_n1308_ = ~new_n1276_ & ~new_n1279_;
  assign new_n1309_ = ~new_n1307_ & ~new_n1308_;
  assign new_n1310_ = new_n1294_ & ~new_n1309_;
  assign new_n1311_ = ~new_n1291_ & new_n1310_;
  assign new_n1312_ = ~new_n1305_ & ~new_n1311_;
  assign new_n1313_ = ~\b[9]  & ~new_n1312_;
  assign new_n1314_ = ~new_n1180_ & ~\quotient[53] ;
  assign new_n1315_ = ~new_n1190_ & new_n1274_;
  assign new_n1316_ = ~new_n1270_ & new_n1315_;
  assign new_n1317_ = ~new_n1271_ & ~new_n1274_;
  assign new_n1318_ = ~new_n1316_ & ~new_n1317_;
  assign new_n1319_ = new_n1294_ & ~new_n1318_;
  assign new_n1320_ = ~new_n1291_ & new_n1319_;
  assign new_n1321_ = ~new_n1314_ & ~new_n1320_;
  assign new_n1322_ = ~\b[8]  & ~new_n1321_;
  assign new_n1323_ = ~new_n1189_ & ~\quotient[53] ;
  assign new_n1324_ = ~new_n1199_ & new_n1269_;
  assign new_n1325_ = ~new_n1265_ & new_n1324_;
  assign new_n1326_ = ~new_n1266_ & ~new_n1269_;
  assign new_n1327_ = ~new_n1325_ & ~new_n1326_;
  assign new_n1328_ = new_n1294_ & ~new_n1327_;
  assign new_n1329_ = ~new_n1291_ & new_n1328_;
  assign new_n1330_ = ~new_n1323_ & ~new_n1329_;
  assign new_n1331_ = ~\b[7]  & ~new_n1330_;
  assign new_n1332_ = ~new_n1198_ & ~\quotient[53] ;
  assign new_n1333_ = ~new_n1208_ & new_n1264_;
  assign new_n1334_ = ~new_n1260_ & new_n1333_;
  assign new_n1335_ = ~new_n1261_ & ~new_n1264_;
  assign new_n1336_ = ~new_n1334_ & ~new_n1335_;
  assign new_n1337_ = new_n1294_ & ~new_n1336_;
  assign new_n1338_ = ~new_n1291_ & new_n1337_;
  assign new_n1339_ = ~new_n1332_ & ~new_n1338_;
  assign new_n1340_ = ~\b[6]  & ~new_n1339_;
  assign new_n1341_ = ~new_n1207_ & ~\quotient[53] ;
  assign new_n1342_ = ~new_n1217_ & new_n1259_;
  assign new_n1343_ = ~new_n1255_ & new_n1342_;
  assign new_n1344_ = ~new_n1256_ & ~new_n1259_;
  assign new_n1345_ = ~new_n1343_ & ~new_n1344_;
  assign new_n1346_ = new_n1294_ & ~new_n1345_;
  assign new_n1347_ = ~new_n1291_ & new_n1346_;
  assign new_n1348_ = ~new_n1341_ & ~new_n1347_;
  assign new_n1349_ = ~\b[5]  & ~new_n1348_;
  assign new_n1350_ = ~new_n1216_ & ~\quotient[53] ;
  assign new_n1351_ = ~new_n1225_ & new_n1254_;
  assign new_n1352_ = ~new_n1250_ & new_n1351_;
  assign new_n1353_ = ~new_n1251_ & ~new_n1254_;
  assign new_n1354_ = ~new_n1352_ & ~new_n1353_;
  assign new_n1355_ = new_n1294_ & ~new_n1354_;
  assign new_n1356_ = ~new_n1291_ & new_n1355_;
  assign new_n1357_ = ~new_n1350_ & ~new_n1356_;
  assign new_n1358_ = ~\b[4]  & ~new_n1357_;
  assign new_n1359_ = ~new_n1224_ & ~\quotient[53] ;
  assign new_n1360_ = ~new_n1245_ & new_n1249_;
  assign new_n1361_ = ~new_n1244_ & new_n1360_;
  assign new_n1362_ = ~new_n1246_ & ~new_n1249_;
  assign new_n1363_ = ~new_n1361_ & ~new_n1362_;
  assign new_n1364_ = new_n1294_ & ~new_n1363_;
  assign new_n1365_ = ~new_n1291_ & new_n1364_;
  assign new_n1366_ = ~new_n1359_ & ~new_n1365_;
  assign new_n1367_ = ~\b[3]  & ~new_n1366_;
  assign new_n1368_ = ~new_n1238_ & ~\quotient[53] ;
  assign new_n1369_ = ~new_n1241_ & new_n1243_;
  assign new_n1370_ = ~new_n1239_ & new_n1369_;
  assign new_n1371_ = new_n1294_ & ~new_n1370_;
  assign new_n1372_ = ~new_n1244_ & new_n1371_;
  assign new_n1373_ = ~new_n1291_ & new_n1372_;
  assign new_n1374_ = ~new_n1368_ & ~new_n1373_;
  assign new_n1375_ = ~\b[2]  & ~new_n1374_;
  assign new_n1376_ = \b[0]  & ~\b[11] ;
  assign new_n1377_ = new_n274_ & new_n1376_;
  assign new_n1378_ = new_n344_ & new_n1377_;
  assign new_n1379_ = new_n432_ & new_n1378_;
  assign new_n1380_ = ~new_n1291_ & new_n1379_;
  assign new_n1381_ = \a[53]  & ~new_n1380_;
  assign new_n1382_ = new_n390_ & new_n1243_;
  assign new_n1383_ = new_n388_ & new_n1382_;
  assign new_n1384_ = new_n378_ & new_n1383_;
  assign new_n1385_ = new_n424_ & new_n1384_;
  assign new_n1386_ = ~new_n1291_ & new_n1385_;
  assign new_n1387_ = ~new_n1381_ & ~new_n1386_;
  assign new_n1388_ = \b[1]  & ~new_n1387_;
  assign new_n1389_ = ~\b[1]  & ~new_n1386_;
  assign new_n1390_ = ~new_n1381_ & new_n1389_;
  assign new_n1391_ = ~new_n1388_ & ~new_n1390_;
  assign new_n1392_ = ~\a[52]  & \b[0] ;
  assign new_n1393_ = ~new_n1391_ & ~new_n1392_;
  assign new_n1394_ = ~\b[1]  & ~new_n1387_;
  assign new_n1395_ = ~new_n1393_ & ~new_n1394_;
  assign new_n1396_ = \b[2]  & ~new_n1373_;
  assign new_n1397_ = ~new_n1368_ & new_n1396_;
  assign new_n1398_ = ~new_n1375_ & ~new_n1397_;
  assign new_n1399_ = ~new_n1395_ & new_n1398_;
  assign new_n1400_ = ~new_n1375_ & ~new_n1399_;
  assign new_n1401_ = \b[3]  & ~new_n1365_;
  assign new_n1402_ = ~new_n1359_ & new_n1401_;
  assign new_n1403_ = ~new_n1367_ & ~new_n1402_;
  assign new_n1404_ = ~new_n1400_ & new_n1403_;
  assign new_n1405_ = ~new_n1367_ & ~new_n1404_;
  assign new_n1406_ = \b[4]  & ~new_n1356_;
  assign new_n1407_ = ~new_n1350_ & new_n1406_;
  assign new_n1408_ = ~new_n1358_ & ~new_n1407_;
  assign new_n1409_ = ~new_n1405_ & new_n1408_;
  assign new_n1410_ = ~new_n1358_ & ~new_n1409_;
  assign new_n1411_ = \b[5]  & ~new_n1347_;
  assign new_n1412_ = ~new_n1341_ & new_n1411_;
  assign new_n1413_ = ~new_n1349_ & ~new_n1412_;
  assign new_n1414_ = ~new_n1410_ & new_n1413_;
  assign new_n1415_ = ~new_n1349_ & ~new_n1414_;
  assign new_n1416_ = \b[6]  & ~new_n1338_;
  assign new_n1417_ = ~new_n1332_ & new_n1416_;
  assign new_n1418_ = ~new_n1340_ & ~new_n1417_;
  assign new_n1419_ = ~new_n1415_ & new_n1418_;
  assign new_n1420_ = ~new_n1340_ & ~new_n1419_;
  assign new_n1421_ = \b[7]  & ~new_n1329_;
  assign new_n1422_ = ~new_n1323_ & new_n1421_;
  assign new_n1423_ = ~new_n1331_ & ~new_n1422_;
  assign new_n1424_ = ~new_n1420_ & new_n1423_;
  assign new_n1425_ = ~new_n1331_ & ~new_n1424_;
  assign new_n1426_ = \b[8]  & ~new_n1320_;
  assign new_n1427_ = ~new_n1314_ & new_n1426_;
  assign new_n1428_ = ~new_n1322_ & ~new_n1427_;
  assign new_n1429_ = ~new_n1425_ & new_n1428_;
  assign new_n1430_ = ~new_n1322_ & ~new_n1429_;
  assign new_n1431_ = \b[9]  & ~new_n1311_;
  assign new_n1432_ = ~new_n1305_ & new_n1431_;
  assign new_n1433_ = ~new_n1313_ & ~new_n1432_;
  assign new_n1434_ = ~new_n1430_ & new_n1433_;
  assign new_n1435_ = ~new_n1313_ & ~new_n1434_;
  assign new_n1436_ = \b[10]  & ~new_n1302_;
  assign new_n1437_ = ~new_n1296_ & new_n1436_;
  assign new_n1438_ = ~new_n1304_ & ~new_n1437_;
  assign new_n1439_ = ~new_n1435_ & new_n1438_;
  assign new_n1440_ = ~new_n1304_ & ~new_n1439_;
  assign new_n1441_ = ~new_n1161_ & ~\quotient[53] ;
  assign new_n1442_ = ~new_n1163_ & new_n1289_;
  assign new_n1443_ = ~new_n1285_ & new_n1442_;
  assign new_n1444_ = ~new_n1286_ & ~new_n1289_;
  assign new_n1445_ = ~new_n1443_ & ~new_n1444_;
  assign new_n1446_ = \quotient[53]  & ~new_n1445_;
  assign new_n1447_ = ~new_n1441_ & ~new_n1446_;
  assign new_n1448_ = ~\b[11]  & ~new_n1447_;
  assign new_n1449_ = \b[11]  & ~new_n1441_;
  assign new_n1450_ = ~new_n1446_ & new_n1449_;
  assign new_n1451_ = new_n275_ & new_n318_;
  assign new_n1452_ = new_n512_ & new_n1451_;
  assign new_n1453_ = ~new_n1450_ & new_n1452_;
  assign new_n1454_ = ~new_n1448_ & new_n1453_;
  assign new_n1455_ = ~new_n1440_ & new_n1454_;
  assign new_n1456_ = new_n1294_ & ~new_n1447_;
  assign \quotient[52]  = new_n1455_ | new_n1456_;
  assign new_n1458_ = ~new_n1313_ & new_n1438_;
  assign new_n1459_ = ~new_n1434_ & new_n1458_;
  assign new_n1460_ = ~new_n1435_ & ~new_n1438_;
  assign new_n1461_ = ~new_n1459_ & ~new_n1460_;
  assign new_n1462_ = \quotient[52]  & ~new_n1461_;
  assign new_n1463_ = ~new_n1303_ & ~new_n1456_;
  assign new_n1464_ = ~new_n1455_ & new_n1463_;
  assign new_n1465_ = ~new_n1462_ & ~new_n1464_;
  assign new_n1466_ = ~new_n1304_ & ~new_n1450_;
  assign new_n1467_ = ~new_n1448_ & new_n1466_;
  assign new_n1468_ = ~new_n1439_ & new_n1467_;
  assign new_n1469_ = ~new_n1448_ & ~new_n1450_;
  assign new_n1470_ = ~new_n1440_ & ~new_n1469_;
  assign new_n1471_ = ~new_n1468_ & ~new_n1470_;
  assign new_n1472_ = \quotient[52]  & ~new_n1471_;
  assign new_n1473_ = ~new_n1447_ & ~new_n1456_;
  assign new_n1474_ = ~new_n1455_ & new_n1473_;
  assign new_n1475_ = ~new_n1472_ & ~new_n1474_;
  assign new_n1476_ = ~\b[12]  & ~new_n1475_;
  assign new_n1477_ = ~\b[11]  & ~new_n1465_;
  assign new_n1478_ = ~new_n1322_ & new_n1433_;
  assign new_n1479_ = ~new_n1429_ & new_n1478_;
  assign new_n1480_ = ~new_n1430_ & ~new_n1433_;
  assign new_n1481_ = ~new_n1479_ & ~new_n1480_;
  assign new_n1482_ = \quotient[52]  & ~new_n1481_;
  assign new_n1483_ = ~new_n1312_ & ~new_n1456_;
  assign new_n1484_ = ~new_n1455_ & new_n1483_;
  assign new_n1485_ = ~new_n1482_ & ~new_n1484_;
  assign new_n1486_ = ~\b[10]  & ~new_n1485_;
  assign new_n1487_ = ~new_n1331_ & new_n1428_;
  assign new_n1488_ = ~new_n1424_ & new_n1487_;
  assign new_n1489_ = ~new_n1425_ & ~new_n1428_;
  assign new_n1490_ = ~new_n1488_ & ~new_n1489_;
  assign new_n1491_ = \quotient[52]  & ~new_n1490_;
  assign new_n1492_ = ~new_n1321_ & ~new_n1456_;
  assign new_n1493_ = ~new_n1455_ & new_n1492_;
  assign new_n1494_ = ~new_n1491_ & ~new_n1493_;
  assign new_n1495_ = ~\b[9]  & ~new_n1494_;
  assign new_n1496_ = ~new_n1340_ & new_n1423_;
  assign new_n1497_ = ~new_n1419_ & new_n1496_;
  assign new_n1498_ = ~new_n1420_ & ~new_n1423_;
  assign new_n1499_ = ~new_n1497_ & ~new_n1498_;
  assign new_n1500_ = \quotient[52]  & ~new_n1499_;
  assign new_n1501_ = ~new_n1330_ & ~new_n1456_;
  assign new_n1502_ = ~new_n1455_ & new_n1501_;
  assign new_n1503_ = ~new_n1500_ & ~new_n1502_;
  assign new_n1504_ = ~\b[8]  & ~new_n1503_;
  assign new_n1505_ = ~new_n1349_ & new_n1418_;
  assign new_n1506_ = ~new_n1414_ & new_n1505_;
  assign new_n1507_ = ~new_n1415_ & ~new_n1418_;
  assign new_n1508_ = ~new_n1506_ & ~new_n1507_;
  assign new_n1509_ = \quotient[52]  & ~new_n1508_;
  assign new_n1510_ = ~new_n1339_ & ~new_n1456_;
  assign new_n1511_ = ~new_n1455_ & new_n1510_;
  assign new_n1512_ = ~new_n1509_ & ~new_n1511_;
  assign new_n1513_ = ~\b[7]  & ~new_n1512_;
  assign new_n1514_ = ~new_n1358_ & new_n1413_;
  assign new_n1515_ = ~new_n1409_ & new_n1514_;
  assign new_n1516_ = ~new_n1410_ & ~new_n1413_;
  assign new_n1517_ = ~new_n1515_ & ~new_n1516_;
  assign new_n1518_ = \quotient[52]  & ~new_n1517_;
  assign new_n1519_ = ~new_n1348_ & ~new_n1456_;
  assign new_n1520_ = ~new_n1455_ & new_n1519_;
  assign new_n1521_ = ~new_n1518_ & ~new_n1520_;
  assign new_n1522_ = ~\b[6]  & ~new_n1521_;
  assign new_n1523_ = ~new_n1367_ & new_n1408_;
  assign new_n1524_ = ~new_n1404_ & new_n1523_;
  assign new_n1525_ = ~new_n1405_ & ~new_n1408_;
  assign new_n1526_ = ~new_n1524_ & ~new_n1525_;
  assign new_n1527_ = \quotient[52]  & ~new_n1526_;
  assign new_n1528_ = ~new_n1357_ & ~new_n1456_;
  assign new_n1529_ = ~new_n1455_ & new_n1528_;
  assign new_n1530_ = ~new_n1527_ & ~new_n1529_;
  assign new_n1531_ = ~\b[5]  & ~new_n1530_;
  assign new_n1532_ = ~new_n1375_ & new_n1403_;
  assign new_n1533_ = ~new_n1399_ & new_n1532_;
  assign new_n1534_ = ~new_n1400_ & ~new_n1403_;
  assign new_n1535_ = ~new_n1533_ & ~new_n1534_;
  assign new_n1536_ = \quotient[52]  & ~new_n1535_;
  assign new_n1537_ = ~new_n1366_ & ~new_n1456_;
  assign new_n1538_ = ~new_n1455_ & new_n1537_;
  assign new_n1539_ = ~new_n1536_ & ~new_n1538_;
  assign new_n1540_ = ~\b[4]  & ~new_n1539_;
  assign new_n1541_ = ~new_n1394_ & new_n1398_;
  assign new_n1542_ = ~new_n1393_ & new_n1541_;
  assign new_n1543_ = ~new_n1395_ & ~new_n1398_;
  assign new_n1544_ = ~new_n1542_ & ~new_n1543_;
  assign new_n1545_ = \quotient[52]  & ~new_n1544_;
  assign new_n1546_ = ~new_n1374_ & ~new_n1456_;
  assign new_n1547_ = ~new_n1455_ & new_n1546_;
  assign new_n1548_ = ~new_n1545_ & ~new_n1547_;
  assign new_n1549_ = ~\b[3]  & ~new_n1548_;
  assign new_n1550_ = ~new_n1390_ & new_n1392_;
  assign new_n1551_ = ~new_n1388_ & new_n1550_;
  assign new_n1552_ = ~new_n1393_ & ~new_n1551_;
  assign new_n1553_ = \quotient[52]  & new_n1552_;
  assign new_n1554_ = ~new_n1387_ & ~new_n1456_;
  assign new_n1555_ = ~new_n1455_ & new_n1554_;
  assign new_n1556_ = ~new_n1553_ & ~new_n1555_;
  assign new_n1557_ = ~\b[2]  & ~new_n1556_;
  assign new_n1558_ = \b[0]  & \quotient[52] ;
  assign new_n1559_ = \a[52]  & ~new_n1558_;
  assign new_n1560_ = new_n1392_ & \quotient[52] ;
  assign new_n1561_ = ~new_n1559_ & ~new_n1560_;
  assign new_n1562_ = \b[1]  & ~new_n1561_;
  assign new_n1563_ = ~\b[1]  & ~new_n1560_;
  assign new_n1564_ = ~new_n1559_ & new_n1563_;
  assign new_n1565_ = ~new_n1562_ & ~new_n1564_;
  assign new_n1566_ = ~\a[51]  & \b[0] ;
  assign new_n1567_ = ~new_n1565_ & ~new_n1566_;
  assign new_n1568_ = ~\b[1]  & ~new_n1561_;
  assign new_n1569_ = ~new_n1567_ & ~new_n1568_;
  assign new_n1570_ = \b[2]  & ~new_n1555_;
  assign new_n1571_ = ~new_n1553_ & new_n1570_;
  assign new_n1572_ = ~new_n1557_ & ~new_n1571_;
  assign new_n1573_ = ~new_n1569_ & new_n1572_;
  assign new_n1574_ = ~new_n1557_ & ~new_n1573_;
  assign new_n1575_ = \b[3]  & ~new_n1547_;
  assign new_n1576_ = ~new_n1545_ & new_n1575_;
  assign new_n1577_ = ~new_n1549_ & ~new_n1576_;
  assign new_n1578_ = ~new_n1574_ & new_n1577_;
  assign new_n1579_ = ~new_n1549_ & ~new_n1578_;
  assign new_n1580_ = \b[4]  & ~new_n1538_;
  assign new_n1581_ = ~new_n1536_ & new_n1580_;
  assign new_n1582_ = ~new_n1540_ & ~new_n1581_;
  assign new_n1583_ = ~new_n1579_ & new_n1582_;
  assign new_n1584_ = ~new_n1540_ & ~new_n1583_;
  assign new_n1585_ = \b[5]  & ~new_n1529_;
  assign new_n1586_ = ~new_n1527_ & new_n1585_;
  assign new_n1587_ = ~new_n1531_ & ~new_n1586_;
  assign new_n1588_ = ~new_n1584_ & new_n1587_;
  assign new_n1589_ = ~new_n1531_ & ~new_n1588_;
  assign new_n1590_ = \b[6]  & ~new_n1520_;
  assign new_n1591_ = ~new_n1518_ & new_n1590_;
  assign new_n1592_ = ~new_n1522_ & ~new_n1591_;
  assign new_n1593_ = ~new_n1589_ & new_n1592_;
  assign new_n1594_ = ~new_n1522_ & ~new_n1593_;
  assign new_n1595_ = \b[7]  & ~new_n1511_;
  assign new_n1596_ = ~new_n1509_ & new_n1595_;
  assign new_n1597_ = ~new_n1513_ & ~new_n1596_;
  assign new_n1598_ = ~new_n1594_ & new_n1597_;
  assign new_n1599_ = ~new_n1513_ & ~new_n1598_;
  assign new_n1600_ = \b[8]  & ~new_n1502_;
  assign new_n1601_ = ~new_n1500_ & new_n1600_;
  assign new_n1602_ = ~new_n1504_ & ~new_n1601_;
  assign new_n1603_ = ~new_n1599_ & new_n1602_;
  assign new_n1604_ = ~new_n1504_ & ~new_n1603_;
  assign new_n1605_ = \b[9]  & ~new_n1493_;
  assign new_n1606_ = ~new_n1491_ & new_n1605_;
  assign new_n1607_ = ~new_n1495_ & ~new_n1606_;
  assign new_n1608_ = ~new_n1604_ & new_n1607_;
  assign new_n1609_ = ~new_n1495_ & ~new_n1608_;
  assign new_n1610_ = \b[10]  & ~new_n1484_;
  assign new_n1611_ = ~new_n1482_ & new_n1610_;
  assign new_n1612_ = ~new_n1486_ & ~new_n1611_;
  assign new_n1613_ = ~new_n1609_ & new_n1612_;
  assign new_n1614_ = ~new_n1486_ & ~new_n1613_;
  assign new_n1615_ = \b[11]  & ~new_n1464_;
  assign new_n1616_ = ~new_n1462_ & new_n1615_;
  assign new_n1617_ = ~new_n1477_ & ~new_n1616_;
  assign new_n1618_ = ~new_n1614_ & new_n1617_;
  assign new_n1619_ = ~new_n1477_ & ~new_n1618_;
  assign new_n1620_ = \b[12]  & ~new_n1474_;
  assign new_n1621_ = ~new_n1472_ & new_n1620_;
  assign new_n1622_ = ~new_n1476_ & ~new_n1621_;
  assign new_n1623_ = ~new_n1619_ & new_n1622_;
  assign new_n1624_ = ~new_n1476_ & ~new_n1623_;
  assign new_n1625_ = new_n589_ & new_n591_;
  assign new_n1626_ = new_n599_ & new_n1625_;
  assign \quotient[51]  = ~new_n1624_ & new_n1626_;
  assign new_n1628_ = ~new_n1465_ & ~\quotient[51] ;
  assign new_n1629_ = ~new_n1486_ & new_n1617_;
  assign new_n1630_ = ~new_n1613_ & new_n1629_;
  assign new_n1631_ = ~new_n1614_ & ~new_n1617_;
  assign new_n1632_ = ~new_n1630_ & ~new_n1631_;
  assign new_n1633_ = new_n1626_ & ~new_n1632_;
  assign new_n1634_ = ~new_n1624_ & new_n1633_;
  assign new_n1635_ = ~new_n1628_ & ~new_n1634_;
  assign new_n1636_ = ~new_n1475_ & ~\quotient[51] ;
  assign new_n1637_ = ~new_n1477_ & new_n1622_;
  assign new_n1638_ = ~new_n1618_ & new_n1637_;
  assign new_n1639_ = ~new_n1619_ & ~new_n1622_;
  assign new_n1640_ = ~new_n1638_ & ~new_n1639_;
  assign new_n1641_ = \quotient[51]  & ~new_n1640_;
  assign new_n1642_ = ~new_n1636_ & ~new_n1641_;
  assign new_n1643_ = ~\b[13]  & ~new_n1642_;
  assign new_n1644_ = ~\b[12]  & ~new_n1635_;
  assign new_n1645_ = ~new_n1485_ & ~\quotient[51] ;
  assign new_n1646_ = ~new_n1495_ & new_n1612_;
  assign new_n1647_ = ~new_n1608_ & new_n1646_;
  assign new_n1648_ = ~new_n1609_ & ~new_n1612_;
  assign new_n1649_ = ~new_n1647_ & ~new_n1648_;
  assign new_n1650_ = new_n1626_ & ~new_n1649_;
  assign new_n1651_ = ~new_n1624_ & new_n1650_;
  assign new_n1652_ = ~new_n1645_ & ~new_n1651_;
  assign new_n1653_ = ~\b[11]  & ~new_n1652_;
  assign new_n1654_ = ~new_n1494_ & ~\quotient[51] ;
  assign new_n1655_ = ~new_n1504_ & new_n1607_;
  assign new_n1656_ = ~new_n1603_ & new_n1655_;
  assign new_n1657_ = ~new_n1604_ & ~new_n1607_;
  assign new_n1658_ = ~new_n1656_ & ~new_n1657_;
  assign new_n1659_ = new_n1626_ & ~new_n1658_;
  assign new_n1660_ = ~new_n1624_ & new_n1659_;
  assign new_n1661_ = ~new_n1654_ & ~new_n1660_;
  assign new_n1662_ = ~\b[10]  & ~new_n1661_;
  assign new_n1663_ = ~new_n1503_ & ~\quotient[51] ;
  assign new_n1664_ = ~new_n1513_ & new_n1602_;
  assign new_n1665_ = ~new_n1598_ & new_n1664_;
  assign new_n1666_ = ~new_n1599_ & ~new_n1602_;
  assign new_n1667_ = ~new_n1665_ & ~new_n1666_;
  assign new_n1668_ = new_n1626_ & ~new_n1667_;
  assign new_n1669_ = ~new_n1624_ & new_n1668_;
  assign new_n1670_ = ~new_n1663_ & ~new_n1669_;
  assign new_n1671_ = ~\b[9]  & ~new_n1670_;
  assign new_n1672_ = ~new_n1512_ & ~\quotient[51] ;
  assign new_n1673_ = ~new_n1522_ & new_n1597_;
  assign new_n1674_ = ~new_n1593_ & new_n1673_;
  assign new_n1675_ = ~new_n1594_ & ~new_n1597_;
  assign new_n1676_ = ~new_n1674_ & ~new_n1675_;
  assign new_n1677_ = new_n1626_ & ~new_n1676_;
  assign new_n1678_ = ~new_n1624_ & new_n1677_;
  assign new_n1679_ = ~new_n1672_ & ~new_n1678_;
  assign new_n1680_ = ~\b[8]  & ~new_n1679_;
  assign new_n1681_ = ~new_n1521_ & ~\quotient[51] ;
  assign new_n1682_ = ~new_n1531_ & new_n1592_;
  assign new_n1683_ = ~new_n1588_ & new_n1682_;
  assign new_n1684_ = ~new_n1589_ & ~new_n1592_;
  assign new_n1685_ = ~new_n1683_ & ~new_n1684_;
  assign new_n1686_ = new_n1626_ & ~new_n1685_;
  assign new_n1687_ = ~new_n1624_ & new_n1686_;
  assign new_n1688_ = ~new_n1681_ & ~new_n1687_;
  assign new_n1689_ = ~\b[7]  & ~new_n1688_;
  assign new_n1690_ = ~new_n1530_ & ~\quotient[51] ;
  assign new_n1691_ = ~new_n1540_ & new_n1587_;
  assign new_n1692_ = ~new_n1583_ & new_n1691_;
  assign new_n1693_ = ~new_n1584_ & ~new_n1587_;
  assign new_n1694_ = ~new_n1692_ & ~new_n1693_;
  assign new_n1695_ = new_n1626_ & ~new_n1694_;
  assign new_n1696_ = ~new_n1624_ & new_n1695_;
  assign new_n1697_ = ~new_n1690_ & ~new_n1696_;
  assign new_n1698_ = ~\b[6]  & ~new_n1697_;
  assign new_n1699_ = ~new_n1539_ & ~\quotient[51] ;
  assign new_n1700_ = ~new_n1549_ & new_n1582_;
  assign new_n1701_ = ~new_n1578_ & new_n1700_;
  assign new_n1702_ = ~new_n1579_ & ~new_n1582_;
  assign new_n1703_ = ~new_n1701_ & ~new_n1702_;
  assign new_n1704_ = new_n1626_ & ~new_n1703_;
  assign new_n1705_ = ~new_n1624_ & new_n1704_;
  assign new_n1706_ = ~new_n1699_ & ~new_n1705_;
  assign new_n1707_ = ~\b[5]  & ~new_n1706_;
  assign new_n1708_ = ~new_n1548_ & ~\quotient[51] ;
  assign new_n1709_ = ~new_n1557_ & new_n1577_;
  assign new_n1710_ = ~new_n1573_ & new_n1709_;
  assign new_n1711_ = ~new_n1574_ & ~new_n1577_;
  assign new_n1712_ = ~new_n1710_ & ~new_n1711_;
  assign new_n1713_ = new_n1626_ & ~new_n1712_;
  assign new_n1714_ = ~new_n1624_ & new_n1713_;
  assign new_n1715_ = ~new_n1708_ & ~new_n1714_;
  assign new_n1716_ = ~\b[4]  & ~new_n1715_;
  assign new_n1717_ = ~new_n1556_ & ~\quotient[51] ;
  assign new_n1718_ = ~new_n1568_ & new_n1572_;
  assign new_n1719_ = ~new_n1567_ & new_n1718_;
  assign new_n1720_ = ~new_n1569_ & ~new_n1572_;
  assign new_n1721_ = ~new_n1719_ & ~new_n1720_;
  assign new_n1722_ = new_n1626_ & ~new_n1721_;
  assign new_n1723_ = ~new_n1624_ & new_n1722_;
  assign new_n1724_ = ~new_n1717_ & ~new_n1723_;
  assign new_n1725_ = ~\b[3]  & ~new_n1724_;
  assign new_n1726_ = ~new_n1561_ & ~\quotient[51] ;
  assign new_n1727_ = ~new_n1564_ & new_n1566_;
  assign new_n1728_ = ~new_n1562_ & new_n1727_;
  assign new_n1729_ = new_n1626_ & ~new_n1728_;
  assign new_n1730_ = ~new_n1567_ & new_n1729_;
  assign new_n1731_ = ~new_n1624_ & new_n1730_;
  assign new_n1732_ = ~new_n1726_ & ~new_n1731_;
  assign new_n1733_ = ~\b[2]  & ~new_n1732_;
  assign new_n1734_ = \b[0]  & ~\b[13] ;
  assign new_n1735_ = new_n273_ & new_n1734_;
  assign new_n1736_ = new_n271_ & new_n1735_;
  assign new_n1737_ = new_n318_ & new_n1736_;
  assign new_n1738_ = new_n512_ & new_n1737_;
  assign new_n1739_ = ~new_n1624_ & new_n1738_;
  assign new_n1740_ = \a[51]  & ~new_n1739_;
  assign new_n1741_ = new_n388_ & new_n1566_;
  assign new_n1742_ = new_n378_ & new_n1741_;
  assign new_n1743_ = new_n424_ & new_n1742_;
  assign new_n1744_ = ~new_n1624_ & new_n1743_;
  assign new_n1745_ = ~new_n1740_ & ~new_n1744_;
  assign new_n1746_ = \b[1]  & ~new_n1745_;
  assign new_n1747_ = ~\b[1]  & ~new_n1744_;
  assign new_n1748_ = ~new_n1740_ & new_n1747_;
  assign new_n1749_ = ~new_n1746_ & ~new_n1748_;
  assign new_n1750_ = ~\a[50]  & \b[0] ;
  assign new_n1751_ = ~new_n1749_ & ~new_n1750_;
  assign new_n1752_ = ~\b[1]  & ~new_n1745_;
  assign new_n1753_ = ~new_n1751_ & ~new_n1752_;
  assign new_n1754_ = \b[2]  & ~new_n1731_;
  assign new_n1755_ = ~new_n1726_ & new_n1754_;
  assign new_n1756_ = ~new_n1733_ & ~new_n1755_;
  assign new_n1757_ = ~new_n1753_ & new_n1756_;
  assign new_n1758_ = ~new_n1733_ & ~new_n1757_;
  assign new_n1759_ = \b[3]  & ~new_n1723_;
  assign new_n1760_ = ~new_n1717_ & new_n1759_;
  assign new_n1761_ = ~new_n1725_ & ~new_n1760_;
  assign new_n1762_ = ~new_n1758_ & new_n1761_;
  assign new_n1763_ = ~new_n1725_ & ~new_n1762_;
  assign new_n1764_ = \b[4]  & ~new_n1714_;
  assign new_n1765_ = ~new_n1708_ & new_n1764_;
  assign new_n1766_ = ~new_n1716_ & ~new_n1765_;
  assign new_n1767_ = ~new_n1763_ & new_n1766_;
  assign new_n1768_ = ~new_n1716_ & ~new_n1767_;
  assign new_n1769_ = \b[5]  & ~new_n1705_;
  assign new_n1770_ = ~new_n1699_ & new_n1769_;
  assign new_n1771_ = ~new_n1707_ & ~new_n1770_;
  assign new_n1772_ = ~new_n1768_ & new_n1771_;
  assign new_n1773_ = ~new_n1707_ & ~new_n1772_;
  assign new_n1774_ = \b[6]  & ~new_n1696_;
  assign new_n1775_ = ~new_n1690_ & new_n1774_;
  assign new_n1776_ = ~new_n1698_ & ~new_n1775_;
  assign new_n1777_ = ~new_n1773_ & new_n1776_;
  assign new_n1778_ = ~new_n1698_ & ~new_n1777_;
  assign new_n1779_ = \b[7]  & ~new_n1687_;
  assign new_n1780_ = ~new_n1681_ & new_n1779_;
  assign new_n1781_ = ~new_n1689_ & ~new_n1780_;
  assign new_n1782_ = ~new_n1778_ & new_n1781_;
  assign new_n1783_ = ~new_n1689_ & ~new_n1782_;
  assign new_n1784_ = \b[8]  & ~new_n1678_;
  assign new_n1785_ = ~new_n1672_ & new_n1784_;
  assign new_n1786_ = ~new_n1680_ & ~new_n1785_;
  assign new_n1787_ = ~new_n1783_ & new_n1786_;
  assign new_n1788_ = ~new_n1680_ & ~new_n1787_;
  assign new_n1789_ = \b[9]  & ~new_n1669_;
  assign new_n1790_ = ~new_n1663_ & new_n1789_;
  assign new_n1791_ = ~new_n1671_ & ~new_n1790_;
  assign new_n1792_ = ~new_n1788_ & new_n1791_;
  assign new_n1793_ = ~new_n1671_ & ~new_n1792_;
  assign new_n1794_ = \b[10]  & ~new_n1660_;
  assign new_n1795_ = ~new_n1654_ & new_n1794_;
  assign new_n1796_ = ~new_n1662_ & ~new_n1795_;
  assign new_n1797_ = ~new_n1793_ & new_n1796_;
  assign new_n1798_ = ~new_n1662_ & ~new_n1797_;
  assign new_n1799_ = \b[11]  & ~new_n1651_;
  assign new_n1800_ = ~new_n1645_ & new_n1799_;
  assign new_n1801_ = ~new_n1653_ & ~new_n1800_;
  assign new_n1802_ = ~new_n1798_ & new_n1801_;
  assign new_n1803_ = ~new_n1653_ & ~new_n1802_;
  assign new_n1804_ = \b[12]  & ~new_n1634_;
  assign new_n1805_ = ~new_n1628_ & new_n1804_;
  assign new_n1806_ = ~new_n1644_ & ~new_n1805_;
  assign new_n1807_ = ~new_n1803_ & new_n1806_;
  assign new_n1808_ = ~new_n1644_ & ~new_n1807_;
  assign new_n1809_ = \b[13]  & ~new_n1636_;
  assign new_n1810_ = ~new_n1641_ & new_n1809_;
  assign new_n1811_ = ~new_n1643_ & ~new_n1810_;
  assign new_n1812_ = ~new_n1808_ & new_n1811_;
  assign new_n1813_ = ~new_n1643_ & ~new_n1812_;
  assign new_n1814_ = new_n271_ & new_n273_;
  assign new_n1815_ = new_n318_ & new_n1814_;
  assign new_n1816_ = new_n512_ & new_n1815_;
  assign \quotient[50]  = ~new_n1813_ & new_n1816_;
  assign new_n1818_ = ~new_n1635_ & ~\quotient[50] ;
  assign new_n1819_ = ~new_n1653_ & new_n1806_;
  assign new_n1820_ = ~new_n1802_ & new_n1819_;
  assign new_n1821_ = ~new_n1803_ & ~new_n1806_;
  assign new_n1822_ = ~new_n1820_ & ~new_n1821_;
  assign new_n1823_ = new_n1816_ & ~new_n1822_;
  assign new_n1824_ = ~new_n1813_ & new_n1823_;
  assign new_n1825_ = ~new_n1818_ & ~new_n1824_;
  assign new_n1826_ = ~\b[13]  & ~new_n1825_;
  assign new_n1827_ = ~new_n1652_ & ~\quotient[50] ;
  assign new_n1828_ = ~new_n1662_ & new_n1801_;
  assign new_n1829_ = ~new_n1797_ & new_n1828_;
  assign new_n1830_ = ~new_n1798_ & ~new_n1801_;
  assign new_n1831_ = ~new_n1829_ & ~new_n1830_;
  assign new_n1832_ = new_n1816_ & ~new_n1831_;
  assign new_n1833_ = ~new_n1813_ & new_n1832_;
  assign new_n1834_ = ~new_n1827_ & ~new_n1833_;
  assign new_n1835_ = ~\b[12]  & ~new_n1834_;
  assign new_n1836_ = ~new_n1661_ & ~\quotient[50] ;
  assign new_n1837_ = ~new_n1671_ & new_n1796_;
  assign new_n1838_ = ~new_n1792_ & new_n1837_;
  assign new_n1839_ = ~new_n1793_ & ~new_n1796_;
  assign new_n1840_ = ~new_n1838_ & ~new_n1839_;
  assign new_n1841_ = new_n1816_ & ~new_n1840_;
  assign new_n1842_ = ~new_n1813_ & new_n1841_;
  assign new_n1843_ = ~new_n1836_ & ~new_n1842_;
  assign new_n1844_ = ~\b[11]  & ~new_n1843_;
  assign new_n1845_ = ~new_n1670_ & ~\quotient[50] ;
  assign new_n1846_ = ~new_n1680_ & new_n1791_;
  assign new_n1847_ = ~new_n1787_ & new_n1846_;
  assign new_n1848_ = ~new_n1788_ & ~new_n1791_;
  assign new_n1849_ = ~new_n1847_ & ~new_n1848_;
  assign new_n1850_ = new_n1816_ & ~new_n1849_;
  assign new_n1851_ = ~new_n1813_ & new_n1850_;
  assign new_n1852_ = ~new_n1845_ & ~new_n1851_;
  assign new_n1853_ = ~\b[10]  & ~new_n1852_;
  assign new_n1854_ = ~new_n1679_ & ~\quotient[50] ;
  assign new_n1855_ = ~new_n1689_ & new_n1786_;
  assign new_n1856_ = ~new_n1782_ & new_n1855_;
  assign new_n1857_ = ~new_n1783_ & ~new_n1786_;
  assign new_n1858_ = ~new_n1856_ & ~new_n1857_;
  assign new_n1859_ = new_n1816_ & ~new_n1858_;
  assign new_n1860_ = ~new_n1813_ & new_n1859_;
  assign new_n1861_ = ~new_n1854_ & ~new_n1860_;
  assign new_n1862_ = ~\b[9]  & ~new_n1861_;
  assign new_n1863_ = ~new_n1688_ & ~\quotient[50] ;
  assign new_n1864_ = ~new_n1698_ & new_n1781_;
  assign new_n1865_ = ~new_n1777_ & new_n1864_;
  assign new_n1866_ = ~new_n1778_ & ~new_n1781_;
  assign new_n1867_ = ~new_n1865_ & ~new_n1866_;
  assign new_n1868_ = new_n1816_ & ~new_n1867_;
  assign new_n1869_ = ~new_n1813_ & new_n1868_;
  assign new_n1870_ = ~new_n1863_ & ~new_n1869_;
  assign new_n1871_ = ~\b[8]  & ~new_n1870_;
  assign new_n1872_ = ~new_n1697_ & ~\quotient[50] ;
  assign new_n1873_ = ~new_n1707_ & new_n1776_;
  assign new_n1874_ = ~new_n1772_ & new_n1873_;
  assign new_n1875_ = ~new_n1773_ & ~new_n1776_;
  assign new_n1876_ = ~new_n1874_ & ~new_n1875_;
  assign new_n1877_ = new_n1816_ & ~new_n1876_;
  assign new_n1878_ = ~new_n1813_ & new_n1877_;
  assign new_n1879_ = ~new_n1872_ & ~new_n1878_;
  assign new_n1880_ = ~\b[7]  & ~new_n1879_;
  assign new_n1881_ = ~new_n1706_ & ~\quotient[50] ;
  assign new_n1882_ = ~new_n1716_ & new_n1771_;
  assign new_n1883_ = ~new_n1767_ & new_n1882_;
  assign new_n1884_ = ~new_n1768_ & ~new_n1771_;
  assign new_n1885_ = ~new_n1883_ & ~new_n1884_;
  assign new_n1886_ = new_n1816_ & ~new_n1885_;
  assign new_n1887_ = ~new_n1813_ & new_n1886_;
  assign new_n1888_ = ~new_n1881_ & ~new_n1887_;
  assign new_n1889_ = ~\b[6]  & ~new_n1888_;
  assign new_n1890_ = ~new_n1715_ & ~\quotient[50] ;
  assign new_n1891_ = ~new_n1725_ & new_n1766_;
  assign new_n1892_ = ~new_n1762_ & new_n1891_;
  assign new_n1893_ = ~new_n1763_ & ~new_n1766_;
  assign new_n1894_ = ~new_n1892_ & ~new_n1893_;
  assign new_n1895_ = new_n1816_ & ~new_n1894_;
  assign new_n1896_ = ~new_n1813_ & new_n1895_;
  assign new_n1897_ = ~new_n1890_ & ~new_n1896_;
  assign new_n1898_ = ~\b[5]  & ~new_n1897_;
  assign new_n1899_ = ~new_n1724_ & ~\quotient[50] ;
  assign new_n1900_ = ~new_n1733_ & new_n1761_;
  assign new_n1901_ = ~new_n1757_ & new_n1900_;
  assign new_n1902_ = ~new_n1758_ & ~new_n1761_;
  assign new_n1903_ = ~new_n1901_ & ~new_n1902_;
  assign new_n1904_ = new_n1816_ & ~new_n1903_;
  assign new_n1905_ = ~new_n1813_ & new_n1904_;
  assign new_n1906_ = ~new_n1899_ & ~new_n1905_;
  assign new_n1907_ = ~\b[4]  & ~new_n1906_;
  assign new_n1908_ = ~new_n1732_ & ~\quotient[50] ;
  assign new_n1909_ = ~new_n1752_ & new_n1756_;
  assign new_n1910_ = ~new_n1751_ & new_n1909_;
  assign new_n1911_ = ~new_n1753_ & ~new_n1756_;
  assign new_n1912_ = ~new_n1910_ & ~new_n1911_;
  assign new_n1913_ = new_n1816_ & ~new_n1912_;
  assign new_n1914_ = ~new_n1813_ & new_n1913_;
  assign new_n1915_ = ~new_n1908_ & ~new_n1914_;
  assign new_n1916_ = ~\b[3]  & ~new_n1915_;
  assign new_n1917_ = ~new_n1745_ & ~\quotient[50] ;
  assign new_n1918_ = ~new_n1748_ & new_n1750_;
  assign new_n1919_ = ~new_n1746_ & new_n1918_;
  assign new_n1920_ = new_n1816_ & ~new_n1919_;
  assign new_n1921_ = ~new_n1751_ & new_n1920_;
  assign new_n1922_ = ~new_n1813_ & new_n1921_;
  assign new_n1923_ = ~new_n1917_ & ~new_n1922_;
  assign new_n1924_ = ~\b[2]  & ~new_n1923_;
  assign new_n1925_ = \b[0]  & ~\b[14] ;
  assign new_n1926_ = new_n387_ & new_n1925_;
  assign new_n1927_ = new_n369_ & new_n1926_;
  assign new_n1928_ = new_n589_ & new_n1927_;
  assign new_n1929_ = new_n599_ & new_n1928_;
  assign new_n1930_ = ~new_n1813_ & new_n1929_;
  assign new_n1931_ = \a[50]  & ~new_n1930_;
  assign new_n1932_ = new_n273_ & new_n1750_;
  assign new_n1933_ = new_n271_ & new_n1932_;
  assign new_n1934_ = new_n318_ & new_n1933_;
  assign new_n1935_ = new_n512_ & new_n1934_;
  assign new_n1936_ = ~new_n1813_ & new_n1935_;
  assign new_n1937_ = ~new_n1931_ & ~new_n1936_;
  assign new_n1938_ = \b[1]  & ~new_n1937_;
  assign new_n1939_ = ~\b[1]  & ~new_n1936_;
  assign new_n1940_ = ~new_n1931_ & new_n1939_;
  assign new_n1941_ = ~new_n1938_ & ~new_n1940_;
  assign new_n1942_ = ~\a[49]  & \b[0] ;
  assign new_n1943_ = ~new_n1941_ & ~new_n1942_;
  assign new_n1944_ = ~\b[1]  & ~new_n1937_;
  assign new_n1945_ = ~new_n1943_ & ~new_n1944_;
  assign new_n1946_ = \b[2]  & ~new_n1922_;
  assign new_n1947_ = ~new_n1917_ & new_n1946_;
  assign new_n1948_ = ~new_n1924_ & ~new_n1947_;
  assign new_n1949_ = ~new_n1945_ & new_n1948_;
  assign new_n1950_ = ~new_n1924_ & ~new_n1949_;
  assign new_n1951_ = \b[3]  & ~new_n1914_;
  assign new_n1952_ = ~new_n1908_ & new_n1951_;
  assign new_n1953_ = ~new_n1916_ & ~new_n1952_;
  assign new_n1954_ = ~new_n1950_ & new_n1953_;
  assign new_n1955_ = ~new_n1916_ & ~new_n1954_;
  assign new_n1956_ = \b[4]  & ~new_n1905_;
  assign new_n1957_ = ~new_n1899_ & new_n1956_;
  assign new_n1958_ = ~new_n1907_ & ~new_n1957_;
  assign new_n1959_ = ~new_n1955_ & new_n1958_;
  assign new_n1960_ = ~new_n1907_ & ~new_n1959_;
  assign new_n1961_ = \b[5]  & ~new_n1896_;
  assign new_n1962_ = ~new_n1890_ & new_n1961_;
  assign new_n1963_ = ~new_n1898_ & ~new_n1962_;
  assign new_n1964_ = ~new_n1960_ & new_n1963_;
  assign new_n1965_ = ~new_n1898_ & ~new_n1964_;
  assign new_n1966_ = \b[6]  & ~new_n1887_;
  assign new_n1967_ = ~new_n1881_ & new_n1966_;
  assign new_n1968_ = ~new_n1889_ & ~new_n1967_;
  assign new_n1969_ = ~new_n1965_ & new_n1968_;
  assign new_n1970_ = ~new_n1889_ & ~new_n1969_;
  assign new_n1971_ = \b[7]  & ~new_n1878_;
  assign new_n1972_ = ~new_n1872_ & new_n1971_;
  assign new_n1973_ = ~new_n1880_ & ~new_n1972_;
  assign new_n1974_ = ~new_n1970_ & new_n1973_;
  assign new_n1975_ = ~new_n1880_ & ~new_n1974_;
  assign new_n1976_ = \b[8]  & ~new_n1869_;
  assign new_n1977_ = ~new_n1863_ & new_n1976_;
  assign new_n1978_ = ~new_n1871_ & ~new_n1977_;
  assign new_n1979_ = ~new_n1975_ & new_n1978_;
  assign new_n1980_ = ~new_n1871_ & ~new_n1979_;
  assign new_n1981_ = \b[9]  & ~new_n1860_;
  assign new_n1982_ = ~new_n1854_ & new_n1981_;
  assign new_n1983_ = ~new_n1862_ & ~new_n1982_;
  assign new_n1984_ = ~new_n1980_ & new_n1983_;
  assign new_n1985_ = ~new_n1862_ & ~new_n1984_;
  assign new_n1986_ = \b[10]  & ~new_n1851_;
  assign new_n1987_ = ~new_n1845_ & new_n1986_;
  assign new_n1988_ = ~new_n1853_ & ~new_n1987_;
  assign new_n1989_ = ~new_n1985_ & new_n1988_;
  assign new_n1990_ = ~new_n1853_ & ~new_n1989_;
  assign new_n1991_ = \b[11]  & ~new_n1842_;
  assign new_n1992_ = ~new_n1836_ & new_n1991_;
  assign new_n1993_ = ~new_n1844_ & ~new_n1992_;
  assign new_n1994_ = ~new_n1990_ & new_n1993_;
  assign new_n1995_ = ~new_n1844_ & ~new_n1994_;
  assign new_n1996_ = \b[12]  & ~new_n1833_;
  assign new_n1997_ = ~new_n1827_ & new_n1996_;
  assign new_n1998_ = ~new_n1835_ & ~new_n1997_;
  assign new_n1999_ = ~new_n1995_ & new_n1998_;
  assign new_n2000_ = ~new_n1835_ & ~new_n1999_;
  assign new_n2001_ = \b[13]  & ~new_n1824_;
  assign new_n2002_ = ~new_n1818_ & new_n2001_;
  assign new_n2003_ = ~new_n1826_ & ~new_n2002_;
  assign new_n2004_ = ~new_n2000_ & new_n2003_;
  assign new_n2005_ = ~new_n1826_ & ~new_n2004_;
  assign new_n2006_ = ~new_n1642_ & ~\quotient[50] ;
  assign new_n2007_ = ~new_n1644_ & new_n1811_;
  assign new_n2008_ = ~new_n1807_ & new_n2007_;
  assign new_n2009_ = ~new_n1808_ & ~new_n1811_;
  assign new_n2010_ = ~new_n2008_ & ~new_n2009_;
  assign new_n2011_ = \quotient[50]  & ~new_n2010_;
  assign new_n2012_ = ~new_n2006_ & ~new_n2011_;
  assign new_n2013_ = ~\b[14]  & ~new_n2012_;
  assign new_n2014_ = \b[14]  & ~new_n2006_;
  assign new_n2015_ = ~new_n2011_ & new_n2014_;
  assign new_n2016_ = new_n369_ & new_n387_;
  assign new_n2017_ = new_n589_ & new_n2016_;
  assign new_n2018_ = new_n599_ & new_n2017_;
  assign new_n2019_ = ~new_n2015_ & new_n2018_;
  assign new_n2020_ = ~new_n2013_ & new_n2019_;
  assign new_n2021_ = ~new_n2005_ & new_n2020_;
  assign new_n2022_ = new_n1816_ & ~new_n2012_;
  assign \quotient[49]  = new_n2021_ | new_n2022_;
  assign new_n2024_ = ~new_n1835_ & new_n2003_;
  assign new_n2025_ = ~new_n1999_ & new_n2024_;
  assign new_n2026_ = ~new_n2000_ & ~new_n2003_;
  assign new_n2027_ = ~new_n2025_ & ~new_n2026_;
  assign new_n2028_ = \quotient[49]  & ~new_n2027_;
  assign new_n2029_ = ~new_n1825_ & ~new_n2022_;
  assign new_n2030_ = ~new_n2021_ & new_n2029_;
  assign new_n2031_ = ~new_n2028_ & ~new_n2030_;
  assign new_n2032_ = ~new_n1826_ & ~new_n2015_;
  assign new_n2033_ = ~new_n2013_ & new_n2032_;
  assign new_n2034_ = ~new_n2004_ & new_n2033_;
  assign new_n2035_ = ~new_n2013_ & ~new_n2015_;
  assign new_n2036_ = ~new_n2005_ & ~new_n2035_;
  assign new_n2037_ = ~new_n2034_ & ~new_n2036_;
  assign new_n2038_ = \quotient[49]  & ~new_n2037_;
  assign new_n2039_ = ~new_n2012_ & ~new_n2022_;
  assign new_n2040_ = ~new_n2021_ & new_n2039_;
  assign new_n2041_ = ~new_n2038_ & ~new_n2040_;
  assign new_n2042_ = ~\b[15]  & ~new_n2041_;
  assign new_n2043_ = ~\b[14]  & ~new_n2031_;
  assign new_n2044_ = ~new_n1844_ & new_n1998_;
  assign new_n2045_ = ~new_n1994_ & new_n2044_;
  assign new_n2046_ = ~new_n1995_ & ~new_n1998_;
  assign new_n2047_ = ~new_n2045_ & ~new_n2046_;
  assign new_n2048_ = \quotient[49]  & ~new_n2047_;
  assign new_n2049_ = ~new_n1834_ & ~new_n2022_;
  assign new_n2050_ = ~new_n2021_ & new_n2049_;
  assign new_n2051_ = ~new_n2048_ & ~new_n2050_;
  assign new_n2052_ = ~\b[13]  & ~new_n2051_;
  assign new_n2053_ = ~new_n1853_ & new_n1993_;
  assign new_n2054_ = ~new_n1989_ & new_n2053_;
  assign new_n2055_ = ~new_n1990_ & ~new_n1993_;
  assign new_n2056_ = ~new_n2054_ & ~new_n2055_;
  assign new_n2057_ = \quotient[49]  & ~new_n2056_;
  assign new_n2058_ = ~new_n1843_ & ~new_n2022_;
  assign new_n2059_ = ~new_n2021_ & new_n2058_;
  assign new_n2060_ = ~new_n2057_ & ~new_n2059_;
  assign new_n2061_ = ~\b[12]  & ~new_n2060_;
  assign new_n2062_ = ~new_n1862_ & new_n1988_;
  assign new_n2063_ = ~new_n1984_ & new_n2062_;
  assign new_n2064_ = ~new_n1985_ & ~new_n1988_;
  assign new_n2065_ = ~new_n2063_ & ~new_n2064_;
  assign new_n2066_ = \quotient[49]  & ~new_n2065_;
  assign new_n2067_ = ~new_n1852_ & ~new_n2022_;
  assign new_n2068_ = ~new_n2021_ & new_n2067_;
  assign new_n2069_ = ~new_n2066_ & ~new_n2068_;
  assign new_n2070_ = ~\b[11]  & ~new_n2069_;
  assign new_n2071_ = ~new_n1871_ & new_n1983_;
  assign new_n2072_ = ~new_n1979_ & new_n2071_;
  assign new_n2073_ = ~new_n1980_ & ~new_n1983_;
  assign new_n2074_ = ~new_n2072_ & ~new_n2073_;
  assign new_n2075_ = \quotient[49]  & ~new_n2074_;
  assign new_n2076_ = ~new_n1861_ & ~new_n2022_;
  assign new_n2077_ = ~new_n2021_ & new_n2076_;
  assign new_n2078_ = ~new_n2075_ & ~new_n2077_;
  assign new_n2079_ = ~\b[10]  & ~new_n2078_;
  assign new_n2080_ = ~new_n1880_ & new_n1978_;
  assign new_n2081_ = ~new_n1974_ & new_n2080_;
  assign new_n2082_ = ~new_n1975_ & ~new_n1978_;
  assign new_n2083_ = ~new_n2081_ & ~new_n2082_;
  assign new_n2084_ = \quotient[49]  & ~new_n2083_;
  assign new_n2085_ = ~new_n1870_ & ~new_n2022_;
  assign new_n2086_ = ~new_n2021_ & new_n2085_;
  assign new_n2087_ = ~new_n2084_ & ~new_n2086_;
  assign new_n2088_ = ~\b[9]  & ~new_n2087_;
  assign new_n2089_ = ~new_n1889_ & new_n1973_;
  assign new_n2090_ = ~new_n1969_ & new_n2089_;
  assign new_n2091_ = ~new_n1970_ & ~new_n1973_;
  assign new_n2092_ = ~new_n2090_ & ~new_n2091_;
  assign new_n2093_ = \quotient[49]  & ~new_n2092_;
  assign new_n2094_ = ~new_n1879_ & ~new_n2022_;
  assign new_n2095_ = ~new_n2021_ & new_n2094_;
  assign new_n2096_ = ~new_n2093_ & ~new_n2095_;
  assign new_n2097_ = ~\b[8]  & ~new_n2096_;
  assign new_n2098_ = ~new_n1898_ & new_n1968_;
  assign new_n2099_ = ~new_n1964_ & new_n2098_;
  assign new_n2100_ = ~new_n1965_ & ~new_n1968_;
  assign new_n2101_ = ~new_n2099_ & ~new_n2100_;
  assign new_n2102_ = \quotient[49]  & ~new_n2101_;
  assign new_n2103_ = ~new_n1888_ & ~new_n2022_;
  assign new_n2104_ = ~new_n2021_ & new_n2103_;
  assign new_n2105_ = ~new_n2102_ & ~new_n2104_;
  assign new_n2106_ = ~\b[7]  & ~new_n2105_;
  assign new_n2107_ = ~new_n1907_ & new_n1963_;
  assign new_n2108_ = ~new_n1959_ & new_n2107_;
  assign new_n2109_ = ~new_n1960_ & ~new_n1963_;
  assign new_n2110_ = ~new_n2108_ & ~new_n2109_;
  assign new_n2111_ = \quotient[49]  & ~new_n2110_;
  assign new_n2112_ = ~new_n1897_ & ~new_n2022_;
  assign new_n2113_ = ~new_n2021_ & new_n2112_;
  assign new_n2114_ = ~new_n2111_ & ~new_n2113_;
  assign new_n2115_ = ~\b[6]  & ~new_n2114_;
  assign new_n2116_ = ~new_n1916_ & new_n1958_;
  assign new_n2117_ = ~new_n1954_ & new_n2116_;
  assign new_n2118_ = ~new_n1955_ & ~new_n1958_;
  assign new_n2119_ = ~new_n2117_ & ~new_n2118_;
  assign new_n2120_ = \quotient[49]  & ~new_n2119_;
  assign new_n2121_ = ~new_n1906_ & ~new_n2022_;
  assign new_n2122_ = ~new_n2021_ & new_n2121_;
  assign new_n2123_ = ~new_n2120_ & ~new_n2122_;
  assign new_n2124_ = ~\b[5]  & ~new_n2123_;
  assign new_n2125_ = ~new_n1924_ & new_n1953_;
  assign new_n2126_ = ~new_n1949_ & new_n2125_;
  assign new_n2127_ = ~new_n1950_ & ~new_n1953_;
  assign new_n2128_ = ~new_n2126_ & ~new_n2127_;
  assign new_n2129_ = \quotient[49]  & ~new_n2128_;
  assign new_n2130_ = ~new_n1915_ & ~new_n2022_;
  assign new_n2131_ = ~new_n2021_ & new_n2130_;
  assign new_n2132_ = ~new_n2129_ & ~new_n2131_;
  assign new_n2133_ = ~\b[4]  & ~new_n2132_;
  assign new_n2134_ = ~new_n1944_ & new_n1948_;
  assign new_n2135_ = ~new_n1943_ & new_n2134_;
  assign new_n2136_ = ~new_n1945_ & ~new_n1948_;
  assign new_n2137_ = ~new_n2135_ & ~new_n2136_;
  assign new_n2138_ = \quotient[49]  & ~new_n2137_;
  assign new_n2139_ = ~new_n1923_ & ~new_n2022_;
  assign new_n2140_ = ~new_n2021_ & new_n2139_;
  assign new_n2141_ = ~new_n2138_ & ~new_n2140_;
  assign new_n2142_ = ~\b[3]  & ~new_n2141_;
  assign new_n2143_ = ~new_n1940_ & new_n1942_;
  assign new_n2144_ = ~new_n1938_ & new_n2143_;
  assign new_n2145_ = ~new_n1943_ & ~new_n2144_;
  assign new_n2146_ = \quotient[49]  & new_n2145_;
  assign new_n2147_ = ~new_n1937_ & ~new_n2022_;
  assign new_n2148_ = ~new_n2021_ & new_n2147_;
  assign new_n2149_ = ~new_n2146_ & ~new_n2148_;
  assign new_n2150_ = ~\b[2]  & ~new_n2149_;
  assign new_n2151_ = \b[0]  & \quotient[49] ;
  assign new_n2152_ = \a[49]  & ~new_n2151_;
  assign new_n2153_ = new_n1942_ & \quotient[49] ;
  assign new_n2154_ = ~new_n2152_ & ~new_n2153_;
  assign new_n2155_ = \b[1]  & ~new_n2154_;
  assign new_n2156_ = ~\b[1]  & ~new_n2153_;
  assign new_n2157_ = ~new_n2152_ & new_n2156_;
  assign new_n2158_ = ~new_n2155_ & ~new_n2157_;
  assign new_n2159_ = ~\a[48]  & \b[0] ;
  assign new_n2160_ = ~new_n2158_ & ~new_n2159_;
  assign new_n2161_ = ~\b[1]  & ~new_n2154_;
  assign new_n2162_ = ~new_n2160_ & ~new_n2161_;
  assign new_n2163_ = \b[2]  & ~new_n2148_;
  assign new_n2164_ = ~new_n2146_ & new_n2163_;
  assign new_n2165_ = ~new_n2150_ & ~new_n2164_;
  assign new_n2166_ = ~new_n2162_ & new_n2165_;
  assign new_n2167_ = ~new_n2150_ & ~new_n2166_;
  assign new_n2168_ = \b[3]  & ~new_n2140_;
  assign new_n2169_ = ~new_n2138_ & new_n2168_;
  assign new_n2170_ = ~new_n2142_ & ~new_n2169_;
  assign new_n2171_ = ~new_n2167_ & new_n2170_;
  assign new_n2172_ = ~new_n2142_ & ~new_n2171_;
  assign new_n2173_ = \b[4]  & ~new_n2131_;
  assign new_n2174_ = ~new_n2129_ & new_n2173_;
  assign new_n2175_ = ~new_n2133_ & ~new_n2174_;
  assign new_n2176_ = ~new_n2172_ & new_n2175_;
  assign new_n2177_ = ~new_n2133_ & ~new_n2176_;
  assign new_n2178_ = \b[5]  & ~new_n2122_;
  assign new_n2179_ = ~new_n2120_ & new_n2178_;
  assign new_n2180_ = ~new_n2124_ & ~new_n2179_;
  assign new_n2181_ = ~new_n2177_ & new_n2180_;
  assign new_n2182_ = ~new_n2124_ & ~new_n2181_;
  assign new_n2183_ = \b[6]  & ~new_n2113_;
  assign new_n2184_ = ~new_n2111_ & new_n2183_;
  assign new_n2185_ = ~new_n2115_ & ~new_n2184_;
  assign new_n2186_ = ~new_n2182_ & new_n2185_;
  assign new_n2187_ = ~new_n2115_ & ~new_n2186_;
  assign new_n2188_ = \b[7]  & ~new_n2104_;
  assign new_n2189_ = ~new_n2102_ & new_n2188_;
  assign new_n2190_ = ~new_n2106_ & ~new_n2189_;
  assign new_n2191_ = ~new_n2187_ & new_n2190_;
  assign new_n2192_ = ~new_n2106_ & ~new_n2191_;
  assign new_n2193_ = \b[8]  & ~new_n2095_;
  assign new_n2194_ = ~new_n2093_ & new_n2193_;
  assign new_n2195_ = ~new_n2097_ & ~new_n2194_;
  assign new_n2196_ = ~new_n2192_ & new_n2195_;
  assign new_n2197_ = ~new_n2097_ & ~new_n2196_;
  assign new_n2198_ = \b[9]  & ~new_n2086_;
  assign new_n2199_ = ~new_n2084_ & new_n2198_;
  assign new_n2200_ = ~new_n2088_ & ~new_n2199_;
  assign new_n2201_ = ~new_n2197_ & new_n2200_;
  assign new_n2202_ = ~new_n2088_ & ~new_n2201_;
  assign new_n2203_ = \b[10]  & ~new_n2077_;
  assign new_n2204_ = ~new_n2075_ & new_n2203_;
  assign new_n2205_ = ~new_n2079_ & ~new_n2204_;
  assign new_n2206_ = ~new_n2202_ & new_n2205_;
  assign new_n2207_ = ~new_n2079_ & ~new_n2206_;
  assign new_n2208_ = \b[11]  & ~new_n2068_;
  assign new_n2209_ = ~new_n2066_ & new_n2208_;
  assign new_n2210_ = ~new_n2070_ & ~new_n2209_;
  assign new_n2211_ = ~new_n2207_ & new_n2210_;
  assign new_n2212_ = ~new_n2070_ & ~new_n2211_;
  assign new_n2213_ = \b[12]  & ~new_n2059_;
  assign new_n2214_ = ~new_n2057_ & new_n2213_;
  assign new_n2215_ = ~new_n2061_ & ~new_n2214_;
  assign new_n2216_ = ~new_n2212_ & new_n2215_;
  assign new_n2217_ = ~new_n2061_ & ~new_n2216_;
  assign new_n2218_ = \b[13]  & ~new_n2050_;
  assign new_n2219_ = ~new_n2048_ & new_n2218_;
  assign new_n2220_ = ~new_n2052_ & ~new_n2219_;
  assign new_n2221_ = ~new_n2217_ & new_n2220_;
  assign new_n2222_ = ~new_n2052_ & ~new_n2221_;
  assign new_n2223_ = \b[14]  & ~new_n2030_;
  assign new_n2224_ = ~new_n2028_ & new_n2223_;
  assign new_n2225_ = ~new_n2043_ & ~new_n2224_;
  assign new_n2226_ = ~new_n2222_ & new_n2225_;
  assign new_n2227_ = ~new_n2043_ & ~new_n2226_;
  assign new_n2228_ = \b[15]  & ~new_n2040_;
  assign new_n2229_ = ~new_n2038_ & new_n2228_;
  assign new_n2230_ = ~new_n2042_ & ~new_n2229_;
  assign new_n2231_ = ~new_n2227_ & new_n2230_;
  assign new_n2232_ = ~new_n2042_ & ~new_n2231_;
  assign \quotient[48]  = new_n346_ & ~new_n2232_;
  assign new_n2234_ = ~new_n2031_ & ~\quotient[48] ;
  assign new_n2235_ = ~new_n2052_ & new_n2225_;
  assign new_n2236_ = ~new_n2221_ & new_n2235_;
  assign new_n2237_ = ~new_n2222_ & ~new_n2225_;
  assign new_n2238_ = ~new_n2236_ & ~new_n2237_;
  assign new_n2239_ = new_n346_ & ~new_n2238_;
  assign new_n2240_ = ~new_n2232_ & new_n2239_;
  assign new_n2241_ = ~new_n2234_ & ~new_n2240_;
  assign new_n2242_ = ~new_n2041_ & ~\quotient[48] ;
  assign new_n2243_ = ~new_n2043_ & new_n2230_;
  assign new_n2244_ = ~new_n2226_ & new_n2243_;
  assign new_n2245_ = ~new_n2227_ & ~new_n2230_;
  assign new_n2246_ = ~new_n2244_ & ~new_n2245_;
  assign new_n2247_ = \quotient[48]  & ~new_n2246_;
  assign new_n2248_ = ~new_n2242_ & ~new_n2247_;
  assign new_n2249_ = ~\b[16]  & ~new_n2248_;
  assign new_n2250_ = ~\b[15]  & ~new_n2241_;
  assign new_n2251_ = ~new_n2051_ & ~\quotient[48] ;
  assign new_n2252_ = ~new_n2061_ & new_n2220_;
  assign new_n2253_ = ~new_n2216_ & new_n2252_;
  assign new_n2254_ = ~new_n2217_ & ~new_n2220_;
  assign new_n2255_ = ~new_n2253_ & ~new_n2254_;
  assign new_n2256_ = new_n346_ & ~new_n2255_;
  assign new_n2257_ = ~new_n2232_ & new_n2256_;
  assign new_n2258_ = ~new_n2251_ & ~new_n2257_;
  assign new_n2259_ = ~\b[14]  & ~new_n2258_;
  assign new_n2260_ = ~new_n2060_ & ~\quotient[48] ;
  assign new_n2261_ = ~new_n2070_ & new_n2215_;
  assign new_n2262_ = ~new_n2211_ & new_n2261_;
  assign new_n2263_ = ~new_n2212_ & ~new_n2215_;
  assign new_n2264_ = ~new_n2262_ & ~new_n2263_;
  assign new_n2265_ = new_n346_ & ~new_n2264_;
  assign new_n2266_ = ~new_n2232_ & new_n2265_;
  assign new_n2267_ = ~new_n2260_ & ~new_n2266_;
  assign new_n2268_ = ~\b[13]  & ~new_n2267_;
  assign new_n2269_ = ~new_n2069_ & ~\quotient[48] ;
  assign new_n2270_ = ~new_n2079_ & new_n2210_;
  assign new_n2271_ = ~new_n2206_ & new_n2270_;
  assign new_n2272_ = ~new_n2207_ & ~new_n2210_;
  assign new_n2273_ = ~new_n2271_ & ~new_n2272_;
  assign new_n2274_ = new_n346_ & ~new_n2273_;
  assign new_n2275_ = ~new_n2232_ & new_n2274_;
  assign new_n2276_ = ~new_n2269_ & ~new_n2275_;
  assign new_n2277_ = ~\b[12]  & ~new_n2276_;
  assign new_n2278_ = ~new_n2078_ & ~\quotient[48] ;
  assign new_n2279_ = ~new_n2088_ & new_n2205_;
  assign new_n2280_ = ~new_n2201_ & new_n2279_;
  assign new_n2281_ = ~new_n2202_ & ~new_n2205_;
  assign new_n2282_ = ~new_n2280_ & ~new_n2281_;
  assign new_n2283_ = new_n346_ & ~new_n2282_;
  assign new_n2284_ = ~new_n2232_ & new_n2283_;
  assign new_n2285_ = ~new_n2278_ & ~new_n2284_;
  assign new_n2286_ = ~\b[11]  & ~new_n2285_;
  assign new_n2287_ = ~new_n2087_ & ~\quotient[48] ;
  assign new_n2288_ = ~new_n2097_ & new_n2200_;
  assign new_n2289_ = ~new_n2196_ & new_n2288_;
  assign new_n2290_ = ~new_n2197_ & ~new_n2200_;
  assign new_n2291_ = ~new_n2289_ & ~new_n2290_;
  assign new_n2292_ = new_n346_ & ~new_n2291_;
  assign new_n2293_ = ~new_n2232_ & new_n2292_;
  assign new_n2294_ = ~new_n2287_ & ~new_n2293_;
  assign new_n2295_ = ~\b[10]  & ~new_n2294_;
  assign new_n2296_ = ~new_n2096_ & ~\quotient[48] ;
  assign new_n2297_ = ~new_n2106_ & new_n2195_;
  assign new_n2298_ = ~new_n2191_ & new_n2297_;
  assign new_n2299_ = ~new_n2192_ & ~new_n2195_;
  assign new_n2300_ = ~new_n2298_ & ~new_n2299_;
  assign new_n2301_ = new_n346_ & ~new_n2300_;
  assign new_n2302_ = ~new_n2232_ & new_n2301_;
  assign new_n2303_ = ~new_n2296_ & ~new_n2302_;
  assign new_n2304_ = ~\b[9]  & ~new_n2303_;
  assign new_n2305_ = ~new_n2105_ & ~\quotient[48] ;
  assign new_n2306_ = ~new_n2115_ & new_n2190_;
  assign new_n2307_ = ~new_n2186_ & new_n2306_;
  assign new_n2308_ = ~new_n2187_ & ~new_n2190_;
  assign new_n2309_ = ~new_n2307_ & ~new_n2308_;
  assign new_n2310_ = new_n346_ & ~new_n2309_;
  assign new_n2311_ = ~new_n2232_ & new_n2310_;
  assign new_n2312_ = ~new_n2305_ & ~new_n2311_;
  assign new_n2313_ = ~\b[8]  & ~new_n2312_;
  assign new_n2314_ = ~new_n2114_ & ~\quotient[48] ;
  assign new_n2315_ = ~new_n2124_ & new_n2185_;
  assign new_n2316_ = ~new_n2181_ & new_n2315_;
  assign new_n2317_ = ~new_n2182_ & ~new_n2185_;
  assign new_n2318_ = ~new_n2316_ & ~new_n2317_;
  assign new_n2319_ = new_n346_ & ~new_n2318_;
  assign new_n2320_ = ~new_n2232_ & new_n2319_;
  assign new_n2321_ = ~new_n2314_ & ~new_n2320_;
  assign new_n2322_ = ~\b[7]  & ~new_n2321_;
  assign new_n2323_ = ~new_n2123_ & ~\quotient[48] ;
  assign new_n2324_ = ~new_n2133_ & new_n2180_;
  assign new_n2325_ = ~new_n2176_ & new_n2324_;
  assign new_n2326_ = ~new_n2177_ & ~new_n2180_;
  assign new_n2327_ = ~new_n2325_ & ~new_n2326_;
  assign new_n2328_ = new_n346_ & ~new_n2327_;
  assign new_n2329_ = ~new_n2232_ & new_n2328_;
  assign new_n2330_ = ~new_n2323_ & ~new_n2329_;
  assign new_n2331_ = ~\b[6]  & ~new_n2330_;
  assign new_n2332_ = ~new_n2132_ & ~\quotient[48] ;
  assign new_n2333_ = ~new_n2142_ & new_n2175_;
  assign new_n2334_ = ~new_n2171_ & new_n2333_;
  assign new_n2335_ = ~new_n2172_ & ~new_n2175_;
  assign new_n2336_ = ~new_n2334_ & ~new_n2335_;
  assign new_n2337_ = new_n346_ & ~new_n2336_;
  assign new_n2338_ = ~new_n2232_ & new_n2337_;
  assign new_n2339_ = ~new_n2332_ & ~new_n2338_;
  assign new_n2340_ = ~\b[5]  & ~new_n2339_;
  assign new_n2341_ = ~new_n2141_ & ~\quotient[48] ;
  assign new_n2342_ = ~new_n2150_ & new_n2170_;
  assign new_n2343_ = ~new_n2166_ & new_n2342_;
  assign new_n2344_ = ~new_n2167_ & ~new_n2170_;
  assign new_n2345_ = ~new_n2343_ & ~new_n2344_;
  assign new_n2346_ = new_n346_ & ~new_n2345_;
  assign new_n2347_ = ~new_n2232_ & new_n2346_;
  assign new_n2348_ = ~new_n2341_ & ~new_n2347_;
  assign new_n2349_ = ~\b[4]  & ~new_n2348_;
  assign new_n2350_ = ~new_n2149_ & ~\quotient[48] ;
  assign new_n2351_ = ~new_n2161_ & new_n2165_;
  assign new_n2352_ = ~new_n2160_ & new_n2351_;
  assign new_n2353_ = ~new_n2162_ & ~new_n2165_;
  assign new_n2354_ = ~new_n2352_ & ~new_n2353_;
  assign new_n2355_ = new_n346_ & ~new_n2354_;
  assign new_n2356_ = ~new_n2232_ & new_n2355_;
  assign new_n2357_ = ~new_n2350_ & ~new_n2356_;
  assign new_n2358_ = ~\b[3]  & ~new_n2357_;
  assign new_n2359_ = ~new_n2154_ & ~\quotient[48] ;
  assign new_n2360_ = ~new_n2157_ & new_n2159_;
  assign new_n2361_ = ~new_n2155_ & new_n2360_;
  assign new_n2362_ = new_n346_ & ~new_n2361_;
  assign new_n2363_ = ~new_n2160_ & new_n2362_;
  assign new_n2364_ = ~new_n2232_ & new_n2363_;
  assign new_n2365_ = ~new_n2359_ & ~new_n2364_;
  assign new_n2366_ = ~\b[2]  & ~new_n2365_;
  assign new_n2367_ = \b[0]  & ~\b[16] ;
  assign new_n2368_ = new_n369_ & new_n2367_;
  assign new_n2369_ = new_n589_ & new_n2368_;
  assign new_n2370_ = new_n599_ & new_n2369_;
  assign new_n2371_ = ~new_n2232_ & new_n2370_;
  assign new_n2372_ = \a[48]  & ~new_n2371_;
  assign new_n2373_ = new_n271_ & new_n2159_;
  assign new_n2374_ = new_n318_ & new_n2373_;
  assign new_n2375_ = new_n512_ & new_n2374_;
  assign new_n2376_ = ~new_n2232_ & new_n2375_;
  assign new_n2377_ = ~new_n2372_ & ~new_n2376_;
  assign new_n2378_ = \b[1]  & ~new_n2377_;
  assign new_n2379_ = ~\b[1]  & ~new_n2376_;
  assign new_n2380_ = ~new_n2372_ & new_n2379_;
  assign new_n2381_ = ~new_n2378_ & ~new_n2380_;
  assign new_n2382_ = ~\a[47]  & \b[0] ;
  assign new_n2383_ = ~new_n2381_ & ~new_n2382_;
  assign new_n2384_ = ~\b[1]  & ~new_n2377_;
  assign new_n2385_ = ~new_n2383_ & ~new_n2384_;
  assign new_n2386_ = \b[2]  & ~new_n2364_;
  assign new_n2387_ = ~new_n2359_ & new_n2386_;
  assign new_n2388_ = ~new_n2366_ & ~new_n2387_;
  assign new_n2389_ = ~new_n2385_ & new_n2388_;
  assign new_n2390_ = ~new_n2366_ & ~new_n2389_;
  assign new_n2391_ = \b[3]  & ~new_n2356_;
  assign new_n2392_ = ~new_n2350_ & new_n2391_;
  assign new_n2393_ = ~new_n2358_ & ~new_n2392_;
  assign new_n2394_ = ~new_n2390_ & new_n2393_;
  assign new_n2395_ = ~new_n2358_ & ~new_n2394_;
  assign new_n2396_ = \b[4]  & ~new_n2347_;
  assign new_n2397_ = ~new_n2341_ & new_n2396_;
  assign new_n2398_ = ~new_n2349_ & ~new_n2397_;
  assign new_n2399_ = ~new_n2395_ & new_n2398_;
  assign new_n2400_ = ~new_n2349_ & ~new_n2399_;
  assign new_n2401_ = \b[5]  & ~new_n2338_;
  assign new_n2402_ = ~new_n2332_ & new_n2401_;
  assign new_n2403_ = ~new_n2340_ & ~new_n2402_;
  assign new_n2404_ = ~new_n2400_ & new_n2403_;
  assign new_n2405_ = ~new_n2340_ & ~new_n2404_;
  assign new_n2406_ = \b[6]  & ~new_n2329_;
  assign new_n2407_ = ~new_n2323_ & new_n2406_;
  assign new_n2408_ = ~new_n2331_ & ~new_n2407_;
  assign new_n2409_ = ~new_n2405_ & new_n2408_;
  assign new_n2410_ = ~new_n2331_ & ~new_n2409_;
  assign new_n2411_ = \b[7]  & ~new_n2320_;
  assign new_n2412_ = ~new_n2314_ & new_n2411_;
  assign new_n2413_ = ~new_n2322_ & ~new_n2412_;
  assign new_n2414_ = ~new_n2410_ & new_n2413_;
  assign new_n2415_ = ~new_n2322_ & ~new_n2414_;
  assign new_n2416_ = \b[8]  & ~new_n2311_;
  assign new_n2417_ = ~new_n2305_ & new_n2416_;
  assign new_n2418_ = ~new_n2313_ & ~new_n2417_;
  assign new_n2419_ = ~new_n2415_ & new_n2418_;
  assign new_n2420_ = ~new_n2313_ & ~new_n2419_;
  assign new_n2421_ = \b[9]  & ~new_n2302_;
  assign new_n2422_ = ~new_n2296_ & new_n2421_;
  assign new_n2423_ = ~new_n2304_ & ~new_n2422_;
  assign new_n2424_ = ~new_n2420_ & new_n2423_;
  assign new_n2425_ = ~new_n2304_ & ~new_n2424_;
  assign new_n2426_ = \b[10]  & ~new_n2293_;
  assign new_n2427_ = ~new_n2287_ & new_n2426_;
  assign new_n2428_ = ~new_n2295_ & ~new_n2427_;
  assign new_n2429_ = ~new_n2425_ & new_n2428_;
  assign new_n2430_ = ~new_n2295_ & ~new_n2429_;
  assign new_n2431_ = \b[11]  & ~new_n2284_;
  assign new_n2432_ = ~new_n2278_ & new_n2431_;
  assign new_n2433_ = ~new_n2286_ & ~new_n2432_;
  assign new_n2434_ = ~new_n2430_ & new_n2433_;
  assign new_n2435_ = ~new_n2286_ & ~new_n2434_;
  assign new_n2436_ = \b[12]  & ~new_n2275_;
  assign new_n2437_ = ~new_n2269_ & new_n2436_;
  assign new_n2438_ = ~new_n2277_ & ~new_n2437_;
  assign new_n2439_ = ~new_n2435_ & new_n2438_;
  assign new_n2440_ = ~new_n2277_ & ~new_n2439_;
  assign new_n2441_ = \b[13]  & ~new_n2266_;
  assign new_n2442_ = ~new_n2260_ & new_n2441_;
  assign new_n2443_ = ~new_n2268_ & ~new_n2442_;
  assign new_n2444_ = ~new_n2440_ & new_n2443_;
  assign new_n2445_ = ~new_n2268_ & ~new_n2444_;
  assign new_n2446_ = \b[14]  & ~new_n2257_;
  assign new_n2447_ = ~new_n2251_ & new_n2446_;
  assign new_n2448_ = ~new_n2259_ & ~new_n2447_;
  assign new_n2449_ = ~new_n2445_ & new_n2448_;
  assign new_n2450_ = ~new_n2259_ & ~new_n2449_;
  assign new_n2451_ = \b[15]  & ~new_n2240_;
  assign new_n2452_ = ~new_n2234_ & new_n2451_;
  assign new_n2453_ = ~new_n2250_ & ~new_n2452_;
  assign new_n2454_ = ~new_n2450_ & new_n2453_;
  assign new_n2455_ = ~new_n2250_ & ~new_n2454_;
  assign new_n2456_ = \b[16]  & ~new_n2242_;
  assign new_n2457_ = ~new_n2247_ & new_n2456_;
  assign new_n2458_ = ~new_n2249_ & ~new_n2457_;
  assign new_n2459_ = ~new_n2455_ & new_n2458_;
  assign new_n2460_ = ~new_n2249_ & ~new_n2459_;
  assign \quotient[47]  = new_n475_ & ~new_n2460_;
  assign new_n2462_ = ~new_n2241_ & ~\quotient[47] ;
  assign new_n2463_ = ~new_n2259_ & new_n2453_;
  assign new_n2464_ = ~new_n2449_ & new_n2463_;
  assign new_n2465_ = ~new_n2450_ & ~new_n2453_;
  assign new_n2466_ = ~new_n2464_ & ~new_n2465_;
  assign new_n2467_ = new_n475_ & ~new_n2466_;
  assign new_n2468_ = ~new_n2460_ & new_n2467_;
  assign new_n2469_ = ~new_n2462_ & ~new_n2468_;
  assign new_n2470_ = ~\b[16]  & ~new_n2469_;
  assign new_n2471_ = ~new_n2258_ & ~\quotient[47] ;
  assign new_n2472_ = ~new_n2268_ & new_n2448_;
  assign new_n2473_ = ~new_n2444_ & new_n2472_;
  assign new_n2474_ = ~new_n2445_ & ~new_n2448_;
  assign new_n2475_ = ~new_n2473_ & ~new_n2474_;
  assign new_n2476_ = new_n475_ & ~new_n2475_;
  assign new_n2477_ = ~new_n2460_ & new_n2476_;
  assign new_n2478_ = ~new_n2471_ & ~new_n2477_;
  assign new_n2479_ = ~\b[15]  & ~new_n2478_;
  assign new_n2480_ = ~new_n2267_ & ~\quotient[47] ;
  assign new_n2481_ = ~new_n2277_ & new_n2443_;
  assign new_n2482_ = ~new_n2439_ & new_n2481_;
  assign new_n2483_ = ~new_n2440_ & ~new_n2443_;
  assign new_n2484_ = ~new_n2482_ & ~new_n2483_;
  assign new_n2485_ = new_n475_ & ~new_n2484_;
  assign new_n2486_ = ~new_n2460_ & new_n2485_;
  assign new_n2487_ = ~new_n2480_ & ~new_n2486_;
  assign new_n2488_ = ~\b[14]  & ~new_n2487_;
  assign new_n2489_ = ~new_n2276_ & ~\quotient[47] ;
  assign new_n2490_ = ~new_n2286_ & new_n2438_;
  assign new_n2491_ = ~new_n2434_ & new_n2490_;
  assign new_n2492_ = ~new_n2435_ & ~new_n2438_;
  assign new_n2493_ = ~new_n2491_ & ~new_n2492_;
  assign new_n2494_ = new_n475_ & ~new_n2493_;
  assign new_n2495_ = ~new_n2460_ & new_n2494_;
  assign new_n2496_ = ~new_n2489_ & ~new_n2495_;
  assign new_n2497_ = ~\b[13]  & ~new_n2496_;
  assign new_n2498_ = ~new_n2285_ & ~\quotient[47] ;
  assign new_n2499_ = ~new_n2295_ & new_n2433_;
  assign new_n2500_ = ~new_n2429_ & new_n2499_;
  assign new_n2501_ = ~new_n2430_ & ~new_n2433_;
  assign new_n2502_ = ~new_n2500_ & ~new_n2501_;
  assign new_n2503_ = new_n475_ & ~new_n2502_;
  assign new_n2504_ = ~new_n2460_ & new_n2503_;
  assign new_n2505_ = ~new_n2498_ & ~new_n2504_;
  assign new_n2506_ = ~\b[12]  & ~new_n2505_;
  assign new_n2507_ = ~new_n2294_ & ~\quotient[47] ;
  assign new_n2508_ = ~new_n2304_ & new_n2428_;
  assign new_n2509_ = ~new_n2424_ & new_n2508_;
  assign new_n2510_ = ~new_n2425_ & ~new_n2428_;
  assign new_n2511_ = ~new_n2509_ & ~new_n2510_;
  assign new_n2512_ = new_n475_ & ~new_n2511_;
  assign new_n2513_ = ~new_n2460_ & new_n2512_;
  assign new_n2514_ = ~new_n2507_ & ~new_n2513_;
  assign new_n2515_ = ~\b[11]  & ~new_n2514_;
  assign new_n2516_ = ~new_n2303_ & ~\quotient[47] ;
  assign new_n2517_ = ~new_n2313_ & new_n2423_;
  assign new_n2518_ = ~new_n2419_ & new_n2517_;
  assign new_n2519_ = ~new_n2420_ & ~new_n2423_;
  assign new_n2520_ = ~new_n2518_ & ~new_n2519_;
  assign new_n2521_ = new_n475_ & ~new_n2520_;
  assign new_n2522_ = ~new_n2460_ & new_n2521_;
  assign new_n2523_ = ~new_n2516_ & ~new_n2522_;
  assign new_n2524_ = ~\b[10]  & ~new_n2523_;
  assign new_n2525_ = ~new_n2312_ & ~\quotient[47] ;
  assign new_n2526_ = ~new_n2322_ & new_n2418_;
  assign new_n2527_ = ~new_n2414_ & new_n2526_;
  assign new_n2528_ = ~new_n2415_ & ~new_n2418_;
  assign new_n2529_ = ~new_n2527_ & ~new_n2528_;
  assign new_n2530_ = new_n475_ & ~new_n2529_;
  assign new_n2531_ = ~new_n2460_ & new_n2530_;
  assign new_n2532_ = ~new_n2525_ & ~new_n2531_;
  assign new_n2533_ = ~\b[9]  & ~new_n2532_;
  assign new_n2534_ = ~new_n2321_ & ~\quotient[47] ;
  assign new_n2535_ = ~new_n2331_ & new_n2413_;
  assign new_n2536_ = ~new_n2409_ & new_n2535_;
  assign new_n2537_ = ~new_n2410_ & ~new_n2413_;
  assign new_n2538_ = ~new_n2536_ & ~new_n2537_;
  assign new_n2539_ = new_n475_ & ~new_n2538_;
  assign new_n2540_ = ~new_n2460_ & new_n2539_;
  assign new_n2541_ = ~new_n2534_ & ~new_n2540_;
  assign new_n2542_ = ~\b[8]  & ~new_n2541_;
  assign new_n2543_ = ~new_n2330_ & ~\quotient[47] ;
  assign new_n2544_ = ~new_n2340_ & new_n2408_;
  assign new_n2545_ = ~new_n2404_ & new_n2544_;
  assign new_n2546_ = ~new_n2405_ & ~new_n2408_;
  assign new_n2547_ = ~new_n2545_ & ~new_n2546_;
  assign new_n2548_ = new_n475_ & ~new_n2547_;
  assign new_n2549_ = ~new_n2460_ & new_n2548_;
  assign new_n2550_ = ~new_n2543_ & ~new_n2549_;
  assign new_n2551_ = ~\b[7]  & ~new_n2550_;
  assign new_n2552_ = ~new_n2339_ & ~\quotient[47] ;
  assign new_n2553_ = ~new_n2349_ & new_n2403_;
  assign new_n2554_ = ~new_n2399_ & new_n2553_;
  assign new_n2555_ = ~new_n2400_ & ~new_n2403_;
  assign new_n2556_ = ~new_n2554_ & ~new_n2555_;
  assign new_n2557_ = new_n475_ & ~new_n2556_;
  assign new_n2558_ = ~new_n2460_ & new_n2557_;
  assign new_n2559_ = ~new_n2552_ & ~new_n2558_;
  assign new_n2560_ = ~\b[6]  & ~new_n2559_;
  assign new_n2561_ = ~new_n2348_ & ~\quotient[47] ;
  assign new_n2562_ = ~new_n2358_ & new_n2398_;
  assign new_n2563_ = ~new_n2394_ & new_n2562_;
  assign new_n2564_ = ~new_n2395_ & ~new_n2398_;
  assign new_n2565_ = ~new_n2563_ & ~new_n2564_;
  assign new_n2566_ = new_n475_ & ~new_n2565_;
  assign new_n2567_ = ~new_n2460_ & new_n2566_;
  assign new_n2568_ = ~new_n2561_ & ~new_n2567_;
  assign new_n2569_ = ~\b[5]  & ~new_n2568_;
  assign new_n2570_ = ~new_n2357_ & ~\quotient[47] ;
  assign new_n2571_ = ~new_n2366_ & new_n2393_;
  assign new_n2572_ = ~new_n2389_ & new_n2571_;
  assign new_n2573_ = ~new_n2390_ & ~new_n2393_;
  assign new_n2574_ = ~new_n2572_ & ~new_n2573_;
  assign new_n2575_ = new_n475_ & ~new_n2574_;
  assign new_n2576_ = ~new_n2460_ & new_n2575_;
  assign new_n2577_ = ~new_n2570_ & ~new_n2576_;
  assign new_n2578_ = ~\b[4]  & ~new_n2577_;
  assign new_n2579_ = ~new_n2365_ & ~\quotient[47] ;
  assign new_n2580_ = ~new_n2384_ & new_n2388_;
  assign new_n2581_ = ~new_n2383_ & new_n2580_;
  assign new_n2582_ = ~new_n2385_ & ~new_n2388_;
  assign new_n2583_ = ~new_n2581_ & ~new_n2582_;
  assign new_n2584_ = new_n475_ & ~new_n2583_;
  assign new_n2585_ = ~new_n2460_ & new_n2584_;
  assign new_n2586_ = ~new_n2579_ & ~new_n2585_;
  assign new_n2587_ = ~\b[3]  & ~new_n2586_;
  assign new_n2588_ = ~new_n2377_ & ~\quotient[47] ;
  assign new_n2589_ = ~new_n2380_ & new_n2382_;
  assign new_n2590_ = ~new_n2378_ & new_n2589_;
  assign new_n2591_ = new_n475_ & ~new_n2590_;
  assign new_n2592_ = ~new_n2383_ & new_n2591_;
  assign new_n2593_ = ~new_n2460_ & new_n2592_;
  assign new_n2594_ = ~new_n2588_ & ~new_n2593_;
  assign new_n2595_ = ~\b[2]  & ~new_n2594_;
  assign new_n2596_ = \b[0]  & ~\b[17] ;
  assign new_n2597_ = new_n270_ & new_n2596_;
  assign new_n2598_ = new_n309_ & new_n2597_;
  assign new_n2599_ = new_n343_ & new_n2598_;
  assign new_n2600_ = new_n341_ & new_n2599_;
  assign new_n2601_ = new_n338_ & new_n2600_;
  assign new_n2602_ = ~new_n2460_ & new_n2601_;
  assign new_n2603_ = \a[47]  & ~new_n2602_;
  assign new_n2604_ = new_n369_ & new_n2382_;
  assign new_n2605_ = new_n589_ & new_n2604_;
  assign new_n2606_ = new_n599_ & new_n2605_;
  assign new_n2607_ = ~new_n2460_ & new_n2606_;
  assign new_n2608_ = ~new_n2603_ & ~new_n2607_;
  assign new_n2609_ = \b[1]  & ~new_n2608_;
  assign new_n2610_ = ~\b[1]  & ~new_n2607_;
  assign new_n2611_ = ~new_n2603_ & new_n2610_;
  assign new_n2612_ = ~new_n2609_ & ~new_n2611_;
  assign new_n2613_ = ~\a[46]  & \b[0] ;
  assign new_n2614_ = ~new_n2612_ & ~new_n2613_;
  assign new_n2615_ = ~\b[1]  & ~new_n2608_;
  assign new_n2616_ = ~new_n2614_ & ~new_n2615_;
  assign new_n2617_ = \b[2]  & ~new_n2593_;
  assign new_n2618_ = ~new_n2588_ & new_n2617_;
  assign new_n2619_ = ~new_n2595_ & ~new_n2618_;
  assign new_n2620_ = ~new_n2616_ & new_n2619_;
  assign new_n2621_ = ~new_n2595_ & ~new_n2620_;
  assign new_n2622_ = \b[3]  & ~new_n2585_;
  assign new_n2623_ = ~new_n2579_ & new_n2622_;
  assign new_n2624_ = ~new_n2587_ & ~new_n2623_;
  assign new_n2625_ = ~new_n2621_ & new_n2624_;
  assign new_n2626_ = ~new_n2587_ & ~new_n2625_;
  assign new_n2627_ = \b[4]  & ~new_n2576_;
  assign new_n2628_ = ~new_n2570_ & new_n2627_;
  assign new_n2629_ = ~new_n2578_ & ~new_n2628_;
  assign new_n2630_ = ~new_n2626_ & new_n2629_;
  assign new_n2631_ = ~new_n2578_ & ~new_n2630_;
  assign new_n2632_ = \b[5]  & ~new_n2567_;
  assign new_n2633_ = ~new_n2561_ & new_n2632_;
  assign new_n2634_ = ~new_n2569_ & ~new_n2633_;
  assign new_n2635_ = ~new_n2631_ & new_n2634_;
  assign new_n2636_ = ~new_n2569_ & ~new_n2635_;
  assign new_n2637_ = \b[6]  & ~new_n2558_;
  assign new_n2638_ = ~new_n2552_ & new_n2637_;
  assign new_n2639_ = ~new_n2560_ & ~new_n2638_;
  assign new_n2640_ = ~new_n2636_ & new_n2639_;
  assign new_n2641_ = ~new_n2560_ & ~new_n2640_;
  assign new_n2642_ = \b[7]  & ~new_n2549_;
  assign new_n2643_ = ~new_n2543_ & new_n2642_;
  assign new_n2644_ = ~new_n2551_ & ~new_n2643_;
  assign new_n2645_ = ~new_n2641_ & new_n2644_;
  assign new_n2646_ = ~new_n2551_ & ~new_n2645_;
  assign new_n2647_ = \b[8]  & ~new_n2540_;
  assign new_n2648_ = ~new_n2534_ & new_n2647_;
  assign new_n2649_ = ~new_n2542_ & ~new_n2648_;
  assign new_n2650_ = ~new_n2646_ & new_n2649_;
  assign new_n2651_ = ~new_n2542_ & ~new_n2650_;
  assign new_n2652_ = \b[9]  & ~new_n2531_;
  assign new_n2653_ = ~new_n2525_ & new_n2652_;
  assign new_n2654_ = ~new_n2533_ & ~new_n2653_;
  assign new_n2655_ = ~new_n2651_ & new_n2654_;
  assign new_n2656_ = ~new_n2533_ & ~new_n2655_;
  assign new_n2657_ = \b[10]  & ~new_n2522_;
  assign new_n2658_ = ~new_n2516_ & new_n2657_;
  assign new_n2659_ = ~new_n2524_ & ~new_n2658_;
  assign new_n2660_ = ~new_n2656_ & new_n2659_;
  assign new_n2661_ = ~new_n2524_ & ~new_n2660_;
  assign new_n2662_ = \b[11]  & ~new_n2513_;
  assign new_n2663_ = ~new_n2507_ & new_n2662_;
  assign new_n2664_ = ~new_n2515_ & ~new_n2663_;
  assign new_n2665_ = ~new_n2661_ & new_n2664_;
  assign new_n2666_ = ~new_n2515_ & ~new_n2665_;
  assign new_n2667_ = \b[12]  & ~new_n2504_;
  assign new_n2668_ = ~new_n2498_ & new_n2667_;
  assign new_n2669_ = ~new_n2506_ & ~new_n2668_;
  assign new_n2670_ = ~new_n2666_ & new_n2669_;
  assign new_n2671_ = ~new_n2506_ & ~new_n2670_;
  assign new_n2672_ = \b[13]  & ~new_n2495_;
  assign new_n2673_ = ~new_n2489_ & new_n2672_;
  assign new_n2674_ = ~new_n2497_ & ~new_n2673_;
  assign new_n2675_ = ~new_n2671_ & new_n2674_;
  assign new_n2676_ = ~new_n2497_ & ~new_n2675_;
  assign new_n2677_ = \b[14]  & ~new_n2486_;
  assign new_n2678_ = ~new_n2480_ & new_n2677_;
  assign new_n2679_ = ~new_n2488_ & ~new_n2678_;
  assign new_n2680_ = ~new_n2676_ & new_n2679_;
  assign new_n2681_ = ~new_n2488_ & ~new_n2680_;
  assign new_n2682_ = \b[15]  & ~new_n2477_;
  assign new_n2683_ = ~new_n2471_ & new_n2682_;
  assign new_n2684_ = ~new_n2479_ & ~new_n2683_;
  assign new_n2685_ = ~new_n2681_ & new_n2684_;
  assign new_n2686_ = ~new_n2479_ & ~new_n2685_;
  assign new_n2687_ = \b[16]  & ~new_n2468_;
  assign new_n2688_ = ~new_n2462_ & new_n2687_;
  assign new_n2689_ = ~new_n2470_ & ~new_n2688_;
  assign new_n2690_ = ~new_n2686_ & new_n2689_;
  assign new_n2691_ = ~new_n2470_ & ~new_n2690_;
  assign new_n2692_ = ~new_n2248_ & ~\quotient[47] ;
  assign new_n2693_ = ~new_n2250_ & new_n2458_;
  assign new_n2694_ = ~new_n2454_ & new_n2693_;
  assign new_n2695_ = ~new_n2455_ & ~new_n2458_;
  assign new_n2696_ = ~new_n2694_ & ~new_n2695_;
  assign new_n2697_ = \quotient[47]  & ~new_n2696_;
  assign new_n2698_ = ~new_n2692_ & ~new_n2697_;
  assign new_n2699_ = ~\b[17]  & ~new_n2698_;
  assign new_n2700_ = \b[17]  & ~new_n2692_;
  assign new_n2701_ = ~new_n2697_ & new_n2700_;
  assign new_n2702_ = new_n270_ & new_n309_;
  assign new_n2703_ = new_n343_ & new_n2702_;
  assign new_n2704_ = new_n341_ & new_n2703_;
  assign new_n2705_ = new_n338_ & new_n2704_;
  assign new_n2706_ = ~new_n2701_ & new_n2705_;
  assign new_n2707_ = ~new_n2699_ & new_n2706_;
  assign new_n2708_ = ~new_n2691_ & new_n2707_;
  assign new_n2709_ = new_n475_ & ~new_n2698_;
  assign \quotient[46]  = new_n2708_ | new_n2709_;
  assign new_n2711_ = ~new_n2479_ & new_n2689_;
  assign new_n2712_ = ~new_n2685_ & new_n2711_;
  assign new_n2713_ = ~new_n2686_ & ~new_n2689_;
  assign new_n2714_ = ~new_n2712_ & ~new_n2713_;
  assign new_n2715_ = \quotient[46]  & ~new_n2714_;
  assign new_n2716_ = ~new_n2469_ & ~new_n2709_;
  assign new_n2717_ = ~new_n2708_ & new_n2716_;
  assign new_n2718_ = ~new_n2715_ & ~new_n2717_;
  assign new_n2719_ = ~new_n2470_ & ~new_n2701_;
  assign new_n2720_ = ~new_n2699_ & new_n2719_;
  assign new_n2721_ = ~new_n2690_ & new_n2720_;
  assign new_n2722_ = ~new_n2699_ & ~new_n2701_;
  assign new_n2723_ = ~new_n2691_ & ~new_n2722_;
  assign new_n2724_ = ~new_n2721_ & ~new_n2723_;
  assign new_n2725_ = \quotient[46]  & ~new_n2724_;
  assign new_n2726_ = ~new_n2698_ & ~new_n2709_;
  assign new_n2727_ = ~new_n2708_ & new_n2726_;
  assign new_n2728_ = ~new_n2725_ & ~new_n2727_;
  assign new_n2729_ = ~\b[18]  & ~new_n2728_;
  assign new_n2730_ = ~\b[17]  & ~new_n2718_;
  assign new_n2731_ = ~new_n2488_ & new_n2684_;
  assign new_n2732_ = ~new_n2680_ & new_n2731_;
  assign new_n2733_ = ~new_n2681_ & ~new_n2684_;
  assign new_n2734_ = ~new_n2732_ & ~new_n2733_;
  assign new_n2735_ = \quotient[46]  & ~new_n2734_;
  assign new_n2736_ = ~new_n2478_ & ~new_n2709_;
  assign new_n2737_ = ~new_n2708_ & new_n2736_;
  assign new_n2738_ = ~new_n2735_ & ~new_n2737_;
  assign new_n2739_ = ~\b[16]  & ~new_n2738_;
  assign new_n2740_ = ~new_n2497_ & new_n2679_;
  assign new_n2741_ = ~new_n2675_ & new_n2740_;
  assign new_n2742_ = ~new_n2676_ & ~new_n2679_;
  assign new_n2743_ = ~new_n2741_ & ~new_n2742_;
  assign new_n2744_ = \quotient[46]  & ~new_n2743_;
  assign new_n2745_ = ~new_n2487_ & ~new_n2709_;
  assign new_n2746_ = ~new_n2708_ & new_n2745_;
  assign new_n2747_ = ~new_n2744_ & ~new_n2746_;
  assign new_n2748_ = ~\b[15]  & ~new_n2747_;
  assign new_n2749_ = ~new_n2506_ & new_n2674_;
  assign new_n2750_ = ~new_n2670_ & new_n2749_;
  assign new_n2751_ = ~new_n2671_ & ~new_n2674_;
  assign new_n2752_ = ~new_n2750_ & ~new_n2751_;
  assign new_n2753_ = \quotient[46]  & ~new_n2752_;
  assign new_n2754_ = ~new_n2496_ & ~new_n2709_;
  assign new_n2755_ = ~new_n2708_ & new_n2754_;
  assign new_n2756_ = ~new_n2753_ & ~new_n2755_;
  assign new_n2757_ = ~\b[14]  & ~new_n2756_;
  assign new_n2758_ = ~new_n2515_ & new_n2669_;
  assign new_n2759_ = ~new_n2665_ & new_n2758_;
  assign new_n2760_ = ~new_n2666_ & ~new_n2669_;
  assign new_n2761_ = ~new_n2759_ & ~new_n2760_;
  assign new_n2762_ = \quotient[46]  & ~new_n2761_;
  assign new_n2763_ = ~new_n2505_ & ~new_n2709_;
  assign new_n2764_ = ~new_n2708_ & new_n2763_;
  assign new_n2765_ = ~new_n2762_ & ~new_n2764_;
  assign new_n2766_ = ~\b[13]  & ~new_n2765_;
  assign new_n2767_ = ~new_n2524_ & new_n2664_;
  assign new_n2768_ = ~new_n2660_ & new_n2767_;
  assign new_n2769_ = ~new_n2661_ & ~new_n2664_;
  assign new_n2770_ = ~new_n2768_ & ~new_n2769_;
  assign new_n2771_ = \quotient[46]  & ~new_n2770_;
  assign new_n2772_ = ~new_n2514_ & ~new_n2709_;
  assign new_n2773_ = ~new_n2708_ & new_n2772_;
  assign new_n2774_ = ~new_n2771_ & ~new_n2773_;
  assign new_n2775_ = ~\b[12]  & ~new_n2774_;
  assign new_n2776_ = ~new_n2533_ & new_n2659_;
  assign new_n2777_ = ~new_n2655_ & new_n2776_;
  assign new_n2778_ = ~new_n2656_ & ~new_n2659_;
  assign new_n2779_ = ~new_n2777_ & ~new_n2778_;
  assign new_n2780_ = \quotient[46]  & ~new_n2779_;
  assign new_n2781_ = ~new_n2523_ & ~new_n2709_;
  assign new_n2782_ = ~new_n2708_ & new_n2781_;
  assign new_n2783_ = ~new_n2780_ & ~new_n2782_;
  assign new_n2784_ = ~\b[11]  & ~new_n2783_;
  assign new_n2785_ = ~new_n2542_ & new_n2654_;
  assign new_n2786_ = ~new_n2650_ & new_n2785_;
  assign new_n2787_ = ~new_n2651_ & ~new_n2654_;
  assign new_n2788_ = ~new_n2786_ & ~new_n2787_;
  assign new_n2789_ = \quotient[46]  & ~new_n2788_;
  assign new_n2790_ = ~new_n2532_ & ~new_n2709_;
  assign new_n2791_ = ~new_n2708_ & new_n2790_;
  assign new_n2792_ = ~new_n2789_ & ~new_n2791_;
  assign new_n2793_ = ~\b[10]  & ~new_n2792_;
  assign new_n2794_ = ~new_n2551_ & new_n2649_;
  assign new_n2795_ = ~new_n2645_ & new_n2794_;
  assign new_n2796_ = ~new_n2646_ & ~new_n2649_;
  assign new_n2797_ = ~new_n2795_ & ~new_n2796_;
  assign new_n2798_ = \quotient[46]  & ~new_n2797_;
  assign new_n2799_ = ~new_n2541_ & ~new_n2709_;
  assign new_n2800_ = ~new_n2708_ & new_n2799_;
  assign new_n2801_ = ~new_n2798_ & ~new_n2800_;
  assign new_n2802_ = ~\b[9]  & ~new_n2801_;
  assign new_n2803_ = ~new_n2560_ & new_n2644_;
  assign new_n2804_ = ~new_n2640_ & new_n2803_;
  assign new_n2805_ = ~new_n2641_ & ~new_n2644_;
  assign new_n2806_ = ~new_n2804_ & ~new_n2805_;
  assign new_n2807_ = \quotient[46]  & ~new_n2806_;
  assign new_n2808_ = ~new_n2550_ & ~new_n2709_;
  assign new_n2809_ = ~new_n2708_ & new_n2808_;
  assign new_n2810_ = ~new_n2807_ & ~new_n2809_;
  assign new_n2811_ = ~\b[8]  & ~new_n2810_;
  assign new_n2812_ = ~new_n2569_ & new_n2639_;
  assign new_n2813_ = ~new_n2635_ & new_n2812_;
  assign new_n2814_ = ~new_n2636_ & ~new_n2639_;
  assign new_n2815_ = ~new_n2813_ & ~new_n2814_;
  assign new_n2816_ = \quotient[46]  & ~new_n2815_;
  assign new_n2817_ = ~new_n2559_ & ~new_n2709_;
  assign new_n2818_ = ~new_n2708_ & new_n2817_;
  assign new_n2819_ = ~new_n2816_ & ~new_n2818_;
  assign new_n2820_ = ~\b[7]  & ~new_n2819_;
  assign new_n2821_ = ~new_n2578_ & new_n2634_;
  assign new_n2822_ = ~new_n2630_ & new_n2821_;
  assign new_n2823_ = ~new_n2631_ & ~new_n2634_;
  assign new_n2824_ = ~new_n2822_ & ~new_n2823_;
  assign new_n2825_ = \quotient[46]  & ~new_n2824_;
  assign new_n2826_ = ~new_n2568_ & ~new_n2709_;
  assign new_n2827_ = ~new_n2708_ & new_n2826_;
  assign new_n2828_ = ~new_n2825_ & ~new_n2827_;
  assign new_n2829_ = ~\b[6]  & ~new_n2828_;
  assign new_n2830_ = ~new_n2587_ & new_n2629_;
  assign new_n2831_ = ~new_n2625_ & new_n2830_;
  assign new_n2832_ = ~new_n2626_ & ~new_n2629_;
  assign new_n2833_ = ~new_n2831_ & ~new_n2832_;
  assign new_n2834_ = \quotient[46]  & ~new_n2833_;
  assign new_n2835_ = ~new_n2577_ & ~new_n2709_;
  assign new_n2836_ = ~new_n2708_ & new_n2835_;
  assign new_n2837_ = ~new_n2834_ & ~new_n2836_;
  assign new_n2838_ = ~\b[5]  & ~new_n2837_;
  assign new_n2839_ = ~new_n2595_ & new_n2624_;
  assign new_n2840_ = ~new_n2620_ & new_n2839_;
  assign new_n2841_ = ~new_n2621_ & ~new_n2624_;
  assign new_n2842_ = ~new_n2840_ & ~new_n2841_;
  assign new_n2843_ = \quotient[46]  & ~new_n2842_;
  assign new_n2844_ = ~new_n2586_ & ~new_n2709_;
  assign new_n2845_ = ~new_n2708_ & new_n2844_;
  assign new_n2846_ = ~new_n2843_ & ~new_n2845_;
  assign new_n2847_ = ~\b[4]  & ~new_n2846_;
  assign new_n2848_ = ~new_n2615_ & new_n2619_;
  assign new_n2849_ = ~new_n2614_ & new_n2848_;
  assign new_n2850_ = ~new_n2616_ & ~new_n2619_;
  assign new_n2851_ = ~new_n2849_ & ~new_n2850_;
  assign new_n2852_ = \quotient[46]  & ~new_n2851_;
  assign new_n2853_ = ~new_n2594_ & ~new_n2709_;
  assign new_n2854_ = ~new_n2708_ & new_n2853_;
  assign new_n2855_ = ~new_n2852_ & ~new_n2854_;
  assign new_n2856_ = ~\b[3]  & ~new_n2855_;
  assign new_n2857_ = ~new_n2611_ & new_n2613_;
  assign new_n2858_ = ~new_n2609_ & new_n2857_;
  assign new_n2859_ = ~new_n2614_ & ~new_n2858_;
  assign new_n2860_ = \quotient[46]  & new_n2859_;
  assign new_n2861_ = ~new_n2608_ & ~new_n2709_;
  assign new_n2862_ = ~new_n2708_ & new_n2861_;
  assign new_n2863_ = ~new_n2860_ & ~new_n2862_;
  assign new_n2864_ = ~\b[2]  & ~new_n2863_;
  assign new_n2865_ = \b[0]  & \quotient[46] ;
  assign new_n2866_ = \a[46]  & ~new_n2865_;
  assign new_n2867_ = new_n2613_ & \quotient[46] ;
  assign new_n2868_ = ~new_n2866_ & ~new_n2867_;
  assign new_n2869_ = \b[1]  & ~new_n2868_;
  assign new_n2870_ = ~\b[1]  & ~new_n2867_;
  assign new_n2871_ = ~new_n2866_ & new_n2870_;
  assign new_n2872_ = ~new_n2869_ & ~new_n2871_;
  assign new_n2873_ = ~\a[45]  & \b[0] ;
  assign new_n2874_ = ~new_n2872_ & ~new_n2873_;
  assign new_n2875_ = ~\b[1]  & ~new_n2868_;
  assign new_n2876_ = ~new_n2874_ & ~new_n2875_;
  assign new_n2877_ = \b[2]  & ~new_n2862_;
  assign new_n2878_ = ~new_n2860_ & new_n2877_;
  assign new_n2879_ = ~new_n2864_ & ~new_n2878_;
  assign new_n2880_ = ~new_n2876_ & new_n2879_;
  assign new_n2881_ = ~new_n2864_ & ~new_n2880_;
  assign new_n2882_ = \b[3]  & ~new_n2854_;
  assign new_n2883_ = ~new_n2852_ & new_n2882_;
  assign new_n2884_ = ~new_n2856_ & ~new_n2883_;
  assign new_n2885_ = ~new_n2881_ & new_n2884_;
  assign new_n2886_ = ~new_n2856_ & ~new_n2885_;
  assign new_n2887_ = \b[4]  & ~new_n2845_;
  assign new_n2888_ = ~new_n2843_ & new_n2887_;
  assign new_n2889_ = ~new_n2847_ & ~new_n2888_;
  assign new_n2890_ = ~new_n2886_ & new_n2889_;
  assign new_n2891_ = ~new_n2847_ & ~new_n2890_;
  assign new_n2892_ = \b[5]  & ~new_n2836_;
  assign new_n2893_ = ~new_n2834_ & new_n2892_;
  assign new_n2894_ = ~new_n2838_ & ~new_n2893_;
  assign new_n2895_ = ~new_n2891_ & new_n2894_;
  assign new_n2896_ = ~new_n2838_ & ~new_n2895_;
  assign new_n2897_ = \b[6]  & ~new_n2827_;
  assign new_n2898_ = ~new_n2825_ & new_n2897_;
  assign new_n2899_ = ~new_n2829_ & ~new_n2898_;
  assign new_n2900_ = ~new_n2896_ & new_n2899_;
  assign new_n2901_ = ~new_n2829_ & ~new_n2900_;
  assign new_n2902_ = \b[7]  & ~new_n2818_;
  assign new_n2903_ = ~new_n2816_ & new_n2902_;
  assign new_n2904_ = ~new_n2820_ & ~new_n2903_;
  assign new_n2905_ = ~new_n2901_ & new_n2904_;
  assign new_n2906_ = ~new_n2820_ & ~new_n2905_;
  assign new_n2907_ = \b[8]  & ~new_n2809_;
  assign new_n2908_ = ~new_n2807_ & new_n2907_;
  assign new_n2909_ = ~new_n2811_ & ~new_n2908_;
  assign new_n2910_ = ~new_n2906_ & new_n2909_;
  assign new_n2911_ = ~new_n2811_ & ~new_n2910_;
  assign new_n2912_ = \b[9]  & ~new_n2800_;
  assign new_n2913_ = ~new_n2798_ & new_n2912_;
  assign new_n2914_ = ~new_n2802_ & ~new_n2913_;
  assign new_n2915_ = ~new_n2911_ & new_n2914_;
  assign new_n2916_ = ~new_n2802_ & ~new_n2915_;
  assign new_n2917_ = \b[10]  & ~new_n2791_;
  assign new_n2918_ = ~new_n2789_ & new_n2917_;
  assign new_n2919_ = ~new_n2793_ & ~new_n2918_;
  assign new_n2920_ = ~new_n2916_ & new_n2919_;
  assign new_n2921_ = ~new_n2793_ & ~new_n2920_;
  assign new_n2922_ = \b[11]  & ~new_n2782_;
  assign new_n2923_ = ~new_n2780_ & new_n2922_;
  assign new_n2924_ = ~new_n2784_ & ~new_n2923_;
  assign new_n2925_ = ~new_n2921_ & new_n2924_;
  assign new_n2926_ = ~new_n2784_ & ~new_n2925_;
  assign new_n2927_ = \b[12]  & ~new_n2773_;
  assign new_n2928_ = ~new_n2771_ & new_n2927_;
  assign new_n2929_ = ~new_n2775_ & ~new_n2928_;
  assign new_n2930_ = ~new_n2926_ & new_n2929_;
  assign new_n2931_ = ~new_n2775_ & ~new_n2930_;
  assign new_n2932_ = \b[13]  & ~new_n2764_;
  assign new_n2933_ = ~new_n2762_ & new_n2932_;
  assign new_n2934_ = ~new_n2766_ & ~new_n2933_;
  assign new_n2935_ = ~new_n2931_ & new_n2934_;
  assign new_n2936_ = ~new_n2766_ & ~new_n2935_;
  assign new_n2937_ = \b[14]  & ~new_n2755_;
  assign new_n2938_ = ~new_n2753_ & new_n2937_;
  assign new_n2939_ = ~new_n2757_ & ~new_n2938_;
  assign new_n2940_ = ~new_n2936_ & new_n2939_;
  assign new_n2941_ = ~new_n2757_ & ~new_n2940_;
  assign new_n2942_ = \b[15]  & ~new_n2746_;
  assign new_n2943_ = ~new_n2744_ & new_n2942_;
  assign new_n2944_ = ~new_n2748_ & ~new_n2943_;
  assign new_n2945_ = ~new_n2941_ & new_n2944_;
  assign new_n2946_ = ~new_n2748_ & ~new_n2945_;
  assign new_n2947_ = \b[16]  & ~new_n2737_;
  assign new_n2948_ = ~new_n2735_ & new_n2947_;
  assign new_n2949_ = ~new_n2739_ & ~new_n2948_;
  assign new_n2950_ = ~new_n2946_ & new_n2949_;
  assign new_n2951_ = ~new_n2739_ & ~new_n2950_;
  assign new_n2952_ = \b[17]  & ~new_n2717_;
  assign new_n2953_ = ~new_n2715_ & new_n2952_;
  assign new_n2954_ = ~new_n2730_ & ~new_n2953_;
  assign new_n2955_ = ~new_n2951_ & new_n2954_;
  assign new_n2956_ = ~new_n2730_ & ~new_n2955_;
  assign new_n2957_ = \b[18]  & ~new_n2727_;
  assign new_n2958_ = ~new_n2725_ & new_n2957_;
  assign new_n2959_ = ~new_n2729_ & ~new_n2958_;
  assign new_n2960_ = ~new_n2956_ & new_n2959_;
  assign new_n2961_ = ~new_n2729_ & ~new_n2960_;
  assign new_n2962_ = new_n366_ & new_n368_;
  assign new_n2963_ = new_n377_ & new_n2962_;
  assign new_n2964_ = new_n423_ & new_n2963_;
  assign new_n2965_ = new_n408_ & new_n2964_;
  assign \quotient[45]  = ~new_n2961_ & new_n2965_;
  assign new_n2967_ = ~new_n2718_ & ~\quotient[45] ;
  assign new_n2968_ = ~new_n2739_ & new_n2954_;
  assign new_n2969_ = ~new_n2950_ & new_n2968_;
  assign new_n2970_ = ~new_n2951_ & ~new_n2954_;
  assign new_n2971_ = ~new_n2969_ & ~new_n2970_;
  assign new_n2972_ = new_n2965_ & ~new_n2971_;
  assign new_n2973_ = ~new_n2961_ & new_n2972_;
  assign new_n2974_ = ~new_n2967_ & ~new_n2973_;
  assign new_n2975_ = ~new_n2728_ & ~\quotient[45] ;
  assign new_n2976_ = ~new_n2730_ & new_n2959_;
  assign new_n2977_ = ~new_n2955_ & new_n2976_;
  assign new_n2978_ = ~new_n2956_ & ~new_n2959_;
  assign new_n2979_ = ~new_n2977_ & ~new_n2978_;
  assign new_n2980_ = \quotient[45]  & ~new_n2979_;
  assign new_n2981_ = ~new_n2975_ & ~new_n2980_;
  assign new_n2982_ = ~\b[19]  & ~new_n2981_;
  assign new_n2983_ = ~\b[18]  & ~new_n2974_;
  assign new_n2984_ = ~new_n2738_ & ~\quotient[45] ;
  assign new_n2985_ = ~new_n2748_ & new_n2949_;
  assign new_n2986_ = ~new_n2945_ & new_n2985_;
  assign new_n2987_ = ~new_n2946_ & ~new_n2949_;
  assign new_n2988_ = ~new_n2986_ & ~new_n2987_;
  assign new_n2989_ = new_n2965_ & ~new_n2988_;
  assign new_n2990_ = ~new_n2961_ & new_n2989_;
  assign new_n2991_ = ~new_n2984_ & ~new_n2990_;
  assign new_n2992_ = ~\b[17]  & ~new_n2991_;
  assign new_n2993_ = ~new_n2747_ & ~\quotient[45] ;
  assign new_n2994_ = ~new_n2757_ & new_n2944_;
  assign new_n2995_ = ~new_n2940_ & new_n2994_;
  assign new_n2996_ = ~new_n2941_ & ~new_n2944_;
  assign new_n2997_ = ~new_n2995_ & ~new_n2996_;
  assign new_n2998_ = new_n2965_ & ~new_n2997_;
  assign new_n2999_ = ~new_n2961_ & new_n2998_;
  assign new_n3000_ = ~new_n2993_ & ~new_n2999_;
  assign new_n3001_ = ~\b[16]  & ~new_n3000_;
  assign new_n3002_ = ~new_n2756_ & ~\quotient[45] ;
  assign new_n3003_ = ~new_n2766_ & new_n2939_;
  assign new_n3004_ = ~new_n2935_ & new_n3003_;
  assign new_n3005_ = ~new_n2936_ & ~new_n2939_;
  assign new_n3006_ = ~new_n3004_ & ~new_n3005_;
  assign new_n3007_ = new_n2965_ & ~new_n3006_;
  assign new_n3008_ = ~new_n2961_ & new_n3007_;
  assign new_n3009_ = ~new_n3002_ & ~new_n3008_;
  assign new_n3010_ = ~\b[15]  & ~new_n3009_;
  assign new_n3011_ = ~new_n2765_ & ~\quotient[45] ;
  assign new_n3012_ = ~new_n2775_ & new_n2934_;
  assign new_n3013_ = ~new_n2930_ & new_n3012_;
  assign new_n3014_ = ~new_n2931_ & ~new_n2934_;
  assign new_n3015_ = ~new_n3013_ & ~new_n3014_;
  assign new_n3016_ = new_n2965_ & ~new_n3015_;
  assign new_n3017_ = ~new_n2961_ & new_n3016_;
  assign new_n3018_ = ~new_n3011_ & ~new_n3017_;
  assign new_n3019_ = ~\b[14]  & ~new_n3018_;
  assign new_n3020_ = ~new_n2774_ & ~\quotient[45] ;
  assign new_n3021_ = ~new_n2784_ & new_n2929_;
  assign new_n3022_ = ~new_n2925_ & new_n3021_;
  assign new_n3023_ = ~new_n2926_ & ~new_n2929_;
  assign new_n3024_ = ~new_n3022_ & ~new_n3023_;
  assign new_n3025_ = new_n2965_ & ~new_n3024_;
  assign new_n3026_ = ~new_n2961_ & new_n3025_;
  assign new_n3027_ = ~new_n3020_ & ~new_n3026_;
  assign new_n3028_ = ~\b[13]  & ~new_n3027_;
  assign new_n3029_ = ~new_n2783_ & ~\quotient[45] ;
  assign new_n3030_ = ~new_n2793_ & new_n2924_;
  assign new_n3031_ = ~new_n2920_ & new_n3030_;
  assign new_n3032_ = ~new_n2921_ & ~new_n2924_;
  assign new_n3033_ = ~new_n3031_ & ~new_n3032_;
  assign new_n3034_ = new_n2965_ & ~new_n3033_;
  assign new_n3035_ = ~new_n2961_ & new_n3034_;
  assign new_n3036_ = ~new_n3029_ & ~new_n3035_;
  assign new_n3037_ = ~\b[12]  & ~new_n3036_;
  assign new_n3038_ = ~new_n2792_ & ~\quotient[45] ;
  assign new_n3039_ = ~new_n2802_ & new_n2919_;
  assign new_n3040_ = ~new_n2915_ & new_n3039_;
  assign new_n3041_ = ~new_n2916_ & ~new_n2919_;
  assign new_n3042_ = ~new_n3040_ & ~new_n3041_;
  assign new_n3043_ = new_n2965_ & ~new_n3042_;
  assign new_n3044_ = ~new_n2961_ & new_n3043_;
  assign new_n3045_ = ~new_n3038_ & ~new_n3044_;
  assign new_n3046_ = ~\b[11]  & ~new_n3045_;
  assign new_n3047_ = ~new_n2801_ & ~\quotient[45] ;
  assign new_n3048_ = ~new_n2811_ & new_n2914_;
  assign new_n3049_ = ~new_n2910_ & new_n3048_;
  assign new_n3050_ = ~new_n2911_ & ~new_n2914_;
  assign new_n3051_ = ~new_n3049_ & ~new_n3050_;
  assign new_n3052_ = new_n2965_ & ~new_n3051_;
  assign new_n3053_ = ~new_n2961_ & new_n3052_;
  assign new_n3054_ = ~new_n3047_ & ~new_n3053_;
  assign new_n3055_ = ~\b[10]  & ~new_n3054_;
  assign new_n3056_ = ~new_n2810_ & ~\quotient[45] ;
  assign new_n3057_ = ~new_n2820_ & new_n2909_;
  assign new_n3058_ = ~new_n2905_ & new_n3057_;
  assign new_n3059_ = ~new_n2906_ & ~new_n2909_;
  assign new_n3060_ = ~new_n3058_ & ~new_n3059_;
  assign new_n3061_ = new_n2965_ & ~new_n3060_;
  assign new_n3062_ = ~new_n2961_ & new_n3061_;
  assign new_n3063_ = ~new_n3056_ & ~new_n3062_;
  assign new_n3064_ = ~\b[9]  & ~new_n3063_;
  assign new_n3065_ = ~new_n2819_ & ~\quotient[45] ;
  assign new_n3066_ = ~new_n2829_ & new_n2904_;
  assign new_n3067_ = ~new_n2900_ & new_n3066_;
  assign new_n3068_ = ~new_n2901_ & ~new_n2904_;
  assign new_n3069_ = ~new_n3067_ & ~new_n3068_;
  assign new_n3070_ = new_n2965_ & ~new_n3069_;
  assign new_n3071_ = ~new_n2961_ & new_n3070_;
  assign new_n3072_ = ~new_n3065_ & ~new_n3071_;
  assign new_n3073_ = ~\b[8]  & ~new_n3072_;
  assign new_n3074_ = ~new_n2828_ & ~\quotient[45] ;
  assign new_n3075_ = ~new_n2838_ & new_n2899_;
  assign new_n3076_ = ~new_n2895_ & new_n3075_;
  assign new_n3077_ = ~new_n2896_ & ~new_n2899_;
  assign new_n3078_ = ~new_n3076_ & ~new_n3077_;
  assign new_n3079_ = new_n2965_ & ~new_n3078_;
  assign new_n3080_ = ~new_n2961_ & new_n3079_;
  assign new_n3081_ = ~new_n3074_ & ~new_n3080_;
  assign new_n3082_ = ~\b[7]  & ~new_n3081_;
  assign new_n3083_ = ~new_n2837_ & ~\quotient[45] ;
  assign new_n3084_ = ~new_n2847_ & new_n2894_;
  assign new_n3085_ = ~new_n2890_ & new_n3084_;
  assign new_n3086_ = ~new_n2891_ & ~new_n2894_;
  assign new_n3087_ = ~new_n3085_ & ~new_n3086_;
  assign new_n3088_ = new_n2965_ & ~new_n3087_;
  assign new_n3089_ = ~new_n2961_ & new_n3088_;
  assign new_n3090_ = ~new_n3083_ & ~new_n3089_;
  assign new_n3091_ = ~\b[6]  & ~new_n3090_;
  assign new_n3092_ = ~new_n2846_ & ~\quotient[45] ;
  assign new_n3093_ = ~new_n2856_ & new_n2889_;
  assign new_n3094_ = ~new_n2885_ & new_n3093_;
  assign new_n3095_ = ~new_n2886_ & ~new_n2889_;
  assign new_n3096_ = ~new_n3094_ & ~new_n3095_;
  assign new_n3097_ = new_n2965_ & ~new_n3096_;
  assign new_n3098_ = ~new_n2961_ & new_n3097_;
  assign new_n3099_ = ~new_n3092_ & ~new_n3098_;
  assign new_n3100_ = ~\b[5]  & ~new_n3099_;
  assign new_n3101_ = ~new_n2855_ & ~\quotient[45] ;
  assign new_n3102_ = ~new_n2864_ & new_n2884_;
  assign new_n3103_ = ~new_n2880_ & new_n3102_;
  assign new_n3104_ = ~new_n2881_ & ~new_n2884_;
  assign new_n3105_ = ~new_n3103_ & ~new_n3104_;
  assign new_n3106_ = new_n2965_ & ~new_n3105_;
  assign new_n3107_ = ~new_n2961_ & new_n3106_;
  assign new_n3108_ = ~new_n3101_ & ~new_n3107_;
  assign new_n3109_ = ~\b[4]  & ~new_n3108_;
  assign new_n3110_ = ~new_n2863_ & ~\quotient[45] ;
  assign new_n3111_ = ~new_n2875_ & new_n2879_;
  assign new_n3112_ = ~new_n2874_ & new_n3111_;
  assign new_n3113_ = ~new_n2876_ & ~new_n2879_;
  assign new_n3114_ = ~new_n3112_ & ~new_n3113_;
  assign new_n3115_ = new_n2965_ & ~new_n3114_;
  assign new_n3116_ = ~new_n2961_ & new_n3115_;
  assign new_n3117_ = ~new_n3110_ & ~new_n3116_;
  assign new_n3118_ = ~\b[3]  & ~new_n3117_;
  assign new_n3119_ = ~new_n2868_ & ~\quotient[45] ;
  assign new_n3120_ = ~new_n2871_ & new_n2873_;
  assign new_n3121_ = ~new_n2869_ & new_n3120_;
  assign new_n3122_ = new_n2965_ & ~new_n3121_;
  assign new_n3123_ = ~new_n2874_ & new_n3122_;
  assign new_n3124_ = ~new_n2961_ & new_n3123_;
  assign new_n3125_ = ~new_n3119_ & ~new_n3124_;
  assign new_n3126_ = ~\b[2]  & ~new_n3125_;
  assign new_n3127_ = \b[0]  & ~\b[19] ;
  assign new_n3128_ = new_n309_ & new_n3127_;
  assign new_n3129_ = new_n343_ & new_n3128_;
  assign new_n3130_ = new_n341_ & new_n3129_;
  assign new_n3131_ = new_n338_ & new_n3130_;
  assign new_n3132_ = ~new_n2961_ & new_n3131_;
  assign new_n3133_ = \a[45]  & ~new_n3132_;
  assign new_n3134_ = new_n368_ & new_n2873_;
  assign new_n3135_ = new_n366_ & new_n3134_;
  assign new_n3136_ = new_n377_ & new_n3135_;
  assign new_n3137_ = new_n423_ & new_n3136_;
  assign new_n3138_ = new_n408_ & new_n3137_;
  assign new_n3139_ = ~new_n2961_ & new_n3138_;
  assign new_n3140_ = ~new_n3133_ & ~new_n3139_;
  assign new_n3141_ = \b[1]  & ~new_n3140_;
  assign new_n3142_ = ~\b[1]  & ~new_n3139_;
  assign new_n3143_ = ~new_n3133_ & new_n3142_;
  assign new_n3144_ = ~new_n3141_ & ~new_n3143_;
  assign new_n3145_ = ~\a[44]  & \b[0] ;
  assign new_n3146_ = ~new_n3144_ & ~new_n3145_;
  assign new_n3147_ = ~\b[1]  & ~new_n3140_;
  assign new_n3148_ = ~new_n3146_ & ~new_n3147_;
  assign new_n3149_ = \b[2]  & ~new_n3124_;
  assign new_n3150_ = ~new_n3119_ & new_n3149_;
  assign new_n3151_ = ~new_n3126_ & ~new_n3150_;
  assign new_n3152_ = ~new_n3148_ & new_n3151_;
  assign new_n3153_ = ~new_n3126_ & ~new_n3152_;
  assign new_n3154_ = \b[3]  & ~new_n3116_;
  assign new_n3155_ = ~new_n3110_ & new_n3154_;
  assign new_n3156_ = ~new_n3118_ & ~new_n3155_;
  assign new_n3157_ = ~new_n3153_ & new_n3156_;
  assign new_n3158_ = ~new_n3118_ & ~new_n3157_;
  assign new_n3159_ = \b[4]  & ~new_n3107_;
  assign new_n3160_ = ~new_n3101_ & new_n3159_;
  assign new_n3161_ = ~new_n3109_ & ~new_n3160_;
  assign new_n3162_ = ~new_n3158_ & new_n3161_;
  assign new_n3163_ = ~new_n3109_ & ~new_n3162_;
  assign new_n3164_ = \b[5]  & ~new_n3098_;
  assign new_n3165_ = ~new_n3092_ & new_n3164_;
  assign new_n3166_ = ~new_n3100_ & ~new_n3165_;
  assign new_n3167_ = ~new_n3163_ & new_n3166_;
  assign new_n3168_ = ~new_n3100_ & ~new_n3167_;
  assign new_n3169_ = \b[6]  & ~new_n3089_;
  assign new_n3170_ = ~new_n3083_ & new_n3169_;
  assign new_n3171_ = ~new_n3091_ & ~new_n3170_;
  assign new_n3172_ = ~new_n3168_ & new_n3171_;
  assign new_n3173_ = ~new_n3091_ & ~new_n3172_;
  assign new_n3174_ = \b[7]  & ~new_n3080_;
  assign new_n3175_ = ~new_n3074_ & new_n3174_;
  assign new_n3176_ = ~new_n3082_ & ~new_n3175_;
  assign new_n3177_ = ~new_n3173_ & new_n3176_;
  assign new_n3178_ = ~new_n3082_ & ~new_n3177_;
  assign new_n3179_ = \b[8]  & ~new_n3071_;
  assign new_n3180_ = ~new_n3065_ & new_n3179_;
  assign new_n3181_ = ~new_n3073_ & ~new_n3180_;
  assign new_n3182_ = ~new_n3178_ & new_n3181_;
  assign new_n3183_ = ~new_n3073_ & ~new_n3182_;
  assign new_n3184_ = \b[9]  & ~new_n3062_;
  assign new_n3185_ = ~new_n3056_ & new_n3184_;
  assign new_n3186_ = ~new_n3064_ & ~new_n3185_;
  assign new_n3187_ = ~new_n3183_ & new_n3186_;
  assign new_n3188_ = ~new_n3064_ & ~new_n3187_;
  assign new_n3189_ = \b[10]  & ~new_n3053_;
  assign new_n3190_ = ~new_n3047_ & new_n3189_;
  assign new_n3191_ = ~new_n3055_ & ~new_n3190_;
  assign new_n3192_ = ~new_n3188_ & new_n3191_;
  assign new_n3193_ = ~new_n3055_ & ~new_n3192_;
  assign new_n3194_ = \b[11]  & ~new_n3044_;
  assign new_n3195_ = ~new_n3038_ & new_n3194_;
  assign new_n3196_ = ~new_n3046_ & ~new_n3195_;
  assign new_n3197_ = ~new_n3193_ & new_n3196_;
  assign new_n3198_ = ~new_n3046_ & ~new_n3197_;
  assign new_n3199_ = \b[12]  & ~new_n3035_;
  assign new_n3200_ = ~new_n3029_ & new_n3199_;
  assign new_n3201_ = ~new_n3037_ & ~new_n3200_;
  assign new_n3202_ = ~new_n3198_ & new_n3201_;
  assign new_n3203_ = ~new_n3037_ & ~new_n3202_;
  assign new_n3204_ = \b[13]  & ~new_n3026_;
  assign new_n3205_ = ~new_n3020_ & new_n3204_;
  assign new_n3206_ = ~new_n3028_ & ~new_n3205_;
  assign new_n3207_ = ~new_n3203_ & new_n3206_;
  assign new_n3208_ = ~new_n3028_ & ~new_n3207_;
  assign new_n3209_ = \b[14]  & ~new_n3017_;
  assign new_n3210_ = ~new_n3011_ & new_n3209_;
  assign new_n3211_ = ~new_n3019_ & ~new_n3210_;
  assign new_n3212_ = ~new_n3208_ & new_n3211_;
  assign new_n3213_ = ~new_n3019_ & ~new_n3212_;
  assign new_n3214_ = \b[15]  & ~new_n3008_;
  assign new_n3215_ = ~new_n3002_ & new_n3214_;
  assign new_n3216_ = ~new_n3010_ & ~new_n3215_;
  assign new_n3217_ = ~new_n3213_ & new_n3216_;
  assign new_n3218_ = ~new_n3010_ & ~new_n3217_;
  assign new_n3219_ = \b[16]  & ~new_n2999_;
  assign new_n3220_ = ~new_n2993_ & new_n3219_;
  assign new_n3221_ = ~new_n3001_ & ~new_n3220_;
  assign new_n3222_ = ~new_n3218_ & new_n3221_;
  assign new_n3223_ = ~new_n3001_ & ~new_n3222_;
  assign new_n3224_ = \b[17]  & ~new_n2990_;
  assign new_n3225_ = ~new_n2984_ & new_n3224_;
  assign new_n3226_ = ~new_n2992_ & ~new_n3225_;
  assign new_n3227_ = ~new_n3223_ & new_n3226_;
  assign new_n3228_ = ~new_n2992_ & ~new_n3227_;
  assign new_n3229_ = \b[18]  & ~new_n2973_;
  assign new_n3230_ = ~new_n2967_ & new_n3229_;
  assign new_n3231_ = ~new_n2983_ & ~new_n3230_;
  assign new_n3232_ = ~new_n3228_ & new_n3231_;
  assign new_n3233_ = ~new_n2983_ & ~new_n3232_;
  assign new_n3234_ = \b[19]  & ~new_n2975_;
  assign new_n3235_ = ~new_n2980_ & new_n3234_;
  assign new_n3236_ = ~new_n2982_ & ~new_n3235_;
  assign new_n3237_ = ~new_n3233_ & new_n3236_;
  assign new_n3238_ = ~new_n2982_ & ~new_n3237_;
  assign \quotient[44]  = new_n320_ & ~new_n3238_;
  assign new_n3240_ = ~new_n2974_ & ~\quotient[44] ;
  assign new_n3241_ = ~new_n2992_ & new_n3231_;
  assign new_n3242_ = ~new_n3227_ & new_n3241_;
  assign new_n3243_ = ~new_n3228_ & ~new_n3231_;
  assign new_n3244_ = ~new_n3242_ & ~new_n3243_;
  assign new_n3245_ = new_n320_ & ~new_n3244_;
  assign new_n3246_ = ~new_n3238_ & new_n3245_;
  assign new_n3247_ = ~new_n3240_ & ~new_n3246_;
  assign new_n3248_ = ~\b[19]  & ~new_n3247_;
  assign new_n3249_ = ~new_n2991_ & ~\quotient[44] ;
  assign new_n3250_ = ~new_n3001_ & new_n3226_;
  assign new_n3251_ = ~new_n3222_ & new_n3250_;
  assign new_n3252_ = ~new_n3223_ & ~new_n3226_;
  assign new_n3253_ = ~new_n3251_ & ~new_n3252_;
  assign new_n3254_ = new_n320_ & ~new_n3253_;
  assign new_n3255_ = ~new_n3238_ & new_n3254_;
  assign new_n3256_ = ~new_n3249_ & ~new_n3255_;
  assign new_n3257_ = ~\b[18]  & ~new_n3256_;
  assign new_n3258_ = ~new_n3000_ & ~\quotient[44] ;
  assign new_n3259_ = ~new_n3010_ & new_n3221_;
  assign new_n3260_ = ~new_n3217_ & new_n3259_;
  assign new_n3261_ = ~new_n3218_ & ~new_n3221_;
  assign new_n3262_ = ~new_n3260_ & ~new_n3261_;
  assign new_n3263_ = new_n320_ & ~new_n3262_;
  assign new_n3264_ = ~new_n3238_ & new_n3263_;
  assign new_n3265_ = ~new_n3258_ & ~new_n3264_;
  assign new_n3266_ = ~\b[17]  & ~new_n3265_;
  assign new_n3267_ = ~new_n3009_ & ~\quotient[44] ;
  assign new_n3268_ = ~new_n3019_ & new_n3216_;
  assign new_n3269_ = ~new_n3212_ & new_n3268_;
  assign new_n3270_ = ~new_n3213_ & ~new_n3216_;
  assign new_n3271_ = ~new_n3269_ & ~new_n3270_;
  assign new_n3272_ = new_n320_ & ~new_n3271_;
  assign new_n3273_ = ~new_n3238_ & new_n3272_;
  assign new_n3274_ = ~new_n3267_ & ~new_n3273_;
  assign new_n3275_ = ~\b[16]  & ~new_n3274_;
  assign new_n3276_ = ~new_n3018_ & ~\quotient[44] ;
  assign new_n3277_ = ~new_n3028_ & new_n3211_;
  assign new_n3278_ = ~new_n3207_ & new_n3277_;
  assign new_n3279_ = ~new_n3208_ & ~new_n3211_;
  assign new_n3280_ = ~new_n3278_ & ~new_n3279_;
  assign new_n3281_ = new_n320_ & ~new_n3280_;
  assign new_n3282_ = ~new_n3238_ & new_n3281_;
  assign new_n3283_ = ~new_n3276_ & ~new_n3282_;
  assign new_n3284_ = ~\b[15]  & ~new_n3283_;
  assign new_n3285_ = ~new_n3027_ & ~\quotient[44] ;
  assign new_n3286_ = ~new_n3037_ & new_n3206_;
  assign new_n3287_ = ~new_n3202_ & new_n3286_;
  assign new_n3288_ = ~new_n3203_ & ~new_n3206_;
  assign new_n3289_ = ~new_n3287_ & ~new_n3288_;
  assign new_n3290_ = new_n320_ & ~new_n3289_;
  assign new_n3291_ = ~new_n3238_ & new_n3290_;
  assign new_n3292_ = ~new_n3285_ & ~new_n3291_;
  assign new_n3293_ = ~\b[14]  & ~new_n3292_;
  assign new_n3294_ = ~new_n3036_ & ~\quotient[44] ;
  assign new_n3295_ = ~new_n3046_ & new_n3201_;
  assign new_n3296_ = ~new_n3197_ & new_n3295_;
  assign new_n3297_ = ~new_n3198_ & ~new_n3201_;
  assign new_n3298_ = ~new_n3296_ & ~new_n3297_;
  assign new_n3299_ = new_n320_ & ~new_n3298_;
  assign new_n3300_ = ~new_n3238_ & new_n3299_;
  assign new_n3301_ = ~new_n3294_ & ~new_n3300_;
  assign new_n3302_ = ~\b[13]  & ~new_n3301_;
  assign new_n3303_ = ~new_n3045_ & ~\quotient[44] ;
  assign new_n3304_ = ~new_n3055_ & new_n3196_;
  assign new_n3305_ = ~new_n3192_ & new_n3304_;
  assign new_n3306_ = ~new_n3193_ & ~new_n3196_;
  assign new_n3307_ = ~new_n3305_ & ~new_n3306_;
  assign new_n3308_ = new_n320_ & ~new_n3307_;
  assign new_n3309_ = ~new_n3238_ & new_n3308_;
  assign new_n3310_ = ~new_n3303_ & ~new_n3309_;
  assign new_n3311_ = ~\b[12]  & ~new_n3310_;
  assign new_n3312_ = ~new_n3054_ & ~\quotient[44] ;
  assign new_n3313_ = ~new_n3064_ & new_n3191_;
  assign new_n3314_ = ~new_n3187_ & new_n3313_;
  assign new_n3315_ = ~new_n3188_ & ~new_n3191_;
  assign new_n3316_ = ~new_n3314_ & ~new_n3315_;
  assign new_n3317_ = new_n320_ & ~new_n3316_;
  assign new_n3318_ = ~new_n3238_ & new_n3317_;
  assign new_n3319_ = ~new_n3312_ & ~new_n3318_;
  assign new_n3320_ = ~\b[11]  & ~new_n3319_;
  assign new_n3321_ = ~new_n3063_ & ~\quotient[44] ;
  assign new_n3322_ = ~new_n3073_ & new_n3186_;
  assign new_n3323_ = ~new_n3182_ & new_n3322_;
  assign new_n3324_ = ~new_n3183_ & ~new_n3186_;
  assign new_n3325_ = ~new_n3323_ & ~new_n3324_;
  assign new_n3326_ = new_n320_ & ~new_n3325_;
  assign new_n3327_ = ~new_n3238_ & new_n3326_;
  assign new_n3328_ = ~new_n3321_ & ~new_n3327_;
  assign new_n3329_ = ~\b[10]  & ~new_n3328_;
  assign new_n3330_ = ~new_n3072_ & ~\quotient[44] ;
  assign new_n3331_ = ~new_n3082_ & new_n3181_;
  assign new_n3332_ = ~new_n3177_ & new_n3331_;
  assign new_n3333_ = ~new_n3178_ & ~new_n3181_;
  assign new_n3334_ = ~new_n3332_ & ~new_n3333_;
  assign new_n3335_ = new_n320_ & ~new_n3334_;
  assign new_n3336_ = ~new_n3238_ & new_n3335_;
  assign new_n3337_ = ~new_n3330_ & ~new_n3336_;
  assign new_n3338_ = ~\b[9]  & ~new_n3337_;
  assign new_n3339_ = ~new_n3081_ & ~\quotient[44] ;
  assign new_n3340_ = ~new_n3091_ & new_n3176_;
  assign new_n3341_ = ~new_n3172_ & new_n3340_;
  assign new_n3342_ = ~new_n3173_ & ~new_n3176_;
  assign new_n3343_ = ~new_n3341_ & ~new_n3342_;
  assign new_n3344_ = new_n320_ & ~new_n3343_;
  assign new_n3345_ = ~new_n3238_ & new_n3344_;
  assign new_n3346_ = ~new_n3339_ & ~new_n3345_;
  assign new_n3347_ = ~\b[8]  & ~new_n3346_;
  assign new_n3348_ = ~new_n3090_ & ~\quotient[44] ;
  assign new_n3349_ = ~new_n3100_ & new_n3171_;
  assign new_n3350_ = ~new_n3167_ & new_n3349_;
  assign new_n3351_ = ~new_n3168_ & ~new_n3171_;
  assign new_n3352_ = ~new_n3350_ & ~new_n3351_;
  assign new_n3353_ = new_n320_ & ~new_n3352_;
  assign new_n3354_ = ~new_n3238_ & new_n3353_;
  assign new_n3355_ = ~new_n3348_ & ~new_n3354_;
  assign new_n3356_ = ~\b[7]  & ~new_n3355_;
  assign new_n3357_ = ~new_n3099_ & ~\quotient[44] ;
  assign new_n3358_ = ~new_n3109_ & new_n3166_;
  assign new_n3359_ = ~new_n3162_ & new_n3358_;
  assign new_n3360_ = ~new_n3163_ & ~new_n3166_;
  assign new_n3361_ = ~new_n3359_ & ~new_n3360_;
  assign new_n3362_ = new_n320_ & ~new_n3361_;
  assign new_n3363_ = ~new_n3238_ & new_n3362_;
  assign new_n3364_ = ~new_n3357_ & ~new_n3363_;
  assign new_n3365_ = ~\b[6]  & ~new_n3364_;
  assign new_n3366_ = ~new_n3108_ & ~\quotient[44] ;
  assign new_n3367_ = ~new_n3118_ & new_n3161_;
  assign new_n3368_ = ~new_n3157_ & new_n3367_;
  assign new_n3369_ = ~new_n3158_ & ~new_n3161_;
  assign new_n3370_ = ~new_n3368_ & ~new_n3369_;
  assign new_n3371_ = new_n320_ & ~new_n3370_;
  assign new_n3372_ = ~new_n3238_ & new_n3371_;
  assign new_n3373_ = ~new_n3366_ & ~new_n3372_;
  assign new_n3374_ = ~\b[5]  & ~new_n3373_;
  assign new_n3375_ = ~new_n3117_ & ~\quotient[44] ;
  assign new_n3376_ = ~new_n3126_ & new_n3156_;
  assign new_n3377_ = ~new_n3152_ & new_n3376_;
  assign new_n3378_ = ~new_n3153_ & ~new_n3156_;
  assign new_n3379_ = ~new_n3377_ & ~new_n3378_;
  assign new_n3380_ = new_n320_ & ~new_n3379_;
  assign new_n3381_ = ~new_n3238_ & new_n3380_;
  assign new_n3382_ = ~new_n3375_ & ~new_n3381_;
  assign new_n3383_ = ~\b[4]  & ~new_n3382_;
  assign new_n3384_ = ~new_n3125_ & ~\quotient[44] ;
  assign new_n3385_ = ~new_n3147_ & new_n3151_;
  assign new_n3386_ = ~new_n3146_ & new_n3385_;
  assign new_n3387_ = ~new_n3148_ & ~new_n3151_;
  assign new_n3388_ = ~new_n3386_ & ~new_n3387_;
  assign new_n3389_ = new_n320_ & ~new_n3388_;
  assign new_n3390_ = ~new_n3238_ & new_n3389_;
  assign new_n3391_ = ~new_n3384_ & ~new_n3390_;
  assign new_n3392_ = ~\b[3]  & ~new_n3391_;
  assign new_n3393_ = ~new_n3140_ & ~\quotient[44] ;
  assign new_n3394_ = ~new_n3143_ & new_n3145_;
  assign new_n3395_ = ~new_n3141_ & new_n3394_;
  assign new_n3396_ = new_n320_ & ~new_n3395_;
  assign new_n3397_ = ~new_n3146_ & new_n3396_;
  assign new_n3398_ = ~new_n3238_ & new_n3397_;
  assign new_n3399_ = ~new_n3393_ & ~new_n3398_;
  assign new_n3400_ = ~\b[2]  & ~new_n3399_;
  assign new_n3401_ = \b[0]  & ~\b[20] ;
  assign new_n3402_ = new_n366_ & new_n3401_;
  assign new_n3403_ = new_n377_ & new_n3402_;
  assign new_n3404_ = new_n423_ & new_n3403_;
  assign new_n3405_ = new_n408_ & new_n3404_;
  assign new_n3406_ = ~new_n3238_ & new_n3405_;
  assign new_n3407_ = \a[44]  & ~new_n3406_;
  assign new_n3408_ = new_n309_ & new_n3145_;
  assign new_n3409_ = new_n343_ & new_n3408_;
  assign new_n3410_ = new_n341_ & new_n3409_;
  assign new_n3411_ = new_n338_ & new_n3410_;
  assign new_n3412_ = ~new_n3238_ & new_n3411_;
  assign new_n3413_ = ~new_n3407_ & ~new_n3412_;
  assign new_n3414_ = \b[1]  & ~new_n3413_;
  assign new_n3415_ = ~\b[1]  & ~new_n3412_;
  assign new_n3416_ = ~new_n3407_ & new_n3415_;
  assign new_n3417_ = ~new_n3414_ & ~new_n3416_;
  assign new_n3418_ = ~\a[43]  & \b[0] ;
  assign new_n3419_ = ~new_n3417_ & ~new_n3418_;
  assign new_n3420_ = ~\b[1]  & ~new_n3413_;
  assign new_n3421_ = ~new_n3419_ & ~new_n3420_;
  assign new_n3422_ = \b[2]  & ~new_n3398_;
  assign new_n3423_ = ~new_n3393_ & new_n3422_;
  assign new_n3424_ = ~new_n3400_ & ~new_n3423_;
  assign new_n3425_ = ~new_n3421_ & new_n3424_;
  assign new_n3426_ = ~new_n3400_ & ~new_n3425_;
  assign new_n3427_ = \b[3]  & ~new_n3390_;
  assign new_n3428_ = ~new_n3384_ & new_n3427_;
  assign new_n3429_ = ~new_n3392_ & ~new_n3428_;
  assign new_n3430_ = ~new_n3426_ & new_n3429_;
  assign new_n3431_ = ~new_n3392_ & ~new_n3430_;
  assign new_n3432_ = \b[4]  & ~new_n3381_;
  assign new_n3433_ = ~new_n3375_ & new_n3432_;
  assign new_n3434_ = ~new_n3383_ & ~new_n3433_;
  assign new_n3435_ = ~new_n3431_ & new_n3434_;
  assign new_n3436_ = ~new_n3383_ & ~new_n3435_;
  assign new_n3437_ = \b[5]  & ~new_n3372_;
  assign new_n3438_ = ~new_n3366_ & new_n3437_;
  assign new_n3439_ = ~new_n3374_ & ~new_n3438_;
  assign new_n3440_ = ~new_n3436_ & new_n3439_;
  assign new_n3441_ = ~new_n3374_ & ~new_n3440_;
  assign new_n3442_ = \b[6]  & ~new_n3363_;
  assign new_n3443_ = ~new_n3357_ & new_n3442_;
  assign new_n3444_ = ~new_n3365_ & ~new_n3443_;
  assign new_n3445_ = ~new_n3441_ & new_n3444_;
  assign new_n3446_ = ~new_n3365_ & ~new_n3445_;
  assign new_n3447_ = \b[7]  & ~new_n3354_;
  assign new_n3448_ = ~new_n3348_ & new_n3447_;
  assign new_n3449_ = ~new_n3356_ & ~new_n3448_;
  assign new_n3450_ = ~new_n3446_ & new_n3449_;
  assign new_n3451_ = ~new_n3356_ & ~new_n3450_;
  assign new_n3452_ = \b[8]  & ~new_n3345_;
  assign new_n3453_ = ~new_n3339_ & new_n3452_;
  assign new_n3454_ = ~new_n3347_ & ~new_n3453_;
  assign new_n3455_ = ~new_n3451_ & new_n3454_;
  assign new_n3456_ = ~new_n3347_ & ~new_n3455_;
  assign new_n3457_ = \b[9]  & ~new_n3336_;
  assign new_n3458_ = ~new_n3330_ & new_n3457_;
  assign new_n3459_ = ~new_n3338_ & ~new_n3458_;
  assign new_n3460_ = ~new_n3456_ & new_n3459_;
  assign new_n3461_ = ~new_n3338_ & ~new_n3460_;
  assign new_n3462_ = \b[10]  & ~new_n3327_;
  assign new_n3463_ = ~new_n3321_ & new_n3462_;
  assign new_n3464_ = ~new_n3329_ & ~new_n3463_;
  assign new_n3465_ = ~new_n3461_ & new_n3464_;
  assign new_n3466_ = ~new_n3329_ & ~new_n3465_;
  assign new_n3467_ = \b[11]  & ~new_n3318_;
  assign new_n3468_ = ~new_n3312_ & new_n3467_;
  assign new_n3469_ = ~new_n3320_ & ~new_n3468_;
  assign new_n3470_ = ~new_n3466_ & new_n3469_;
  assign new_n3471_ = ~new_n3320_ & ~new_n3470_;
  assign new_n3472_ = \b[12]  & ~new_n3309_;
  assign new_n3473_ = ~new_n3303_ & new_n3472_;
  assign new_n3474_ = ~new_n3311_ & ~new_n3473_;
  assign new_n3475_ = ~new_n3471_ & new_n3474_;
  assign new_n3476_ = ~new_n3311_ & ~new_n3475_;
  assign new_n3477_ = \b[13]  & ~new_n3300_;
  assign new_n3478_ = ~new_n3294_ & new_n3477_;
  assign new_n3479_ = ~new_n3302_ & ~new_n3478_;
  assign new_n3480_ = ~new_n3476_ & new_n3479_;
  assign new_n3481_ = ~new_n3302_ & ~new_n3480_;
  assign new_n3482_ = \b[14]  & ~new_n3291_;
  assign new_n3483_ = ~new_n3285_ & new_n3482_;
  assign new_n3484_ = ~new_n3293_ & ~new_n3483_;
  assign new_n3485_ = ~new_n3481_ & new_n3484_;
  assign new_n3486_ = ~new_n3293_ & ~new_n3485_;
  assign new_n3487_ = \b[15]  & ~new_n3282_;
  assign new_n3488_ = ~new_n3276_ & new_n3487_;
  assign new_n3489_ = ~new_n3284_ & ~new_n3488_;
  assign new_n3490_ = ~new_n3486_ & new_n3489_;
  assign new_n3491_ = ~new_n3284_ & ~new_n3490_;
  assign new_n3492_ = \b[16]  & ~new_n3273_;
  assign new_n3493_ = ~new_n3267_ & new_n3492_;
  assign new_n3494_ = ~new_n3275_ & ~new_n3493_;
  assign new_n3495_ = ~new_n3491_ & new_n3494_;
  assign new_n3496_ = ~new_n3275_ & ~new_n3495_;
  assign new_n3497_ = \b[17]  & ~new_n3264_;
  assign new_n3498_ = ~new_n3258_ & new_n3497_;
  assign new_n3499_ = ~new_n3266_ & ~new_n3498_;
  assign new_n3500_ = ~new_n3496_ & new_n3499_;
  assign new_n3501_ = ~new_n3266_ & ~new_n3500_;
  assign new_n3502_ = \b[18]  & ~new_n3255_;
  assign new_n3503_ = ~new_n3249_ & new_n3502_;
  assign new_n3504_ = ~new_n3257_ & ~new_n3503_;
  assign new_n3505_ = ~new_n3501_ & new_n3504_;
  assign new_n3506_ = ~new_n3257_ & ~new_n3505_;
  assign new_n3507_ = \b[19]  & ~new_n3246_;
  assign new_n3508_ = ~new_n3240_ & new_n3507_;
  assign new_n3509_ = ~new_n3248_ & ~new_n3508_;
  assign new_n3510_ = ~new_n3506_ & new_n3509_;
  assign new_n3511_ = ~new_n3248_ & ~new_n3510_;
  assign new_n3512_ = ~new_n2981_ & ~\quotient[44] ;
  assign new_n3513_ = ~new_n2983_ & new_n3236_;
  assign new_n3514_ = ~new_n3232_ & new_n3513_;
  assign new_n3515_ = ~new_n3233_ & ~new_n3236_;
  assign new_n3516_ = ~new_n3514_ & ~new_n3515_;
  assign new_n3517_ = \quotient[44]  & ~new_n3516_;
  assign new_n3518_ = ~new_n3512_ & ~new_n3517_;
  assign new_n3519_ = ~\b[20]  & ~new_n3518_;
  assign new_n3520_ = \b[20]  & ~new_n3512_;
  assign new_n3521_ = ~new_n3517_ & new_n3520_;
  assign new_n3522_ = new_n643_ & ~new_n3521_;
  assign new_n3523_ = ~new_n3519_ & new_n3522_;
  assign new_n3524_ = ~new_n3511_ & new_n3523_;
  assign new_n3525_ = new_n320_ & ~new_n3518_;
  assign \quotient[43]  = new_n3524_ | new_n3525_;
  assign new_n3527_ = ~new_n3257_ & new_n3509_;
  assign new_n3528_ = ~new_n3505_ & new_n3527_;
  assign new_n3529_ = ~new_n3506_ & ~new_n3509_;
  assign new_n3530_ = ~new_n3528_ & ~new_n3529_;
  assign new_n3531_ = \quotient[43]  & ~new_n3530_;
  assign new_n3532_ = ~new_n3247_ & ~new_n3525_;
  assign new_n3533_ = ~new_n3524_ & new_n3532_;
  assign new_n3534_ = ~new_n3531_ & ~new_n3533_;
  assign new_n3535_ = ~new_n3248_ & ~new_n3521_;
  assign new_n3536_ = ~new_n3519_ & new_n3535_;
  assign new_n3537_ = ~new_n3510_ & new_n3536_;
  assign new_n3538_ = ~new_n3519_ & ~new_n3521_;
  assign new_n3539_ = ~new_n3511_ & ~new_n3538_;
  assign new_n3540_ = ~new_n3537_ & ~new_n3539_;
  assign new_n3541_ = \quotient[43]  & ~new_n3540_;
  assign new_n3542_ = ~new_n3518_ & ~new_n3525_;
  assign new_n3543_ = ~new_n3524_ & new_n3542_;
  assign new_n3544_ = ~new_n3541_ & ~new_n3543_;
  assign new_n3545_ = ~\b[21]  & ~new_n3544_;
  assign new_n3546_ = ~\b[20]  & ~new_n3534_;
  assign new_n3547_ = ~new_n3266_ & new_n3504_;
  assign new_n3548_ = ~new_n3500_ & new_n3547_;
  assign new_n3549_ = ~new_n3501_ & ~new_n3504_;
  assign new_n3550_ = ~new_n3548_ & ~new_n3549_;
  assign new_n3551_ = \quotient[43]  & ~new_n3550_;
  assign new_n3552_ = ~new_n3256_ & ~new_n3525_;
  assign new_n3553_ = ~new_n3524_ & new_n3552_;
  assign new_n3554_ = ~new_n3551_ & ~new_n3553_;
  assign new_n3555_ = ~\b[19]  & ~new_n3554_;
  assign new_n3556_ = ~new_n3275_ & new_n3499_;
  assign new_n3557_ = ~new_n3495_ & new_n3556_;
  assign new_n3558_ = ~new_n3496_ & ~new_n3499_;
  assign new_n3559_ = ~new_n3557_ & ~new_n3558_;
  assign new_n3560_ = \quotient[43]  & ~new_n3559_;
  assign new_n3561_ = ~new_n3265_ & ~new_n3525_;
  assign new_n3562_ = ~new_n3524_ & new_n3561_;
  assign new_n3563_ = ~new_n3560_ & ~new_n3562_;
  assign new_n3564_ = ~\b[18]  & ~new_n3563_;
  assign new_n3565_ = ~new_n3284_ & new_n3494_;
  assign new_n3566_ = ~new_n3490_ & new_n3565_;
  assign new_n3567_ = ~new_n3491_ & ~new_n3494_;
  assign new_n3568_ = ~new_n3566_ & ~new_n3567_;
  assign new_n3569_ = \quotient[43]  & ~new_n3568_;
  assign new_n3570_ = ~new_n3274_ & ~new_n3525_;
  assign new_n3571_ = ~new_n3524_ & new_n3570_;
  assign new_n3572_ = ~new_n3569_ & ~new_n3571_;
  assign new_n3573_ = ~\b[17]  & ~new_n3572_;
  assign new_n3574_ = ~new_n3293_ & new_n3489_;
  assign new_n3575_ = ~new_n3485_ & new_n3574_;
  assign new_n3576_ = ~new_n3486_ & ~new_n3489_;
  assign new_n3577_ = ~new_n3575_ & ~new_n3576_;
  assign new_n3578_ = \quotient[43]  & ~new_n3577_;
  assign new_n3579_ = ~new_n3283_ & ~new_n3525_;
  assign new_n3580_ = ~new_n3524_ & new_n3579_;
  assign new_n3581_ = ~new_n3578_ & ~new_n3580_;
  assign new_n3582_ = ~\b[16]  & ~new_n3581_;
  assign new_n3583_ = ~new_n3302_ & new_n3484_;
  assign new_n3584_ = ~new_n3480_ & new_n3583_;
  assign new_n3585_ = ~new_n3481_ & ~new_n3484_;
  assign new_n3586_ = ~new_n3584_ & ~new_n3585_;
  assign new_n3587_ = \quotient[43]  & ~new_n3586_;
  assign new_n3588_ = ~new_n3292_ & ~new_n3525_;
  assign new_n3589_ = ~new_n3524_ & new_n3588_;
  assign new_n3590_ = ~new_n3587_ & ~new_n3589_;
  assign new_n3591_ = ~\b[15]  & ~new_n3590_;
  assign new_n3592_ = ~new_n3311_ & new_n3479_;
  assign new_n3593_ = ~new_n3475_ & new_n3592_;
  assign new_n3594_ = ~new_n3476_ & ~new_n3479_;
  assign new_n3595_ = ~new_n3593_ & ~new_n3594_;
  assign new_n3596_ = \quotient[43]  & ~new_n3595_;
  assign new_n3597_ = ~new_n3301_ & ~new_n3525_;
  assign new_n3598_ = ~new_n3524_ & new_n3597_;
  assign new_n3599_ = ~new_n3596_ & ~new_n3598_;
  assign new_n3600_ = ~\b[14]  & ~new_n3599_;
  assign new_n3601_ = ~new_n3320_ & new_n3474_;
  assign new_n3602_ = ~new_n3470_ & new_n3601_;
  assign new_n3603_ = ~new_n3471_ & ~new_n3474_;
  assign new_n3604_ = ~new_n3602_ & ~new_n3603_;
  assign new_n3605_ = \quotient[43]  & ~new_n3604_;
  assign new_n3606_ = ~new_n3310_ & ~new_n3525_;
  assign new_n3607_ = ~new_n3524_ & new_n3606_;
  assign new_n3608_ = ~new_n3605_ & ~new_n3607_;
  assign new_n3609_ = ~\b[13]  & ~new_n3608_;
  assign new_n3610_ = ~new_n3329_ & new_n3469_;
  assign new_n3611_ = ~new_n3465_ & new_n3610_;
  assign new_n3612_ = ~new_n3466_ & ~new_n3469_;
  assign new_n3613_ = ~new_n3611_ & ~new_n3612_;
  assign new_n3614_ = \quotient[43]  & ~new_n3613_;
  assign new_n3615_ = ~new_n3319_ & ~new_n3525_;
  assign new_n3616_ = ~new_n3524_ & new_n3615_;
  assign new_n3617_ = ~new_n3614_ & ~new_n3616_;
  assign new_n3618_ = ~\b[12]  & ~new_n3617_;
  assign new_n3619_ = ~new_n3338_ & new_n3464_;
  assign new_n3620_ = ~new_n3460_ & new_n3619_;
  assign new_n3621_ = ~new_n3461_ & ~new_n3464_;
  assign new_n3622_ = ~new_n3620_ & ~new_n3621_;
  assign new_n3623_ = \quotient[43]  & ~new_n3622_;
  assign new_n3624_ = ~new_n3328_ & ~new_n3525_;
  assign new_n3625_ = ~new_n3524_ & new_n3624_;
  assign new_n3626_ = ~new_n3623_ & ~new_n3625_;
  assign new_n3627_ = ~\b[11]  & ~new_n3626_;
  assign new_n3628_ = ~new_n3347_ & new_n3459_;
  assign new_n3629_ = ~new_n3455_ & new_n3628_;
  assign new_n3630_ = ~new_n3456_ & ~new_n3459_;
  assign new_n3631_ = ~new_n3629_ & ~new_n3630_;
  assign new_n3632_ = \quotient[43]  & ~new_n3631_;
  assign new_n3633_ = ~new_n3337_ & ~new_n3525_;
  assign new_n3634_ = ~new_n3524_ & new_n3633_;
  assign new_n3635_ = ~new_n3632_ & ~new_n3634_;
  assign new_n3636_ = ~\b[10]  & ~new_n3635_;
  assign new_n3637_ = ~new_n3356_ & new_n3454_;
  assign new_n3638_ = ~new_n3450_ & new_n3637_;
  assign new_n3639_ = ~new_n3451_ & ~new_n3454_;
  assign new_n3640_ = ~new_n3638_ & ~new_n3639_;
  assign new_n3641_ = \quotient[43]  & ~new_n3640_;
  assign new_n3642_ = ~new_n3346_ & ~new_n3525_;
  assign new_n3643_ = ~new_n3524_ & new_n3642_;
  assign new_n3644_ = ~new_n3641_ & ~new_n3643_;
  assign new_n3645_ = ~\b[9]  & ~new_n3644_;
  assign new_n3646_ = ~new_n3365_ & new_n3449_;
  assign new_n3647_ = ~new_n3445_ & new_n3646_;
  assign new_n3648_ = ~new_n3446_ & ~new_n3449_;
  assign new_n3649_ = ~new_n3647_ & ~new_n3648_;
  assign new_n3650_ = \quotient[43]  & ~new_n3649_;
  assign new_n3651_ = ~new_n3355_ & ~new_n3525_;
  assign new_n3652_ = ~new_n3524_ & new_n3651_;
  assign new_n3653_ = ~new_n3650_ & ~new_n3652_;
  assign new_n3654_ = ~\b[8]  & ~new_n3653_;
  assign new_n3655_ = ~new_n3374_ & new_n3444_;
  assign new_n3656_ = ~new_n3440_ & new_n3655_;
  assign new_n3657_ = ~new_n3441_ & ~new_n3444_;
  assign new_n3658_ = ~new_n3656_ & ~new_n3657_;
  assign new_n3659_ = \quotient[43]  & ~new_n3658_;
  assign new_n3660_ = ~new_n3364_ & ~new_n3525_;
  assign new_n3661_ = ~new_n3524_ & new_n3660_;
  assign new_n3662_ = ~new_n3659_ & ~new_n3661_;
  assign new_n3663_ = ~\b[7]  & ~new_n3662_;
  assign new_n3664_ = ~new_n3383_ & new_n3439_;
  assign new_n3665_ = ~new_n3435_ & new_n3664_;
  assign new_n3666_ = ~new_n3436_ & ~new_n3439_;
  assign new_n3667_ = ~new_n3665_ & ~new_n3666_;
  assign new_n3668_ = \quotient[43]  & ~new_n3667_;
  assign new_n3669_ = ~new_n3373_ & ~new_n3525_;
  assign new_n3670_ = ~new_n3524_ & new_n3669_;
  assign new_n3671_ = ~new_n3668_ & ~new_n3670_;
  assign new_n3672_ = ~\b[6]  & ~new_n3671_;
  assign new_n3673_ = ~new_n3392_ & new_n3434_;
  assign new_n3674_ = ~new_n3430_ & new_n3673_;
  assign new_n3675_ = ~new_n3431_ & ~new_n3434_;
  assign new_n3676_ = ~new_n3674_ & ~new_n3675_;
  assign new_n3677_ = \quotient[43]  & ~new_n3676_;
  assign new_n3678_ = ~new_n3382_ & ~new_n3525_;
  assign new_n3679_ = ~new_n3524_ & new_n3678_;
  assign new_n3680_ = ~new_n3677_ & ~new_n3679_;
  assign new_n3681_ = ~\b[5]  & ~new_n3680_;
  assign new_n3682_ = ~new_n3400_ & new_n3429_;
  assign new_n3683_ = ~new_n3425_ & new_n3682_;
  assign new_n3684_ = ~new_n3426_ & ~new_n3429_;
  assign new_n3685_ = ~new_n3683_ & ~new_n3684_;
  assign new_n3686_ = \quotient[43]  & ~new_n3685_;
  assign new_n3687_ = ~new_n3391_ & ~new_n3525_;
  assign new_n3688_ = ~new_n3524_ & new_n3687_;
  assign new_n3689_ = ~new_n3686_ & ~new_n3688_;
  assign new_n3690_ = ~\b[4]  & ~new_n3689_;
  assign new_n3691_ = ~new_n3420_ & new_n3424_;
  assign new_n3692_ = ~new_n3419_ & new_n3691_;
  assign new_n3693_ = ~new_n3421_ & ~new_n3424_;
  assign new_n3694_ = ~new_n3692_ & ~new_n3693_;
  assign new_n3695_ = \quotient[43]  & ~new_n3694_;
  assign new_n3696_ = ~new_n3399_ & ~new_n3525_;
  assign new_n3697_ = ~new_n3524_ & new_n3696_;
  assign new_n3698_ = ~new_n3695_ & ~new_n3697_;
  assign new_n3699_ = ~\b[3]  & ~new_n3698_;
  assign new_n3700_ = ~new_n3416_ & new_n3418_;
  assign new_n3701_ = ~new_n3414_ & new_n3700_;
  assign new_n3702_ = ~new_n3419_ & ~new_n3701_;
  assign new_n3703_ = \quotient[43]  & new_n3702_;
  assign new_n3704_ = ~new_n3413_ & ~new_n3525_;
  assign new_n3705_ = ~new_n3524_ & new_n3704_;
  assign new_n3706_ = ~new_n3703_ & ~new_n3705_;
  assign new_n3707_ = ~\b[2]  & ~new_n3706_;
  assign new_n3708_ = \b[0]  & \quotient[43] ;
  assign new_n3709_ = \a[43]  & ~new_n3708_;
  assign new_n3710_ = new_n3418_ & \quotient[43] ;
  assign new_n3711_ = ~new_n3709_ & ~new_n3710_;
  assign new_n3712_ = \b[1]  & ~new_n3711_;
  assign new_n3713_ = ~\b[1]  & ~new_n3710_;
  assign new_n3714_ = ~new_n3709_ & new_n3713_;
  assign new_n3715_ = ~new_n3712_ & ~new_n3714_;
  assign new_n3716_ = ~\a[42]  & \b[0] ;
  assign new_n3717_ = ~new_n3715_ & ~new_n3716_;
  assign new_n3718_ = ~\b[1]  & ~new_n3711_;
  assign new_n3719_ = ~new_n3717_ & ~new_n3718_;
  assign new_n3720_ = \b[2]  & ~new_n3705_;
  assign new_n3721_ = ~new_n3703_ & new_n3720_;
  assign new_n3722_ = ~new_n3707_ & ~new_n3721_;
  assign new_n3723_ = ~new_n3719_ & new_n3722_;
  assign new_n3724_ = ~new_n3707_ & ~new_n3723_;
  assign new_n3725_ = \b[3]  & ~new_n3697_;
  assign new_n3726_ = ~new_n3695_ & new_n3725_;
  assign new_n3727_ = ~new_n3699_ & ~new_n3726_;
  assign new_n3728_ = ~new_n3724_ & new_n3727_;
  assign new_n3729_ = ~new_n3699_ & ~new_n3728_;
  assign new_n3730_ = \b[4]  & ~new_n3688_;
  assign new_n3731_ = ~new_n3686_ & new_n3730_;
  assign new_n3732_ = ~new_n3690_ & ~new_n3731_;
  assign new_n3733_ = ~new_n3729_ & new_n3732_;
  assign new_n3734_ = ~new_n3690_ & ~new_n3733_;
  assign new_n3735_ = \b[5]  & ~new_n3679_;
  assign new_n3736_ = ~new_n3677_ & new_n3735_;
  assign new_n3737_ = ~new_n3681_ & ~new_n3736_;
  assign new_n3738_ = ~new_n3734_ & new_n3737_;
  assign new_n3739_ = ~new_n3681_ & ~new_n3738_;
  assign new_n3740_ = \b[6]  & ~new_n3670_;
  assign new_n3741_ = ~new_n3668_ & new_n3740_;
  assign new_n3742_ = ~new_n3672_ & ~new_n3741_;
  assign new_n3743_ = ~new_n3739_ & new_n3742_;
  assign new_n3744_ = ~new_n3672_ & ~new_n3743_;
  assign new_n3745_ = \b[7]  & ~new_n3661_;
  assign new_n3746_ = ~new_n3659_ & new_n3745_;
  assign new_n3747_ = ~new_n3663_ & ~new_n3746_;
  assign new_n3748_ = ~new_n3744_ & new_n3747_;
  assign new_n3749_ = ~new_n3663_ & ~new_n3748_;
  assign new_n3750_ = \b[8]  & ~new_n3652_;
  assign new_n3751_ = ~new_n3650_ & new_n3750_;
  assign new_n3752_ = ~new_n3654_ & ~new_n3751_;
  assign new_n3753_ = ~new_n3749_ & new_n3752_;
  assign new_n3754_ = ~new_n3654_ & ~new_n3753_;
  assign new_n3755_ = \b[9]  & ~new_n3643_;
  assign new_n3756_ = ~new_n3641_ & new_n3755_;
  assign new_n3757_ = ~new_n3645_ & ~new_n3756_;
  assign new_n3758_ = ~new_n3754_ & new_n3757_;
  assign new_n3759_ = ~new_n3645_ & ~new_n3758_;
  assign new_n3760_ = \b[10]  & ~new_n3634_;
  assign new_n3761_ = ~new_n3632_ & new_n3760_;
  assign new_n3762_ = ~new_n3636_ & ~new_n3761_;
  assign new_n3763_ = ~new_n3759_ & new_n3762_;
  assign new_n3764_ = ~new_n3636_ & ~new_n3763_;
  assign new_n3765_ = \b[11]  & ~new_n3625_;
  assign new_n3766_ = ~new_n3623_ & new_n3765_;
  assign new_n3767_ = ~new_n3627_ & ~new_n3766_;
  assign new_n3768_ = ~new_n3764_ & new_n3767_;
  assign new_n3769_ = ~new_n3627_ & ~new_n3768_;
  assign new_n3770_ = \b[12]  & ~new_n3616_;
  assign new_n3771_ = ~new_n3614_ & new_n3770_;
  assign new_n3772_ = ~new_n3618_ & ~new_n3771_;
  assign new_n3773_ = ~new_n3769_ & new_n3772_;
  assign new_n3774_ = ~new_n3618_ & ~new_n3773_;
  assign new_n3775_ = \b[13]  & ~new_n3607_;
  assign new_n3776_ = ~new_n3605_ & new_n3775_;
  assign new_n3777_ = ~new_n3609_ & ~new_n3776_;
  assign new_n3778_ = ~new_n3774_ & new_n3777_;
  assign new_n3779_ = ~new_n3609_ & ~new_n3778_;
  assign new_n3780_ = \b[14]  & ~new_n3598_;
  assign new_n3781_ = ~new_n3596_ & new_n3780_;
  assign new_n3782_ = ~new_n3600_ & ~new_n3781_;
  assign new_n3783_ = ~new_n3779_ & new_n3782_;
  assign new_n3784_ = ~new_n3600_ & ~new_n3783_;
  assign new_n3785_ = \b[15]  & ~new_n3589_;
  assign new_n3786_ = ~new_n3587_ & new_n3785_;
  assign new_n3787_ = ~new_n3591_ & ~new_n3786_;
  assign new_n3788_ = ~new_n3784_ & new_n3787_;
  assign new_n3789_ = ~new_n3591_ & ~new_n3788_;
  assign new_n3790_ = \b[16]  & ~new_n3580_;
  assign new_n3791_ = ~new_n3578_ & new_n3790_;
  assign new_n3792_ = ~new_n3582_ & ~new_n3791_;
  assign new_n3793_ = ~new_n3789_ & new_n3792_;
  assign new_n3794_ = ~new_n3582_ & ~new_n3793_;
  assign new_n3795_ = \b[17]  & ~new_n3571_;
  assign new_n3796_ = ~new_n3569_ & new_n3795_;
  assign new_n3797_ = ~new_n3573_ & ~new_n3796_;
  assign new_n3798_ = ~new_n3794_ & new_n3797_;
  assign new_n3799_ = ~new_n3573_ & ~new_n3798_;
  assign new_n3800_ = \b[18]  & ~new_n3562_;
  assign new_n3801_ = ~new_n3560_ & new_n3800_;
  assign new_n3802_ = ~new_n3564_ & ~new_n3801_;
  assign new_n3803_ = ~new_n3799_ & new_n3802_;
  assign new_n3804_ = ~new_n3564_ & ~new_n3803_;
  assign new_n3805_ = \b[19]  & ~new_n3553_;
  assign new_n3806_ = ~new_n3551_ & new_n3805_;
  assign new_n3807_ = ~new_n3555_ & ~new_n3806_;
  assign new_n3808_ = ~new_n3804_ & new_n3807_;
  assign new_n3809_ = ~new_n3555_ & ~new_n3808_;
  assign new_n3810_ = \b[20]  & ~new_n3533_;
  assign new_n3811_ = ~new_n3531_ & new_n3810_;
  assign new_n3812_ = ~new_n3546_ & ~new_n3811_;
  assign new_n3813_ = ~new_n3809_ & new_n3812_;
  assign new_n3814_ = ~new_n3546_ & ~new_n3813_;
  assign new_n3815_ = \b[21]  & ~new_n3543_;
  assign new_n3816_ = ~new_n3541_ & new_n3815_;
  assign new_n3817_ = ~new_n3545_ & ~new_n3816_;
  assign new_n3818_ = ~new_n3814_ & new_n3817_;
  assign new_n3819_ = ~new_n3545_ & ~new_n3818_;
  assign new_n3820_ = new_n306_ & new_n308_;
  assign new_n3821_ = new_n317_ & new_n3820_;
  assign new_n3822_ = new_n303_ & new_n3821_;
  assign new_n3823_ = new_n288_ & new_n3822_;
  assign \quotient[42]  = ~new_n3819_ & new_n3823_;
  assign new_n3825_ = ~new_n3534_ & ~\quotient[42] ;
  assign new_n3826_ = ~new_n3555_ & new_n3812_;
  assign new_n3827_ = ~new_n3808_ & new_n3826_;
  assign new_n3828_ = ~new_n3809_ & ~new_n3812_;
  assign new_n3829_ = ~new_n3827_ & ~new_n3828_;
  assign new_n3830_ = new_n3823_ & ~new_n3829_;
  assign new_n3831_ = ~new_n3819_ & new_n3830_;
  assign new_n3832_ = ~new_n3825_ & ~new_n3831_;
  assign new_n3833_ = ~new_n3544_ & ~\quotient[42] ;
  assign new_n3834_ = ~new_n3546_ & new_n3817_;
  assign new_n3835_ = ~new_n3813_ & new_n3834_;
  assign new_n3836_ = ~new_n3814_ & ~new_n3817_;
  assign new_n3837_ = ~new_n3835_ & ~new_n3836_;
  assign new_n3838_ = \quotient[42]  & ~new_n3837_;
  assign new_n3839_ = ~new_n3833_ & ~new_n3838_;
  assign new_n3840_ = ~\b[22]  & ~new_n3839_;
  assign new_n3841_ = ~\b[21]  & ~new_n3832_;
  assign new_n3842_ = ~new_n3554_ & ~\quotient[42] ;
  assign new_n3843_ = ~new_n3564_ & new_n3807_;
  assign new_n3844_ = ~new_n3803_ & new_n3843_;
  assign new_n3845_ = ~new_n3804_ & ~new_n3807_;
  assign new_n3846_ = ~new_n3844_ & ~new_n3845_;
  assign new_n3847_ = new_n3823_ & ~new_n3846_;
  assign new_n3848_ = ~new_n3819_ & new_n3847_;
  assign new_n3849_ = ~new_n3842_ & ~new_n3848_;
  assign new_n3850_ = ~\b[20]  & ~new_n3849_;
  assign new_n3851_ = ~new_n3563_ & ~\quotient[42] ;
  assign new_n3852_ = ~new_n3573_ & new_n3802_;
  assign new_n3853_ = ~new_n3798_ & new_n3852_;
  assign new_n3854_ = ~new_n3799_ & ~new_n3802_;
  assign new_n3855_ = ~new_n3853_ & ~new_n3854_;
  assign new_n3856_ = new_n3823_ & ~new_n3855_;
  assign new_n3857_ = ~new_n3819_ & new_n3856_;
  assign new_n3858_ = ~new_n3851_ & ~new_n3857_;
  assign new_n3859_ = ~\b[19]  & ~new_n3858_;
  assign new_n3860_ = ~new_n3572_ & ~\quotient[42] ;
  assign new_n3861_ = ~new_n3582_ & new_n3797_;
  assign new_n3862_ = ~new_n3793_ & new_n3861_;
  assign new_n3863_ = ~new_n3794_ & ~new_n3797_;
  assign new_n3864_ = ~new_n3862_ & ~new_n3863_;
  assign new_n3865_ = new_n3823_ & ~new_n3864_;
  assign new_n3866_ = ~new_n3819_ & new_n3865_;
  assign new_n3867_ = ~new_n3860_ & ~new_n3866_;
  assign new_n3868_ = ~\b[18]  & ~new_n3867_;
  assign new_n3869_ = ~new_n3581_ & ~\quotient[42] ;
  assign new_n3870_ = ~new_n3591_ & new_n3792_;
  assign new_n3871_ = ~new_n3788_ & new_n3870_;
  assign new_n3872_ = ~new_n3789_ & ~new_n3792_;
  assign new_n3873_ = ~new_n3871_ & ~new_n3872_;
  assign new_n3874_ = new_n3823_ & ~new_n3873_;
  assign new_n3875_ = ~new_n3819_ & new_n3874_;
  assign new_n3876_ = ~new_n3869_ & ~new_n3875_;
  assign new_n3877_ = ~\b[17]  & ~new_n3876_;
  assign new_n3878_ = ~new_n3590_ & ~\quotient[42] ;
  assign new_n3879_ = ~new_n3600_ & new_n3787_;
  assign new_n3880_ = ~new_n3783_ & new_n3879_;
  assign new_n3881_ = ~new_n3784_ & ~new_n3787_;
  assign new_n3882_ = ~new_n3880_ & ~new_n3881_;
  assign new_n3883_ = new_n3823_ & ~new_n3882_;
  assign new_n3884_ = ~new_n3819_ & new_n3883_;
  assign new_n3885_ = ~new_n3878_ & ~new_n3884_;
  assign new_n3886_ = ~\b[16]  & ~new_n3885_;
  assign new_n3887_ = ~new_n3599_ & ~\quotient[42] ;
  assign new_n3888_ = ~new_n3609_ & new_n3782_;
  assign new_n3889_ = ~new_n3778_ & new_n3888_;
  assign new_n3890_ = ~new_n3779_ & ~new_n3782_;
  assign new_n3891_ = ~new_n3889_ & ~new_n3890_;
  assign new_n3892_ = new_n3823_ & ~new_n3891_;
  assign new_n3893_ = ~new_n3819_ & new_n3892_;
  assign new_n3894_ = ~new_n3887_ & ~new_n3893_;
  assign new_n3895_ = ~\b[15]  & ~new_n3894_;
  assign new_n3896_ = ~new_n3608_ & ~\quotient[42] ;
  assign new_n3897_ = ~new_n3618_ & new_n3777_;
  assign new_n3898_ = ~new_n3773_ & new_n3897_;
  assign new_n3899_ = ~new_n3774_ & ~new_n3777_;
  assign new_n3900_ = ~new_n3898_ & ~new_n3899_;
  assign new_n3901_ = new_n3823_ & ~new_n3900_;
  assign new_n3902_ = ~new_n3819_ & new_n3901_;
  assign new_n3903_ = ~new_n3896_ & ~new_n3902_;
  assign new_n3904_ = ~\b[14]  & ~new_n3903_;
  assign new_n3905_ = ~new_n3617_ & ~\quotient[42] ;
  assign new_n3906_ = ~new_n3627_ & new_n3772_;
  assign new_n3907_ = ~new_n3768_ & new_n3906_;
  assign new_n3908_ = ~new_n3769_ & ~new_n3772_;
  assign new_n3909_ = ~new_n3907_ & ~new_n3908_;
  assign new_n3910_ = new_n3823_ & ~new_n3909_;
  assign new_n3911_ = ~new_n3819_ & new_n3910_;
  assign new_n3912_ = ~new_n3905_ & ~new_n3911_;
  assign new_n3913_ = ~\b[13]  & ~new_n3912_;
  assign new_n3914_ = ~new_n3626_ & ~\quotient[42] ;
  assign new_n3915_ = ~new_n3636_ & new_n3767_;
  assign new_n3916_ = ~new_n3763_ & new_n3915_;
  assign new_n3917_ = ~new_n3764_ & ~new_n3767_;
  assign new_n3918_ = ~new_n3916_ & ~new_n3917_;
  assign new_n3919_ = new_n3823_ & ~new_n3918_;
  assign new_n3920_ = ~new_n3819_ & new_n3919_;
  assign new_n3921_ = ~new_n3914_ & ~new_n3920_;
  assign new_n3922_ = ~\b[12]  & ~new_n3921_;
  assign new_n3923_ = ~new_n3635_ & ~\quotient[42] ;
  assign new_n3924_ = ~new_n3645_ & new_n3762_;
  assign new_n3925_ = ~new_n3758_ & new_n3924_;
  assign new_n3926_ = ~new_n3759_ & ~new_n3762_;
  assign new_n3927_ = ~new_n3925_ & ~new_n3926_;
  assign new_n3928_ = new_n3823_ & ~new_n3927_;
  assign new_n3929_ = ~new_n3819_ & new_n3928_;
  assign new_n3930_ = ~new_n3923_ & ~new_n3929_;
  assign new_n3931_ = ~\b[11]  & ~new_n3930_;
  assign new_n3932_ = ~new_n3644_ & ~\quotient[42] ;
  assign new_n3933_ = ~new_n3654_ & new_n3757_;
  assign new_n3934_ = ~new_n3753_ & new_n3933_;
  assign new_n3935_ = ~new_n3754_ & ~new_n3757_;
  assign new_n3936_ = ~new_n3934_ & ~new_n3935_;
  assign new_n3937_ = new_n3823_ & ~new_n3936_;
  assign new_n3938_ = ~new_n3819_ & new_n3937_;
  assign new_n3939_ = ~new_n3932_ & ~new_n3938_;
  assign new_n3940_ = ~\b[10]  & ~new_n3939_;
  assign new_n3941_ = ~new_n3653_ & ~\quotient[42] ;
  assign new_n3942_ = ~new_n3663_ & new_n3752_;
  assign new_n3943_ = ~new_n3748_ & new_n3942_;
  assign new_n3944_ = ~new_n3749_ & ~new_n3752_;
  assign new_n3945_ = ~new_n3943_ & ~new_n3944_;
  assign new_n3946_ = new_n3823_ & ~new_n3945_;
  assign new_n3947_ = ~new_n3819_ & new_n3946_;
  assign new_n3948_ = ~new_n3941_ & ~new_n3947_;
  assign new_n3949_ = ~\b[9]  & ~new_n3948_;
  assign new_n3950_ = ~new_n3662_ & ~\quotient[42] ;
  assign new_n3951_ = ~new_n3672_ & new_n3747_;
  assign new_n3952_ = ~new_n3743_ & new_n3951_;
  assign new_n3953_ = ~new_n3744_ & ~new_n3747_;
  assign new_n3954_ = ~new_n3952_ & ~new_n3953_;
  assign new_n3955_ = new_n3823_ & ~new_n3954_;
  assign new_n3956_ = ~new_n3819_ & new_n3955_;
  assign new_n3957_ = ~new_n3950_ & ~new_n3956_;
  assign new_n3958_ = ~\b[8]  & ~new_n3957_;
  assign new_n3959_ = ~new_n3671_ & ~\quotient[42] ;
  assign new_n3960_ = ~new_n3681_ & new_n3742_;
  assign new_n3961_ = ~new_n3738_ & new_n3960_;
  assign new_n3962_ = ~new_n3739_ & ~new_n3742_;
  assign new_n3963_ = ~new_n3961_ & ~new_n3962_;
  assign new_n3964_ = new_n3823_ & ~new_n3963_;
  assign new_n3965_ = ~new_n3819_ & new_n3964_;
  assign new_n3966_ = ~new_n3959_ & ~new_n3965_;
  assign new_n3967_ = ~\b[7]  & ~new_n3966_;
  assign new_n3968_ = ~new_n3680_ & ~\quotient[42] ;
  assign new_n3969_ = ~new_n3690_ & new_n3737_;
  assign new_n3970_ = ~new_n3733_ & new_n3969_;
  assign new_n3971_ = ~new_n3734_ & ~new_n3737_;
  assign new_n3972_ = ~new_n3970_ & ~new_n3971_;
  assign new_n3973_ = new_n3823_ & ~new_n3972_;
  assign new_n3974_ = ~new_n3819_ & new_n3973_;
  assign new_n3975_ = ~new_n3968_ & ~new_n3974_;
  assign new_n3976_ = ~\b[6]  & ~new_n3975_;
  assign new_n3977_ = ~new_n3689_ & ~\quotient[42] ;
  assign new_n3978_ = ~new_n3699_ & new_n3732_;
  assign new_n3979_ = ~new_n3728_ & new_n3978_;
  assign new_n3980_ = ~new_n3729_ & ~new_n3732_;
  assign new_n3981_ = ~new_n3979_ & ~new_n3980_;
  assign new_n3982_ = new_n3823_ & ~new_n3981_;
  assign new_n3983_ = ~new_n3819_ & new_n3982_;
  assign new_n3984_ = ~new_n3977_ & ~new_n3983_;
  assign new_n3985_ = ~\b[5]  & ~new_n3984_;
  assign new_n3986_ = ~new_n3698_ & ~\quotient[42] ;
  assign new_n3987_ = ~new_n3707_ & new_n3727_;
  assign new_n3988_ = ~new_n3723_ & new_n3987_;
  assign new_n3989_ = ~new_n3724_ & ~new_n3727_;
  assign new_n3990_ = ~new_n3988_ & ~new_n3989_;
  assign new_n3991_ = new_n3823_ & ~new_n3990_;
  assign new_n3992_ = ~new_n3819_ & new_n3991_;
  assign new_n3993_ = ~new_n3986_ & ~new_n3992_;
  assign new_n3994_ = ~\b[4]  & ~new_n3993_;
  assign new_n3995_ = ~new_n3706_ & ~\quotient[42] ;
  assign new_n3996_ = ~new_n3718_ & new_n3722_;
  assign new_n3997_ = ~new_n3717_ & new_n3996_;
  assign new_n3998_ = ~new_n3719_ & ~new_n3722_;
  assign new_n3999_ = ~new_n3997_ & ~new_n3998_;
  assign new_n4000_ = new_n3823_ & ~new_n3999_;
  assign new_n4001_ = ~new_n3819_ & new_n4000_;
  assign new_n4002_ = ~new_n3995_ & ~new_n4001_;
  assign new_n4003_ = ~\b[3]  & ~new_n4002_;
  assign new_n4004_ = ~new_n3711_ & ~\quotient[42] ;
  assign new_n4005_ = ~new_n3714_ & new_n3716_;
  assign new_n4006_ = ~new_n3712_ & new_n4005_;
  assign new_n4007_ = new_n3823_ & ~new_n4006_;
  assign new_n4008_ = ~new_n3717_ & new_n4007_;
  assign new_n4009_ = ~new_n3819_ & new_n4008_;
  assign new_n4010_ = ~new_n4004_ & ~new_n4009_;
  assign new_n4011_ = ~\b[2]  & ~new_n4010_;
  assign new_n4012_ = \b[0]  & ~\b[22] ;
  assign new_n4013_ = new_n365_ & new_n4012_;
  assign new_n4014_ = new_n376_ & new_n4013_;
  assign new_n4015_ = new_n588_ & new_n4014_;
  assign new_n4016_ = new_n598_ & new_n4015_;
  assign new_n4017_ = new_n595_ & new_n4016_;
  assign new_n4018_ = ~new_n3819_ & new_n4017_;
  assign new_n4019_ = \a[42]  & ~new_n4018_;
  assign new_n4020_ = new_n308_ & new_n3716_;
  assign new_n4021_ = new_n306_ & new_n4020_;
  assign new_n4022_ = new_n317_ & new_n4021_;
  assign new_n4023_ = new_n303_ & new_n4022_;
  assign new_n4024_ = new_n288_ & new_n4023_;
  assign new_n4025_ = ~new_n3819_ & new_n4024_;
  assign new_n4026_ = ~new_n4019_ & ~new_n4025_;
  assign new_n4027_ = \b[1]  & ~new_n4026_;
  assign new_n4028_ = ~\b[1]  & ~new_n4025_;
  assign new_n4029_ = ~new_n4019_ & new_n4028_;
  assign new_n4030_ = ~new_n4027_ & ~new_n4029_;
  assign new_n4031_ = ~\a[41]  & \b[0] ;
  assign new_n4032_ = ~new_n4030_ & ~new_n4031_;
  assign new_n4033_ = ~\b[1]  & ~new_n4026_;
  assign new_n4034_ = ~new_n4032_ & ~new_n4033_;
  assign new_n4035_ = \b[2]  & ~new_n4009_;
  assign new_n4036_ = ~new_n4004_ & new_n4035_;
  assign new_n4037_ = ~new_n4011_ & ~new_n4036_;
  assign new_n4038_ = ~new_n4034_ & new_n4037_;
  assign new_n4039_ = ~new_n4011_ & ~new_n4038_;
  assign new_n4040_ = \b[3]  & ~new_n4001_;
  assign new_n4041_ = ~new_n3995_ & new_n4040_;
  assign new_n4042_ = ~new_n4003_ & ~new_n4041_;
  assign new_n4043_ = ~new_n4039_ & new_n4042_;
  assign new_n4044_ = ~new_n4003_ & ~new_n4043_;
  assign new_n4045_ = \b[4]  & ~new_n3992_;
  assign new_n4046_ = ~new_n3986_ & new_n4045_;
  assign new_n4047_ = ~new_n3994_ & ~new_n4046_;
  assign new_n4048_ = ~new_n4044_ & new_n4047_;
  assign new_n4049_ = ~new_n3994_ & ~new_n4048_;
  assign new_n4050_ = \b[5]  & ~new_n3983_;
  assign new_n4051_ = ~new_n3977_ & new_n4050_;
  assign new_n4052_ = ~new_n3985_ & ~new_n4051_;
  assign new_n4053_ = ~new_n4049_ & new_n4052_;
  assign new_n4054_ = ~new_n3985_ & ~new_n4053_;
  assign new_n4055_ = \b[6]  & ~new_n3974_;
  assign new_n4056_ = ~new_n3968_ & new_n4055_;
  assign new_n4057_ = ~new_n3976_ & ~new_n4056_;
  assign new_n4058_ = ~new_n4054_ & new_n4057_;
  assign new_n4059_ = ~new_n3976_ & ~new_n4058_;
  assign new_n4060_ = \b[7]  & ~new_n3965_;
  assign new_n4061_ = ~new_n3959_ & new_n4060_;
  assign new_n4062_ = ~new_n3967_ & ~new_n4061_;
  assign new_n4063_ = ~new_n4059_ & new_n4062_;
  assign new_n4064_ = ~new_n3967_ & ~new_n4063_;
  assign new_n4065_ = \b[8]  & ~new_n3956_;
  assign new_n4066_ = ~new_n3950_ & new_n4065_;
  assign new_n4067_ = ~new_n3958_ & ~new_n4066_;
  assign new_n4068_ = ~new_n4064_ & new_n4067_;
  assign new_n4069_ = ~new_n3958_ & ~new_n4068_;
  assign new_n4070_ = \b[9]  & ~new_n3947_;
  assign new_n4071_ = ~new_n3941_ & new_n4070_;
  assign new_n4072_ = ~new_n3949_ & ~new_n4071_;
  assign new_n4073_ = ~new_n4069_ & new_n4072_;
  assign new_n4074_ = ~new_n3949_ & ~new_n4073_;
  assign new_n4075_ = \b[10]  & ~new_n3938_;
  assign new_n4076_ = ~new_n3932_ & new_n4075_;
  assign new_n4077_ = ~new_n3940_ & ~new_n4076_;
  assign new_n4078_ = ~new_n4074_ & new_n4077_;
  assign new_n4079_ = ~new_n3940_ & ~new_n4078_;
  assign new_n4080_ = \b[11]  & ~new_n3929_;
  assign new_n4081_ = ~new_n3923_ & new_n4080_;
  assign new_n4082_ = ~new_n3931_ & ~new_n4081_;
  assign new_n4083_ = ~new_n4079_ & new_n4082_;
  assign new_n4084_ = ~new_n3931_ & ~new_n4083_;
  assign new_n4085_ = \b[12]  & ~new_n3920_;
  assign new_n4086_ = ~new_n3914_ & new_n4085_;
  assign new_n4087_ = ~new_n3922_ & ~new_n4086_;
  assign new_n4088_ = ~new_n4084_ & new_n4087_;
  assign new_n4089_ = ~new_n3922_ & ~new_n4088_;
  assign new_n4090_ = \b[13]  & ~new_n3911_;
  assign new_n4091_ = ~new_n3905_ & new_n4090_;
  assign new_n4092_ = ~new_n3913_ & ~new_n4091_;
  assign new_n4093_ = ~new_n4089_ & new_n4092_;
  assign new_n4094_ = ~new_n3913_ & ~new_n4093_;
  assign new_n4095_ = \b[14]  & ~new_n3902_;
  assign new_n4096_ = ~new_n3896_ & new_n4095_;
  assign new_n4097_ = ~new_n3904_ & ~new_n4096_;
  assign new_n4098_ = ~new_n4094_ & new_n4097_;
  assign new_n4099_ = ~new_n3904_ & ~new_n4098_;
  assign new_n4100_ = \b[15]  & ~new_n3893_;
  assign new_n4101_ = ~new_n3887_ & new_n4100_;
  assign new_n4102_ = ~new_n3895_ & ~new_n4101_;
  assign new_n4103_ = ~new_n4099_ & new_n4102_;
  assign new_n4104_ = ~new_n3895_ & ~new_n4103_;
  assign new_n4105_ = \b[16]  & ~new_n3884_;
  assign new_n4106_ = ~new_n3878_ & new_n4105_;
  assign new_n4107_ = ~new_n3886_ & ~new_n4106_;
  assign new_n4108_ = ~new_n4104_ & new_n4107_;
  assign new_n4109_ = ~new_n3886_ & ~new_n4108_;
  assign new_n4110_ = \b[17]  & ~new_n3875_;
  assign new_n4111_ = ~new_n3869_ & new_n4110_;
  assign new_n4112_ = ~new_n3877_ & ~new_n4111_;
  assign new_n4113_ = ~new_n4109_ & new_n4112_;
  assign new_n4114_ = ~new_n3877_ & ~new_n4113_;
  assign new_n4115_ = \b[18]  & ~new_n3866_;
  assign new_n4116_ = ~new_n3860_ & new_n4115_;
  assign new_n4117_ = ~new_n3868_ & ~new_n4116_;
  assign new_n4118_ = ~new_n4114_ & new_n4117_;
  assign new_n4119_ = ~new_n3868_ & ~new_n4118_;
  assign new_n4120_ = \b[19]  & ~new_n3857_;
  assign new_n4121_ = ~new_n3851_ & new_n4120_;
  assign new_n4122_ = ~new_n3859_ & ~new_n4121_;
  assign new_n4123_ = ~new_n4119_ & new_n4122_;
  assign new_n4124_ = ~new_n3859_ & ~new_n4123_;
  assign new_n4125_ = \b[20]  & ~new_n3848_;
  assign new_n4126_ = ~new_n3842_ & new_n4125_;
  assign new_n4127_ = ~new_n3850_ & ~new_n4126_;
  assign new_n4128_ = ~new_n4124_ & new_n4127_;
  assign new_n4129_ = ~new_n3850_ & ~new_n4128_;
  assign new_n4130_ = \b[21]  & ~new_n3831_;
  assign new_n4131_ = ~new_n3825_ & new_n4130_;
  assign new_n4132_ = ~new_n3841_ & ~new_n4131_;
  assign new_n4133_ = ~new_n4129_ & new_n4132_;
  assign new_n4134_ = ~new_n3841_ & ~new_n4133_;
  assign new_n4135_ = \b[22]  & ~new_n3833_;
  assign new_n4136_ = ~new_n3838_ & new_n4135_;
  assign new_n4137_ = ~new_n3840_ & ~new_n4136_;
  assign new_n4138_ = ~new_n4134_ & new_n4137_;
  assign new_n4139_ = ~new_n3840_ & ~new_n4138_;
  assign new_n4140_ = new_n365_ & new_n376_;
  assign new_n4141_ = new_n588_ & new_n4140_;
  assign new_n4142_ = new_n598_ & new_n4141_;
  assign new_n4143_ = new_n595_ & new_n4142_;
  assign \quotient[41]  = ~new_n4139_ & new_n4143_;
  assign new_n4145_ = ~new_n3832_ & ~\quotient[41] ;
  assign new_n4146_ = ~new_n3850_ & new_n4132_;
  assign new_n4147_ = ~new_n4128_ & new_n4146_;
  assign new_n4148_ = ~new_n4129_ & ~new_n4132_;
  assign new_n4149_ = ~new_n4147_ & ~new_n4148_;
  assign new_n4150_ = new_n4143_ & ~new_n4149_;
  assign new_n4151_ = ~new_n4139_ & new_n4150_;
  assign new_n4152_ = ~new_n4145_ & ~new_n4151_;
  assign new_n4153_ = ~\b[22]  & ~new_n4152_;
  assign new_n4154_ = ~new_n3849_ & ~\quotient[41] ;
  assign new_n4155_ = ~new_n3859_ & new_n4127_;
  assign new_n4156_ = ~new_n4123_ & new_n4155_;
  assign new_n4157_ = ~new_n4124_ & ~new_n4127_;
  assign new_n4158_ = ~new_n4156_ & ~new_n4157_;
  assign new_n4159_ = new_n4143_ & ~new_n4158_;
  assign new_n4160_ = ~new_n4139_ & new_n4159_;
  assign new_n4161_ = ~new_n4154_ & ~new_n4160_;
  assign new_n4162_ = ~\b[21]  & ~new_n4161_;
  assign new_n4163_ = ~new_n3858_ & ~\quotient[41] ;
  assign new_n4164_ = ~new_n3868_ & new_n4122_;
  assign new_n4165_ = ~new_n4118_ & new_n4164_;
  assign new_n4166_ = ~new_n4119_ & ~new_n4122_;
  assign new_n4167_ = ~new_n4165_ & ~new_n4166_;
  assign new_n4168_ = new_n4143_ & ~new_n4167_;
  assign new_n4169_ = ~new_n4139_ & new_n4168_;
  assign new_n4170_ = ~new_n4163_ & ~new_n4169_;
  assign new_n4171_ = ~\b[20]  & ~new_n4170_;
  assign new_n4172_ = ~new_n3867_ & ~\quotient[41] ;
  assign new_n4173_ = ~new_n3877_ & new_n4117_;
  assign new_n4174_ = ~new_n4113_ & new_n4173_;
  assign new_n4175_ = ~new_n4114_ & ~new_n4117_;
  assign new_n4176_ = ~new_n4174_ & ~new_n4175_;
  assign new_n4177_ = new_n4143_ & ~new_n4176_;
  assign new_n4178_ = ~new_n4139_ & new_n4177_;
  assign new_n4179_ = ~new_n4172_ & ~new_n4178_;
  assign new_n4180_ = ~\b[19]  & ~new_n4179_;
  assign new_n4181_ = ~new_n3876_ & ~\quotient[41] ;
  assign new_n4182_ = ~new_n3886_ & new_n4112_;
  assign new_n4183_ = ~new_n4108_ & new_n4182_;
  assign new_n4184_ = ~new_n4109_ & ~new_n4112_;
  assign new_n4185_ = ~new_n4183_ & ~new_n4184_;
  assign new_n4186_ = new_n4143_ & ~new_n4185_;
  assign new_n4187_ = ~new_n4139_ & new_n4186_;
  assign new_n4188_ = ~new_n4181_ & ~new_n4187_;
  assign new_n4189_ = ~\b[18]  & ~new_n4188_;
  assign new_n4190_ = ~new_n3885_ & ~\quotient[41] ;
  assign new_n4191_ = ~new_n3895_ & new_n4107_;
  assign new_n4192_ = ~new_n4103_ & new_n4191_;
  assign new_n4193_ = ~new_n4104_ & ~new_n4107_;
  assign new_n4194_ = ~new_n4192_ & ~new_n4193_;
  assign new_n4195_ = new_n4143_ & ~new_n4194_;
  assign new_n4196_ = ~new_n4139_ & new_n4195_;
  assign new_n4197_ = ~new_n4190_ & ~new_n4196_;
  assign new_n4198_ = ~\b[17]  & ~new_n4197_;
  assign new_n4199_ = ~new_n3894_ & ~\quotient[41] ;
  assign new_n4200_ = ~new_n3904_ & new_n4102_;
  assign new_n4201_ = ~new_n4098_ & new_n4200_;
  assign new_n4202_ = ~new_n4099_ & ~new_n4102_;
  assign new_n4203_ = ~new_n4201_ & ~new_n4202_;
  assign new_n4204_ = new_n4143_ & ~new_n4203_;
  assign new_n4205_ = ~new_n4139_ & new_n4204_;
  assign new_n4206_ = ~new_n4199_ & ~new_n4205_;
  assign new_n4207_ = ~\b[16]  & ~new_n4206_;
  assign new_n4208_ = ~new_n3903_ & ~\quotient[41] ;
  assign new_n4209_ = ~new_n3913_ & new_n4097_;
  assign new_n4210_ = ~new_n4093_ & new_n4209_;
  assign new_n4211_ = ~new_n4094_ & ~new_n4097_;
  assign new_n4212_ = ~new_n4210_ & ~new_n4211_;
  assign new_n4213_ = new_n4143_ & ~new_n4212_;
  assign new_n4214_ = ~new_n4139_ & new_n4213_;
  assign new_n4215_ = ~new_n4208_ & ~new_n4214_;
  assign new_n4216_ = ~\b[15]  & ~new_n4215_;
  assign new_n4217_ = ~new_n3912_ & ~\quotient[41] ;
  assign new_n4218_ = ~new_n3922_ & new_n4092_;
  assign new_n4219_ = ~new_n4088_ & new_n4218_;
  assign new_n4220_ = ~new_n4089_ & ~new_n4092_;
  assign new_n4221_ = ~new_n4219_ & ~new_n4220_;
  assign new_n4222_ = new_n4143_ & ~new_n4221_;
  assign new_n4223_ = ~new_n4139_ & new_n4222_;
  assign new_n4224_ = ~new_n4217_ & ~new_n4223_;
  assign new_n4225_ = ~\b[14]  & ~new_n4224_;
  assign new_n4226_ = ~new_n3921_ & ~\quotient[41] ;
  assign new_n4227_ = ~new_n3931_ & new_n4087_;
  assign new_n4228_ = ~new_n4083_ & new_n4227_;
  assign new_n4229_ = ~new_n4084_ & ~new_n4087_;
  assign new_n4230_ = ~new_n4228_ & ~new_n4229_;
  assign new_n4231_ = new_n4143_ & ~new_n4230_;
  assign new_n4232_ = ~new_n4139_ & new_n4231_;
  assign new_n4233_ = ~new_n4226_ & ~new_n4232_;
  assign new_n4234_ = ~\b[13]  & ~new_n4233_;
  assign new_n4235_ = ~new_n3930_ & ~\quotient[41] ;
  assign new_n4236_ = ~new_n3940_ & new_n4082_;
  assign new_n4237_ = ~new_n4078_ & new_n4236_;
  assign new_n4238_ = ~new_n4079_ & ~new_n4082_;
  assign new_n4239_ = ~new_n4237_ & ~new_n4238_;
  assign new_n4240_ = new_n4143_ & ~new_n4239_;
  assign new_n4241_ = ~new_n4139_ & new_n4240_;
  assign new_n4242_ = ~new_n4235_ & ~new_n4241_;
  assign new_n4243_ = ~\b[12]  & ~new_n4242_;
  assign new_n4244_ = ~new_n3939_ & ~\quotient[41] ;
  assign new_n4245_ = ~new_n3949_ & new_n4077_;
  assign new_n4246_ = ~new_n4073_ & new_n4245_;
  assign new_n4247_ = ~new_n4074_ & ~new_n4077_;
  assign new_n4248_ = ~new_n4246_ & ~new_n4247_;
  assign new_n4249_ = new_n4143_ & ~new_n4248_;
  assign new_n4250_ = ~new_n4139_ & new_n4249_;
  assign new_n4251_ = ~new_n4244_ & ~new_n4250_;
  assign new_n4252_ = ~\b[11]  & ~new_n4251_;
  assign new_n4253_ = ~new_n3948_ & ~\quotient[41] ;
  assign new_n4254_ = ~new_n3958_ & new_n4072_;
  assign new_n4255_ = ~new_n4068_ & new_n4254_;
  assign new_n4256_ = ~new_n4069_ & ~new_n4072_;
  assign new_n4257_ = ~new_n4255_ & ~new_n4256_;
  assign new_n4258_ = new_n4143_ & ~new_n4257_;
  assign new_n4259_ = ~new_n4139_ & new_n4258_;
  assign new_n4260_ = ~new_n4253_ & ~new_n4259_;
  assign new_n4261_ = ~\b[10]  & ~new_n4260_;
  assign new_n4262_ = ~new_n3957_ & ~\quotient[41] ;
  assign new_n4263_ = ~new_n3967_ & new_n4067_;
  assign new_n4264_ = ~new_n4063_ & new_n4263_;
  assign new_n4265_ = ~new_n4064_ & ~new_n4067_;
  assign new_n4266_ = ~new_n4264_ & ~new_n4265_;
  assign new_n4267_ = new_n4143_ & ~new_n4266_;
  assign new_n4268_ = ~new_n4139_ & new_n4267_;
  assign new_n4269_ = ~new_n4262_ & ~new_n4268_;
  assign new_n4270_ = ~\b[9]  & ~new_n4269_;
  assign new_n4271_ = ~new_n3966_ & ~\quotient[41] ;
  assign new_n4272_ = ~new_n3976_ & new_n4062_;
  assign new_n4273_ = ~new_n4058_ & new_n4272_;
  assign new_n4274_ = ~new_n4059_ & ~new_n4062_;
  assign new_n4275_ = ~new_n4273_ & ~new_n4274_;
  assign new_n4276_ = new_n4143_ & ~new_n4275_;
  assign new_n4277_ = ~new_n4139_ & new_n4276_;
  assign new_n4278_ = ~new_n4271_ & ~new_n4277_;
  assign new_n4279_ = ~\b[8]  & ~new_n4278_;
  assign new_n4280_ = ~new_n3975_ & ~\quotient[41] ;
  assign new_n4281_ = ~new_n3985_ & new_n4057_;
  assign new_n4282_ = ~new_n4053_ & new_n4281_;
  assign new_n4283_ = ~new_n4054_ & ~new_n4057_;
  assign new_n4284_ = ~new_n4282_ & ~new_n4283_;
  assign new_n4285_ = new_n4143_ & ~new_n4284_;
  assign new_n4286_ = ~new_n4139_ & new_n4285_;
  assign new_n4287_ = ~new_n4280_ & ~new_n4286_;
  assign new_n4288_ = ~\b[7]  & ~new_n4287_;
  assign new_n4289_ = ~new_n3984_ & ~\quotient[41] ;
  assign new_n4290_ = ~new_n3994_ & new_n4052_;
  assign new_n4291_ = ~new_n4048_ & new_n4290_;
  assign new_n4292_ = ~new_n4049_ & ~new_n4052_;
  assign new_n4293_ = ~new_n4291_ & ~new_n4292_;
  assign new_n4294_ = new_n4143_ & ~new_n4293_;
  assign new_n4295_ = ~new_n4139_ & new_n4294_;
  assign new_n4296_ = ~new_n4289_ & ~new_n4295_;
  assign new_n4297_ = ~\b[6]  & ~new_n4296_;
  assign new_n4298_ = ~new_n3993_ & ~\quotient[41] ;
  assign new_n4299_ = ~new_n4003_ & new_n4047_;
  assign new_n4300_ = ~new_n4043_ & new_n4299_;
  assign new_n4301_ = ~new_n4044_ & ~new_n4047_;
  assign new_n4302_ = ~new_n4300_ & ~new_n4301_;
  assign new_n4303_ = new_n4143_ & ~new_n4302_;
  assign new_n4304_ = ~new_n4139_ & new_n4303_;
  assign new_n4305_ = ~new_n4298_ & ~new_n4304_;
  assign new_n4306_ = ~\b[5]  & ~new_n4305_;
  assign new_n4307_ = ~new_n4002_ & ~\quotient[41] ;
  assign new_n4308_ = ~new_n4011_ & new_n4042_;
  assign new_n4309_ = ~new_n4038_ & new_n4308_;
  assign new_n4310_ = ~new_n4039_ & ~new_n4042_;
  assign new_n4311_ = ~new_n4309_ & ~new_n4310_;
  assign new_n4312_ = new_n4143_ & ~new_n4311_;
  assign new_n4313_ = ~new_n4139_ & new_n4312_;
  assign new_n4314_ = ~new_n4307_ & ~new_n4313_;
  assign new_n4315_ = ~\b[4]  & ~new_n4314_;
  assign new_n4316_ = ~new_n4010_ & ~\quotient[41] ;
  assign new_n4317_ = ~new_n4033_ & new_n4037_;
  assign new_n4318_ = ~new_n4032_ & new_n4317_;
  assign new_n4319_ = ~new_n4034_ & ~new_n4037_;
  assign new_n4320_ = ~new_n4318_ & ~new_n4319_;
  assign new_n4321_ = new_n4143_ & ~new_n4320_;
  assign new_n4322_ = ~new_n4139_ & new_n4321_;
  assign new_n4323_ = ~new_n4316_ & ~new_n4322_;
  assign new_n4324_ = ~\b[3]  & ~new_n4323_;
  assign new_n4325_ = ~new_n4026_ & ~\quotient[41] ;
  assign new_n4326_ = ~new_n4029_ & new_n4031_;
  assign new_n4327_ = ~new_n4027_ & new_n4326_;
  assign new_n4328_ = new_n4143_ & ~new_n4327_;
  assign new_n4329_ = ~new_n4032_ & new_n4328_;
  assign new_n4330_ = ~new_n4139_ & new_n4329_;
  assign new_n4331_ = ~new_n4325_ & ~new_n4330_;
  assign new_n4332_ = ~\b[2]  & ~new_n4331_;
  assign new_n4333_ = \b[0]  & ~\b[23] ;
  assign new_n4334_ = new_n306_ & new_n4333_;
  assign new_n4335_ = new_n317_ & new_n4334_;
  assign new_n4336_ = new_n303_ & new_n4335_;
  assign new_n4337_ = new_n288_ & new_n4336_;
  assign new_n4338_ = ~new_n4139_ & new_n4337_;
  assign new_n4339_ = \a[41]  & ~new_n4338_;
  assign new_n4340_ = new_n365_ & new_n4031_;
  assign new_n4341_ = new_n376_ & new_n4340_;
  assign new_n4342_ = new_n588_ & new_n4341_;
  assign new_n4343_ = new_n598_ & new_n4342_;
  assign new_n4344_ = new_n595_ & new_n4343_;
  assign new_n4345_ = ~new_n4139_ & new_n4344_;
  assign new_n4346_ = ~new_n4339_ & ~new_n4345_;
  assign new_n4347_ = \b[1]  & ~new_n4346_;
  assign new_n4348_ = ~\b[1]  & ~new_n4345_;
  assign new_n4349_ = ~new_n4339_ & new_n4348_;
  assign new_n4350_ = ~new_n4347_ & ~new_n4349_;
  assign new_n4351_ = ~\a[40]  & \b[0] ;
  assign new_n4352_ = ~new_n4350_ & ~new_n4351_;
  assign new_n4353_ = ~\b[1]  & ~new_n4346_;
  assign new_n4354_ = ~new_n4352_ & ~new_n4353_;
  assign new_n4355_ = \b[2]  & ~new_n4330_;
  assign new_n4356_ = ~new_n4325_ & new_n4355_;
  assign new_n4357_ = ~new_n4332_ & ~new_n4356_;
  assign new_n4358_ = ~new_n4354_ & new_n4357_;
  assign new_n4359_ = ~new_n4332_ & ~new_n4358_;
  assign new_n4360_ = \b[3]  & ~new_n4322_;
  assign new_n4361_ = ~new_n4316_ & new_n4360_;
  assign new_n4362_ = ~new_n4324_ & ~new_n4361_;
  assign new_n4363_ = ~new_n4359_ & new_n4362_;
  assign new_n4364_ = ~new_n4324_ & ~new_n4363_;
  assign new_n4365_ = \b[4]  & ~new_n4313_;
  assign new_n4366_ = ~new_n4307_ & new_n4365_;
  assign new_n4367_ = ~new_n4315_ & ~new_n4366_;
  assign new_n4368_ = ~new_n4364_ & new_n4367_;
  assign new_n4369_ = ~new_n4315_ & ~new_n4368_;
  assign new_n4370_ = \b[5]  & ~new_n4304_;
  assign new_n4371_ = ~new_n4298_ & new_n4370_;
  assign new_n4372_ = ~new_n4306_ & ~new_n4371_;
  assign new_n4373_ = ~new_n4369_ & new_n4372_;
  assign new_n4374_ = ~new_n4306_ & ~new_n4373_;
  assign new_n4375_ = \b[6]  & ~new_n4295_;
  assign new_n4376_ = ~new_n4289_ & new_n4375_;
  assign new_n4377_ = ~new_n4297_ & ~new_n4376_;
  assign new_n4378_ = ~new_n4374_ & new_n4377_;
  assign new_n4379_ = ~new_n4297_ & ~new_n4378_;
  assign new_n4380_ = \b[7]  & ~new_n4286_;
  assign new_n4381_ = ~new_n4280_ & new_n4380_;
  assign new_n4382_ = ~new_n4288_ & ~new_n4381_;
  assign new_n4383_ = ~new_n4379_ & new_n4382_;
  assign new_n4384_ = ~new_n4288_ & ~new_n4383_;
  assign new_n4385_ = \b[8]  & ~new_n4277_;
  assign new_n4386_ = ~new_n4271_ & new_n4385_;
  assign new_n4387_ = ~new_n4279_ & ~new_n4386_;
  assign new_n4388_ = ~new_n4384_ & new_n4387_;
  assign new_n4389_ = ~new_n4279_ & ~new_n4388_;
  assign new_n4390_ = \b[9]  & ~new_n4268_;
  assign new_n4391_ = ~new_n4262_ & new_n4390_;
  assign new_n4392_ = ~new_n4270_ & ~new_n4391_;
  assign new_n4393_ = ~new_n4389_ & new_n4392_;
  assign new_n4394_ = ~new_n4270_ & ~new_n4393_;
  assign new_n4395_ = \b[10]  & ~new_n4259_;
  assign new_n4396_ = ~new_n4253_ & new_n4395_;
  assign new_n4397_ = ~new_n4261_ & ~new_n4396_;
  assign new_n4398_ = ~new_n4394_ & new_n4397_;
  assign new_n4399_ = ~new_n4261_ & ~new_n4398_;
  assign new_n4400_ = \b[11]  & ~new_n4250_;
  assign new_n4401_ = ~new_n4244_ & new_n4400_;
  assign new_n4402_ = ~new_n4252_ & ~new_n4401_;
  assign new_n4403_ = ~new_n4399_ & new_n4402_;
  assign new_n4404_ = ~new_n4252_ & ~new_n4403_;
  assign new_n4405_ = \b[12]  & ~new_n4241_;
  assign new_n4406_ = ~new_n4235_ & new_n4405_;
  assign new_n4407_ = ~new_n4243_ & ~new_n4406_;
  assign new_n4408_ = ~new_n4404_ & new_n4407_;
  assign new_n4409_ = ~new_n4243_ & ~new_n4408_;
  assign new_n4410_ = \b[13]  & ~new_n4232_;
  assign new_n4411_ = ~new_n4226_ & new_n4410_;
  assign new_n4412_ = ~new_n4234_ & ~new_n4411_;
  assign new_n4413_ = ~new_n4409_ & new_n4412_;
  assign new_n4414_ = ~new_n4234_ & ~new_n4413_;
  assign new_n4415_ = \b[14]  & ~new_n4223_;
  assign new_n4416_ = ~new_n4217_ & new_n4415_;
  assign new_n4417_ = ~new_n4225_ & ~new_n4416_;
  assign new_n4418_ = ~new_n4414_ & new_n4417_;
  assign new_n4419_ = ~new_n4225_ & ~new_n4418_;
  assign new_n4420_ = \b[15]  & ~new_n4214_;
  assign new_n4421_ = ~new_n4208_ & new_n4420_;
  assign new_n4422_ = ~new_n4216_ & ~new_n4421_;
  assign new_n4423_ = ~new_n4419_ & new_n4422_;
  assign new_n4424_ = ~new_n4216_ & ~new_n4423_;
  assign new_n4425_ = \b[16]  & ~new_n4205_;
  assign new_n4426_ = ~new_n4199_ & new_n4425_;
  assign new_n4427_ = ~new_n4207_ & ~new_n4426_;
  assign new_n4428_ = ~new_n4424_ & new_n4427_;
  assign new_n4429_ = ~new_n4207_ & ~new_n4428_;
  assign new_n4430_ = \b[17]  & ~new_n4196_;
  assign new_n4431_ = ~new_n4190_ & new_n4430_;
  assign new_n4432_ = ~new_n4198_ & ~new_n4431_;
  assign new_n4433_ = ~new_n4429_ & new_n4432_;
  assign new_n4434_ = ~new_n4198_ & ~new_n4433_;
  assign new_n4435_ = \b[18]  & ~new_n4187_;
  assign new_n4436_ = ~new_n4181_ & new_n4435_;
  assign new_n4437_ = ~new_n4189_ & ~new_n4436_;
  assign new_n4438_ = ~new_n4434_ & new_n4437_;
  assign new_n4439_ = ~new_n4189_ & ~new_n4438_;
  assign new_n4440_ = \b[19]  & ~new_n4178_;
  assign new_n4441_ = ~new_n4172_ & new_n4440_;
  assign new_n4442_ = ~new_n4180_ & ~new_n4441_;
  assign new_n4443_ = ~new_n4439_ & new_n4442_;
  assign new_n4444_ = ~new_n4180_ & ~new_n4443_;
  assign new_n4445_ = \b[20]  & ~new_n4169_;
  assign new_n4446_ = ~new_n4163_ & new_n4445_;
  assign new_n4447_ = ~new_n4171_ & ~new_n4446_;
  assign new_n4448_ = ~new_n4444_ & new_n4447_;
  assign new_n4449_ = ~new_n4171_ & ~new_n4448_;
  assign new_n4450_ = \b[21]  & ~new_n4160_;
  assign new_n4451_ = ~new_n4154_ & new_n4450_;
  assign new_n4452_ = ~new_n4162_ & ~new_n4451_;
  assign new_n4453_ = ~new_n4449_ & new_n4452_;
  assign new_n4454_ = ~new_n4162_ & ~new_n4453_;
  assign new_n4455_ = \b[22]  & ~new_n4151_;
  assign new_n4456_ = ~new_n4145_ & new_n4455_;
  assign new_n4457_ = ~new_n4153_ & ~new_n4456_;
  assign new_n4458_ = ~new_n4454_ & new_n4457_;
  assign new_n4459_ = ~new_n4153_ & ~new_n4458_;
  assign new_n4460_ = ~new_n3839_ & ~\quotient[41] ;
  assign new_n4461_ = ~new_n3841_ & new_n4137_;
  assign new_n4462_ = ~new_n4133_ & new_n4461_;
  assign new_n4463_ = ~new_n4134_ & ~new_n4137_;
  assign new_n4464_ = ~new_n4462_ & ~new_n4463_;
  assign new_n4465_ = \quotient[41]  & ~new_n4464_;
  assign new_n4466_ = ~new_n4460_ & ~new_n4465_;
  assign new_n4467_ = ~\b[23]  & ~new_n4466_;
  assign new_n4468_ = \b[23]  & ~new_n4460_;
  assign new_n4469_ = ~new_n4465_ & new_n4468_;
  assign new_n4470_ = new_n341_ & new_n343_;
  assign new_n4471_ = new_n338_ & new_n4470_;
  assign new_n4472_ = ~new_n4469_ & new_n4471_;
  assign new_n4473_ = ~new_n4467_ & new_n4472_;
  assign new_n4474_ = ~new_n4459_ & new_n4473_;
  assign new_n4475_ = new_n4143_ & ~new_n4466_;
  assign \quotient[40]  = new_n4474_ | new_n4475_;
  assign new_n4477_ = ~new_n4162_ & new_n4457_;
  assign new_n4478_ = ~new_n4453_ & new_n4477_;
  assign new_n4479_ = ~new_n4454_ & ~new_n4457_;
  assign new_n4480_ = ~new_n4478_ & ~new_n4479_;
  assign new_n4481_ = \quotient[40]  & ~new_n4480_;
  assign new_n4482_ = ~new_n4152_ & ~new_n4475_;
  assign new_n4483_ = ~new_n4474_ & new_n4482_;
  assign new_n4484_ = ~new_n4481_ & ~new_n4483_;
  assign new_n4485_ = ~new_n4153_ & ~new_n4469_;
  assign new_n4486_ = ~new_n4467_ & new_n4485_;
  assign new_n4487_ = ~new_n4458_ & new_n4486_;
  assign new_n4488_ = ~new_n4467_ & ~new_n4469_;
  assign new_n4489_ = ~new_n4459_ & ~new_n4488_;
  assign new_n4490_ = ~new_n4487_ & ~new_n4489_;
  assign new_n4491_ = \quotient[40]  & ~new_n4490_;
  assign new_n4492_ = ~new_n4466_ & ~new_n4475_;
  assign new_n4493_ = ~new_n4474_ & new_n4492_;
  assign new_n4494_ = ~new_n4491_ & ~new_n4493_;
  assign new_n4495_ = ~\b[24]  & ~new_n4494_;
  assign new_n4496_ = ~\b[23]  & ~new_n4484_;
  assign new_n4497_ = ~new_n4171_ & new_n4452_;
  assign new_n4498_ = ~new_n4448_ & new_n4497_;
  assign new_n4499_ = ~new_n4449_ & ~new_n4452_;
  assign new_n4500_ = ~new_n4498_ & ~new_n4499_;
  assign new_n4501_ = \quotient[40]  & ~new_n4500_;
  assign new_n4502_ = ~new_n4161_ & ~new_n4475_;
  assign new_n4503_ = ~new_n4474_ & new_n4502_;
  assign new_n4504_ = ~new_n4501_ & ~new_n4503_;
  assign new_n4505_ = ~\b[22]  & ~new_n4504_;
  assign new_n4506_ = ~new_n4180_ & new_n4447_;
  assign new_n4507_ = ~new_n4443_ & new_n4506_;
  assign new_n4508_ = ~new_n4444_ & ~new_n4447_;
  assign new_n4509_ = ~new_n4507_ & ~new_n4508_;
  assign new_n4510_ = \quotient[40]  & ~new_n4509_;
  assign new_n4511_ = ~new_n4170_ & ~new_n4475_;
  assign new_n4512_ = ~new_n4474_ & new_n4511_;
  assign new_n4513_ = ~new_n4510_ & ~new_n4512_;
  assign new_n4514_ = ~\b[21]  & ~new_n4513_;
  assign new_n4515_ = ~new_n4189_ & new_n4442_;
  assign new_n4516_ = ~new_n4438_ & new_n4515_;
  assign new_n4517_ = ~new_n4439_ & ~new_n4442_;
  assign new_n4518_ = ~new_n4516_ & ~new_n4517_;
  assign new_n4519_ = \quotient[40]  & ~new_n4518_;
  assign new_n4520_ = ~new_n4179_ & ~new_n4475_;
  assign new_n4521_ = ~new_n4474_ & new_n4520_;
  assign new_n4522_ = ~new_n4519_ & ~new_n4521_;
  assign new_n4523_ = ~\b[20]  & ~new_n4522_;
  assign new_n4524_ = ~new_n4198_ & new_n4437_;
  assign new_n4525_ = ~new_n4433_ & new_n4524_;
  assign new_n4526_ = ~new_n4434_ & ~new_n4437_;
  assign new_n4527_ = ~new_n4525_ & ~new_n4526_;
  assign new_n4528_ = \quotient[40]  & ~new_n4527_;
  assign new_n4529_ = ~new_n4188_ & ~new_n4475_;
  assign new_n4530_ = ~new_n4474_ & new_n4529_;
  assign new_n4531_ = ~new_n4528_ & ~new_n4530_;
  assign new_n4532_ = ~\b[19]  & ~new_n4531_;
  assign new_n4533_ = ~new_n4207_ & new_n4432_;
  assign new_n4534_ = ~new_n4428_ & new_n4533_;
  assign new_n4535_ = ~new_n4429_ & ~new_n4432_;
  assign new_n4536_ = ~new_n4534_ & ~new_n4535_;
  assign new_n4537_ = \quotient[40]  & ~new_n4536_;
  assign new_n4538_ = ~new_n4197_ & ~new_n4475_;
  assign new_n4539_ = ~new_n4474_ & new_n4538_;
  assign new_n4540_ = ~new_n4537_ & ~new_n4539_;
  assign new_n4541_ = ~\b[18]  & ~new_n4540_;
  assign new_n4542_ = ~new_n4216_ & new_n4427_;
  assign new_n4543_ = ~new_n4423_ & new_n4542_;
  assign new_n4544_ = ~new_n4424_ & ~new_n4427_;
  assign new_n4545_ = ~new_n4543_ & ~new_n4544_;
  assign new_n4546_ = \quotient[40]  & ~new_n4545_;
  assign new_n4547_ = ~new_n4206_ & ~new_n4475_;
  assign new_n4548_ = ~new_n4474_ & new_n4547_;
  assign new_n4549_ = ~new_n4546_ & ~new_n4548_;
  assign new_n4550_ = ~\b[17]  & ~new_n4549_;
  assign new_n4551_ = ~new_n4225_ & new_n4422_;
  assign new_n4552_ = ~new_n4418_ & new_n4551_;
  assign new_n4553_ = ~new_n4419_ & ~new_n4422_;
  assign new_n4554_ = ~new_n4552_ & ~new_n4553_;
  assign new_n4555_ = \quotient[40]  & ~new_n4554_;
  assign new_n4556_ = ~new_n4215_ & ~new_n4475_;
  assign new_n4557_ = ~new_n4474_ & new_n4556_;
  assign new_n4558_ = ~new_n4555_ & ~new_n4557_;
  assign new_n4559_ = ~\b[16]  & ~new_n4558_;
  assign new_n4560_ = ~new_n4234_ & new_n4417_;
  assign new_n4561_ = ~new_n4413_ & new_n4560_;
  assign new_n4562_ = ~new_n4414_ & ~new_n4417_;
  assign new_n4563_ = ~new_n4561_ & ~new_n4562_;
  assign new_n4564_ = \quotient[40]  & ~new_n4563_;
  assign new_n4565_ = ~new_n4224_ & ~new_n4475_;
  assign new_n4566_ = ~new_n4474_ & new_n4565_;
  assign new_n4567_ = ~new_n4564_ & ~new_n4566_;
  assign new_n4568_ = ~\b[15]  & ~new_n4567_;
  assign new_n4569_ = ~new_n4243_ & new_n4412_;
  assign new_n4570_ = ~new_n4408_ & new_n4569_;
  assign new_n4571_ = ~new_n4409_ & ~new_n4412_;
  assign new_n4572_ = ~new_n4570_ & ~new_n4571_;
  assign new_n4573_ = \quotient[40]  & ~new_n4572_;
  assign new_n4574_ = ~new_n4233_ & ~new_n4475_;
  assign new_n4575_ = ~new_n4474_ & new_n4574_;
  assign new_n4576_ = ~new_n4573_ & ~new_n4575_;
  assign new_n4577_ = ~\b[14]  & ~new_n4576_;
  assign new_n4578_ = ~new_n4252_ & new_n4407_;
  assign new_n4579_ = ~new_n4403_ & new_n4578_;
  assign new_n4580_ = ~new_n4404_ & ~new_n4407_;
  assign new_n4581_ = ~new_n4579_ & ~new_n4580_;
  assign new_n4582_ = \quotient[40]  & ~new_n4581_;
  assign new_n4583_ = ~new_n4242_ & ~new_n4475_;
  assign new_n4584_ = ~new_n4474_ & new_n4583_;
  assign new_n4585_ = ~new_n4582_ & ~new_n4584_;
  assign new_n4586_ = ~\b[13]  & ~new_n4585_;
  assign new_n4587_ = ~new_n4261_ & new_n4402_;
  assign new_n4588_ = ~new_n4398_ & new_n4587_;
  assign new_n4589_ = ~new_n4399_ & ~new_n4402_;
  assign new_n4590_ = ~new_n4588_ & ~new_n4589_;
  assign new_n4591_ = \quotient[40]  & ~new_n4590_;
  assign new_n4592_ = ~new_n4251_ & ~new_n4475_;
  assign new_n4593_ = ~new_n4474_ & new_n4592_;
  assign new_n4594_ = ~new_n4591_ & ~new_n4593_;
  assign new_n4595_ = ~\b[12]  & ~new_n4594_;
  assign new_n4596_ = ~new_n4270_ & new_n4397_;
  assign new_n4597_ = ~new_n4393_ & new_n4596_;
  assign new_n4598_ = ~new_n4394_ & ~new_n4397_;
  assign new_n4599_ = ~new_n4597_ & ~new_n4598_;
  assign new_n4600_ = \quotient[40]  & ~new_n4599_;
  assign new_n4601_ = ~new_n4260_ & ~new_n4475_;
  assign new_n4602_ = ~new_n4474_ & new_n4601_;
  assign new_n4603_ = ~new_n4600_ & ~new_n4602_;
  assign new_n4604_ = ~\b[11]  & ~new_n4603_;
  assign new_n4605_ = ~new_n4279_ & new_n4392_;
  assign new_n4606_ = ~new_n4388_ & new_n4605_;
  assign new_n4607_ = ~new_n4389_ & ~new_n4392_;
  assign new_n4608_ = ~new_n4606_ & ~new_n4607_;
  assign new_n4609_ = \quotient[40]  & ~new_n4608_;
  assign new_n4610_ = ~new_n4269_ & ~new_n4475_;
  assign new_n4611_ = ~new_n4474_ & new_n4610_;
  assign new_n4612_ = ~new_n4609_ & ~new_n4611_;
  assign new_n4613_ = ~\b[10]  & ~new_n4612_;
  assign new_n4614_ = ~new_n4288_ & new_n4387_;
  assign new_n4615_ = ~new_n4383_ & new_n4614_;
  assign new_n4616_ = ~new_n4384_ & ~new_n4387_;
  assign new_n4617_ = ~new_n4615_ & ~new_n4616_;
  assign new_n4618_ = \quotient[40]  & ~new_n4617_;
  assign new_n4619_ = ~new_n4278_ & ~new_n4475_;
  assign new_n4620_ = ~new_n4474_ & new_n4619_;
  assign new_n4621_ = ~new_n4618_ & ~new_n4620_;
  assign new_n4622_ = ~\b[9]  & ~new_n4621_;
  assign new_n4623_ = ~new_n4297_ & new_n4382_;
  assign new_n4624_ = ~new_n4378_ & new_n4623_;
  assign new_n4625_ = ~new_n4379_ & ~new_n4382_;
  assign new_n4626_ = ~new_n4624_ & ~new_n4625_;
  assign new_n4627_ = \quotient[40]  & ~new_n4626_;
  assign new_n4628_ = ~new_n4287_ & ~new_n4475_;
  assign new_n4629_ = ~new_n4474_ & new_n4628_;
  assign new_n4630_ = ~new_n4627_ & ~new_n4629_;
  assign new_n4631_ = ~\b[8]  & ~new_n4630_;
  assign new_n4632_ = ~new_n4306_ & new_n4377_;
  assign new_n4633_ = ~new_n4373_ & new_n4632_;
  assign new_n4634_ = ~new_n4374_ & ~new_n4377_;
  assign new_n4635_ = ~new_n4633_ & ~new_n4634_;
  assign new_n4636_ = \quotient[40]  & ~new_n4635_;
  assign new_n4637_ = ~new_n4296_ & ~new_n4475_;
  assign new_n4638_ = ~new_n4474_ & new_n4637_;
  assign new_n4639_ = ~new_n4636_ & ~new_n4638_;
  assign new_n4640_ = ~\b[7]  & ~new_n4639_;
  assign new_n4641_ = ~new_n4315_ & new_n4372_;
  assign new_n4642_ = ~new_n4368_ & new_n4641_;
  assign new_n4643_ = ~new_n4369_ & ~new_n4372_;
  assign new_n4644_ = ~new_n4642_ & ~new_n4643_;
  assign new_n4645_ = \quotient[40]  & ~new_n4644_;
  assign new_n4646_ = ~new_n4305_ & ~new_n4475_;
  assign new_n4647_ = ~new_n4474_ & new_n4646_;
  assign new_n4648_ = ~new_n4645_ & ~new_n4647_;
  assign new_n4649_ = ~\b[6]  & ~new_n4648_;
  assign new_n4650_ = ~new_n4324_ & new_n4367_;
  assign new_n4651_ = ~new_n4363_ & new_n4650_;
  assign new_n4652_ = ~new_n4364_ & ~new_n4367_;
  assign new_n4653_ = ~new_n4651_ & ~new_n4652_;
  assign new_n4654_ = \quotient[40]  & ~new_n4653_;
  assign new_n4655_ = ~new_n4314_ & ~new_n4475_;
  assign new_n4656_ = ~new_n4474_ & new_n4655_;
  assign new_n4657_ = ~new_n4654_ & ~new_n4656_;
  assign new_n4658_ = ~\b[5]  & ~new_n4657_;
  assign new_n4659_ = ~new_n4332_ & new_n4362_;
  assign new_n4660_ = ~new_n4358_ & new_n4659_;
  assign new_n4661_ = ~new_n4359_ & ~new_n4362_;
  assign new_n4662_ = ~new_n4660_ & ~new_n4661_;
  assign new_n4663_ = \quotient[40]  & ~new_n4662_;
  assign new_n4664_ = ~new_n4323_ & ~new_n4475_;
  assign new_n4665_ = ~new_n4474_ & new_n4664_;
  assign new_n4666_ = ~new_n4663_ & ~new_n4665_;
  assign new_n4667_ = ~\b[4]  & ~new_n4666_;
  assign new_n4668_ = ~new_n4353_ & new_n4357_;
  assign new_n4669_ = ~new_n4352_ & new_n4668_;
  assign new_n4670_ = ~new_n4354_ & ~new_n4357_;
  assign new_n4671_ = ~new_n4669_ & ~new_n4670_;
  assign new_n4672_ = \quotient[40]  & ~new_n4671_;
  assign new_n4673_ = ~new_n4331_ & ~new_n4475_;
  assign new_n4674_ = ~new_n4474_ & new_n4673_;
  assign new_n4675_ = ~new_n4672_ & ~new_n4674_;
  assign new_n4676_ = ~\b[3]  & ~new_n4675_;
  assign new_n4677_ = ~new_n4349_ & new_n4351_;
  assign new_n4678_ = ~new_n4347_ & new_n4677_;
  assign new_n4679_ = ~new_n4352_ & ~new_n4678_;
  assign new_n4680_ = \quotient[40]  & new_n4679_;
  assign new_n4681_ = ~new_n4346_ & ~new_n4475_;
  assign new_n4682_ = ~new_n4474_ & new_n4681_;
  assign new_n4683_ = ~new_n4680_ & ~new_n4682_;
  assign new_n4684_ = ~\b[2]  & ~new_n4683_;
  assign new_n4685_ = \b[0]  & \quotient[40] ;
  assign new_n4686_ = \a[40]  & ~new_n4685_;
  assign new_n4687_ = new_n4351_ & \quotient[40] ;
  assign new_n4688_ = ~new_n4686_ & ~new_n4687_;
  assign new_n4689_ = \b[1]  & ~new_n4688_;
  assign new_n4690_ = ~\b[1]  & ~new_n4687_;
  assign new_n4691_ = ~new_n4686_ & new_n4690_;
  assign new_n4692_ = ~new_n4689_ & ~new_n4691_;
  assign new_n4693_ = ~\a[39]  & \b[0] ;
  assign new_n4694_ = ~new_n4692_ & ~new_n4693_;
  assign new_n4695_ = ~\b[1]  & ~new_n4688_;
  assign new_n4696_ = ~new_n4694_ & ~new_n4695_;
  assign new_n4697_ = \b[2]  & ~new_n4682_;
  assign new_n4698_ = ~new_n4680_ & new_n4697_;
  assign new_n4699_ = ~new_n4684_ & ~new_n4698_;
  assign new_n4700_ = ~new_n4696_ & new_n4699_;
  assign new_n4701_ = ~new_n4684_ & ~new_n4700_;
  assign new_n4702_ = \b[3]  & ~new_n4674_;
  assign new_n4703_ = ~new_n4672_ & new_n4702_;
  assign new_n4704_ = ~new_n4676_ & ~new_n4703_;
  assign new_n4705_ = ~new_n4701_ & new_n4704_;
  assign new_n4706_ = ~new_n4676_ & ~new_n4705_;
  assign new_n4707_ = \b[4]  & ~new_n4665_;
  assign new_n4708_ = ~new_n4663_ & new_n4707_;
  assign new_n4709_ = ~new_n4667_ & ~new_n4708_;
  assign new_n4710_ = ~new_n4706_ & new_n4709_;
  assign new_n4711_ = ~new_n4667_ & ~new_n4710_;
  assign new_n4712_ = \b[5]  & ~new_n4656_;
  assign new_n4713_ = ~new_n4654_ & new_n4712_;
  assign new_n4714_ = ~new_n4658_ & ~new_n4713_;
  assign new_n4715_ = ~new_n4711_ & new_n4714_;
  assign new_n4716_ = ~new_n4658_ & ~new_n4715_;
  assign new_n4717_ = \b[6]  & ~new_n4647_;
  assign new_n4718_ = ~new_n4645_ & new_n4717_;
  assign new_n4719_ = ~new_n4649_ & ~new_n4718_;
  assign new_n4720_ = ~new_n4716_ & new_n4719_;
  assign new_n4721_ = ~new_n4649_ & ~new_n4720_;
  assign new_n4722_ = \b[7]  & ~new_n4638_;
  assign new_n4723_ = ~new_n4636_ & new_n4722_;
  assign new_n4724_ = ~new_n4640_ & ~new_n4723_;
  assign new_n4725_ = ~new_n4721_ & new_n4724_;
  assign new_n4726_ = ~new_n4640_ & ~new_n4725_;
  assign new_n4727_ = \b[8]  & ~new_n4629_;
  assign new_n4728_ = ~new_n4627_ & new_n4727_;
  assign new_n4729_ = ~new_n4631_ & ~new_n4728_;
  assign new_n4730_ = ~new_n4726_ & new_n4729_;
  assign new_n4731_ = ~new_n4631_ & ~new_n4730_;
  assign new_n4732_ = \b[9]  & ~new_n4620_;
  assign new_n4733_ = ~new_n4618_ & new_n4732_;
  assign new_n4734_ = ~new_n4622_ & ~new_n4733_;
  assign new_n4735_ = ~new_n4731_ & new_n4734_;
  assign new_n4736_ = ~new_n4622_ & ~new_n4735_;
  assign new_n4737_ = \b[10]  & ~new_n4611_;
  assign new_n4738_ = ~new_n4609_ & new_n4737_;
  assign new_n4739_ = ~new_n4613_ & ~new_n4738_;
  assign new_n4740_ = ~new_n4736_ & new_n4739_;
  assign new_n4741_ = ~new_n4613_ & ~new_n4740_;
  assign new_n4742_ = \b[11]  & ~new_n4602_;
  assign new_n4743_ = ~new_n4600_ & new_n4742_;
  assign new_n4744_ = ~new_n4604_ & ~new_n4743_;
  assign new_n4745_ = ~new_n4741_ & new_n4744_;
  assign new_n4746_ = ~new_n4604_ & ~new_n4745_;
  assign new_n4747_ = \b[12]  & ~new_n4593_;
  assign new_n4748_ = ~new_n4591_ & new_n4747_;
  assign new_n4749_ = ~new_n4595_ & ~new_n4748_;
  assign new_n4750_ = ~new_n4746_ & new_n4749_;
  assign new_n4751_ = ~new_n4595_ & ~new_n4750_;
  assign new_n4752_ = \b[13]  & ~new_n4584_;
  assign new_n4753_ = ~new_n4582_ & new_n4752_;
  assign new_n4754_ = ~new_n4586_ & ~new_n4753_;
  assign new_n4755_ = ~new_n4751_ & new_n4754_;
  assign new_n4756_ = ~new_n4586_ & ~new_n4755_;
  assign new_n4757_ = \b[14]  & ~new_n4575_;
  assign new_n4758_ = ~new_n4573_ & new_n4757_;
  assign new_n4759_ = ~new_n4577_ & ~new_n4758_;
  assign new_n4760_ = ~new_n4756_ & new_n4759_;
  assign new_n4761_ = ~new_n4577_ & ~new_n4760_;
  assign new_n4762_ = \b[15]  & ~new_n4566_;
  assign new_n4763_ = ~new_n4564_ & new_n4762_;
  assign new_n4764_ = ~new_n4568_ & ~new_n4763_;
  assign new_n4765_ = ~new_n4761_ & new_n4764_;
  assign new_n4766_ = ~new_n4568_ & ~new_n4765_;
  assign new_n4767_ = \b[16]  & ~new_n4557_;
  assign new_n4768_ = ~new_n4555_ & new_n4767_;
  assign new_n4769_ = ~new_n4559_ & ~new_n4768_;
  assign new_n4770_ = ~new_n4766_ & new_n4769_;
  assign new_n4771_ = ~new_n4559_ & ~new_n4770_;
  assign new_n4772_ = \b[17]  & ~new_n4548_;
  assign new_n4773_ = ~new_n4546_ & new_n4772_;
  assign new_n4774_ = ~new_n4550_ & ~new_n4773_;
  assign new_n4775_ = ~new_n4771_ & new_n4774_;
  assign new_n4776_ = ~new_n4550_ & ~new_n4775_;
  assign new_n4777_ = \b[18]  & ~new_n4539_;
  assign new_n4778_ = ~new_n4537_ & new_n4777_;
  assign new_n4779_ = ~new_n4541_ & ~new_n4778_;
  assign new_n4780_ = ~new_n4776_ & new_n4779_;
  assign new_n4781_ = ~new_n4541_ & ~new_n4780_;
  assign new_n4782_ = \b[19]  & ~new_n4530_;
  assign new_n4783_ = ~new_n4528_ & new_n4782_;
  assign new_n4784_ = ~new_n4532_ & ~new_n4783_;
  assign new_n4785_ = ~new_n4781_ & new_n4784_;
  assign new_n4786_ = ~new_n4532_ & ~new_n4785_;
  assign new_n4787_ = \b[20]  & ~new_n4521_;
  assign new_n4788_ = ~new_n4519_ & new_n4787_;
  assign new_n4789_ = ~new_n4523_ & ~new_n4788_;
  assign new_n4790_ = ~new_n4786_ & new_n4789_;
  assign new_n4791_ = ~new_n4523_ & ~new_n4790_;
  assign new_n4792_ = \b[21]  & ~new_n4512_;
  assign new_n4793_ = ~new_n4510_ & new_n4792_;
  assign new_n4794_ = ~new_n4514_ & ~new_n4793_;
  assign new_n4795_ = ~new_n4791_ & new_n4794_;
  assign new_n4796_ = ~new_n4514_ & ~new_n4795_;
  assign new_n4797_ = \b[22]  & ~new_n4503_;
  assign new_n4798_ = ~new_n4501_ & new_n4797_;
  assign new_n4799_ = ~new_n4505_ & ~new_n4798_;
  assign new_n4800_ = ~new_n4796_ & new_n4799_;
  assign new_n4801_ = ~new_n4505_ & ~new_n4800_;
  assign new_n4802_ = \b[23]  & ~new_n4483_;
  assign new_n4803_ = ~new_n4481_ & new_n4802_;
  assign new_n4804_ = ~new_n4496_ & ~new_n4803_;
  assign new_n4805_ = ~new_n4801_ & new_n4804_;
  assign new_n4806_ = ~new_n4496_ & ~new_n4805_;
  assign new_n4807_ = \b[24]  & ~new_n4493_;
  assign new_n4808_ = ~new_n4491_ & new_n4807_;
  assign new_n4809_ = ~new_n4495_ & ~new_n4808_;
  assign new_n4810_ = ~new_n4806_ & new_n4809_;
  assign new_n4811_ = ~new_n4495_ & ~new_n4810_;
  assign new_n4812_ = new_n377_ & new_n423_;
  assign new_n4813_ = new_n408_ & new_n4812_;
  assign \quotient[39]  = ~new_n4811_ & new_n4813_;
  assign new_n4815_ = ~new_n4484_ & ~\quotient[39] ;
  assign new_n4816_ = ~new_n4505_ & new_n4804_;
  assign new_n4817_ = ~new_n4800_ & new_n4816_;
  assign new_n4818_ = ~new_n4801_ & ~new_n4804_;
  assign new_n4819_ = ~new_n4817_ & ~new_n4818_;
  assign new_n4820_ = new_n4813_ & ~new_n4819_;
  assign new_n4821_ = ~new_n4811_ & new_n4820_;
  assign new_n4822_ = ~new_n4815_ & ~new_n4821_;
  assign new_n4823_ = ~new_n4494_ & ~\quotient[39] ;
  assign new_n4824_ = ~new_n4496_ & new_n4809_;
  assign new_n4825_ = ~new_n4805_ & new_n4824_;
  assign new_n4826_ = ~new_n4806_ & ~new_n4809_;
  assign new_n4827_ = ~new_n4825_ & ~new_n4826_;
  assign new_n4828_ = \quotient[39]  & ~new_n4827_;
  assign new_n4829_ = ~new_n4823_ & ~new_n4828_;
  assign new_n4830_ = ~\b[25]  & ~new_n4829_;
  assign new_n4831_ = ~\b[24]  & ~new_n4822_;
  assign new_n4832_ = ~new_n4504_ & ~\quotient[39] ;
  assign new_n4833_ = ~new_n4514_ & new_n4799_;
  assign new_n4834_ = ~new_n4795_ & new_n4833_;
  assign new_n4835_ = ~new_n4796_ & ~new_n4799_;
  assign new_n4836_ = ~new_n4834_ & ~new_n4835_;
  assign new_n4837_ = new_n4813_ & ~new_n4836_;
  assign new_n4838_ = ~new_n4811_ & new_n4837_;
  assign new_n4839_ = ~new_n4832_ & ~new_n4838_;
  assign new_n4840_ = ~\b[23]  & ~new_n4839_;
  assign new_n4841_ = ~new_n4513_ & ~\quotient[39] ;
  assign new_n4842_ = ~new_n4523_ & new_n4794_;
  assign new_n4843_ = ~new_n4790_ & new_n4842_;
  assign new_n4844_ = ~new_n4791_ & ~new_n4794_;
  assign new_n4845_ = ~new_n4843_ & ~new_n4844_;
  assign new_n4846_ = new_n4813_ & ~new_n4845_;
  assign new_n4847_ = ~new_n4811_ & new_n4846_;
  assign new_n4848_ = ~new_n4841_ & ~new_n4847_;
  assign new_n4849_ = ~\b[22]  & ~new_n4848_;
  assign new_n4850_ = ~new_n4522_ & ~\quotient[39] ;
  assign new_n4851_ = ~new_n4532_ & new_n4789_;
  assign new_n4852_ = ~new_n4785_ & new_n4851_;
  assign new_n4853_ = ~new_n4786_ & ~new_n4789_;
  assign new_n4854_ = ~new_n4852_ & ~new_n4853_;
  assign new_n4855_ = new_n4813_ & ~new_n4854_;
  assign new_n4856_ = ~new_n4811_ & new_n4855_;
  assign new_n4857_ = ~new_n4850_ & ~new_n4856_;
  assign new_n4858_ = ~\b[21]  & ~new_n4857_;
  assign new_n4859_ = ~new_n4531_ & ~\quotient[39] ;
  assign new_n4860_ = ~new_n4541_ & new_n4784_;
  assign new_n4861_ = ~new_n4780_ & new_n4860_;
  assign new_n4862_ = ~new_n4781_ & ~new_n4784_;
  assign new_n4863_ = ~new_n4861_ & ~new_n4862_;
  assign new_n4864_ = new_n4813_ & ~new_n4863_;
  assign new_n4865_ = ~new_n4811_ & new_n4864_;
  assign new_n4866_ = ~new_n4859_ & ~new_n4865_;
  assign new_n4867_ = ~\b[20]  & ~new_n4866_;
  assign new_n4868_ = ~new_n4540_ & ~\quotient[39] ;
  assign new_n4869_ = ~new_n4550_ & new_n4779_;
  assign new_n4870_ = ~new_n4775_ & new_n4869_;
  assign new_n4871_ = ~new_n4776_ & ~new_n4779_;
  assign new_n4872_ = ~new_n4870_ & ~new_n4871_;
  assign new_n4873_ = new_n4813_ & ~new_n4872_;
  assign new_n4874_ = ~new_n4811_ & new_n4873_;
  assign new_n4875_ = ~new_n4868_ & ~new_n4874_;
  assign new_n4876_ = ~\b[19]  & ~new_n4875_;
  assign new_n4877_ = ~new_n4549_ & ~\quotient[39] ;
  assign new_n4878_ = ~new_n4559_ & new_n4774_;
  assign new_n4879_ = ~new_n4770_ & new_n4878_;
  assign new_n4880_ = ~new_n4771_ & ~new_n4774_;
  assign new_n4881_ = ~new_n4879_ & ~new_n4880_;
  assign new_n4882_ = new_n4813_ & ~new_n4881_;
  assign new_n4883_ = ~new_n4811_ & new_n4882_;
  assign new_n4884_ = ~new_n4877_ & ~new_n4883_;
  assign new_n4885_ = ~\b[18]  & ~new_n4884_;
  assign new_n4886_ = ~new_n4558_ & ~\quotient[39] ;
  assign new_n4887_ = ~new_n4568_ & new_n4769_;
  assign new_n4888_ = ~new_n4765_ & new_n4887_;
  assign new_n4889_ = ~new_n4766_ & ~new_n4769_;
  assign new_n4890_ = ~new_n4888_ & ~new_n4889_;
  assign new_n4891_ = new_n4813_ & ~new_n4890_;
  assign new_n4892_ = ~new_n4811_ & new_n4891_;
  assign new_n4893_ = ~new_n4886_ & ~new_n4892_;
  assign new_n4894_ = ~\b[17]  & ~new_n4893_;
  assign new_n4895_ = ~new_n4567_ & ~\quotient[39] ;
  assign new_n4896_ = ~new_n4577_ & new_n4764_;
  assign new_n4897_ = ~new_n4760_ & new_n4896_;
  assign new_n4898_ = ~new_n4761_ & ~new_n4764_;
  assign new_n4899_ = ~new_n4897_ & ~new_n4898_;
  assign new_n4900_ = new_n4813_ & ~new_n4899_;
  assign new_n4901_ = ~new_n4811_ & new_n4900_;
  assign new_n4902_ = ~new_n4895_ & ~new_n4901_;
  assign new_n4903_ = ~\b[16]  & ~new_n4902_;
  assign new_n4904_ = ~new_n4576_ & ~\quotient[39] ;
  assign new_n4905_ = ~new_n4586_ & new_n4759_;
  assign new_n4906_ = ~new_n4755_ & new_n4905_;
  assign new_n4907_ = ~new_n4756_ & ~new_n4759_;
  assign new_n4908_ = ~new_n4906_ & ~new_n4907_;
  assign new_n4909_ = new_n4813_ & ~new_n4908_;
  assign new_n4910_ = ~new_n4811_ & new_n4909_;
  assign new_n4911_ = ~new_n4904_ & ~new_n4910_;
  assign new_n4912_ = ~\b[15]  & ~new_n4911_;
  assign new_n4913_ = ~new_n4585_ & ~\quotient[39] ;
  assign new_n4914_ = ~new_n4595_ & new_n4754_;
  assign new_n4915_ = ~new_n4750_ & new_n4914_;
  assign new_n4916_ = ~new_n4751_ & ~new_n4754_;
  assign new_n4917_ = ~new_n4915_ & ~new_n4916_;
  assign new_n4918_ = new_n4813_ & ~new_n4917_;
  assign new_n4919_ = ~new_n4811_ & new_n4918_;
  assign new_n4920_ = ~new_n4913_ & ~new_n4919_;
  assign new_n4921_ = ~\b[14]  & ~new_n4920_;
  assign new_n4922_ = ~new_n4594_ & ~\quotient[39] ;
  assign new_n4923_ = ~new_n4604_ & new_n4749_;
  assign new_n4924_ = ~new_n4745_ & new_n4923_;
  assign new_n4925_ = ~new_n4746_ & ~new_n4749_;
  assign new_n4926_ = ~new_n4924_ & ~new_n4925_;
  assign new_n4927_ = new_n4813_ & ~new_n4926_;
  assign new_n4928_ = ~new_n4811_ & new_n4927_;
  assign new_n4929_ = ~new_n4922_ & ~new_n4928_;
  assign new_n4930_ = ~\b[13]  & ~new_n4929_;
  assign new_n4931_ = ~new_n4603_ & ~\quotient[39] ;
  assign new_n4932_ = ~new_n4613_ & new_n4744_;
  assign new_n4933_ = ~new_n4740_ & new_n4932_;
  assign new_n4934_ = ~new_n4741_ & ~new_n4744_;
  assign new_n4935_ = ~new_n4933_ & ~new_n4934_;
  assign new_n4936_ = new_n4813_ & ~new_n4935_;
  assign new_n4937_ = ~new_n4811_ & new_n4936_;
  assign new_n4938_ = ~new_n4931_ & ~new_n4937_;
  assign new_n4939_ = ~\b[12]  & ~new_n4938_;
  assign new_n4940_ = ~new_n4612_ & ~\quotient[39] ;
  assign new_n4941_ = ~new_n4622_ & new_n4739_;
  assign new_n4942_ = ~new_n4735_ & new_n4941_;
  assign new_n4943_ = ~new_n4736_ & ~new_n4739_;
  assign new_n4944_ = ~new_n4942_ & ~new_n4943_;
  assign new_n4945_ = new_n4813_ & ~new_n4944_;
  assign new_n4946_ = ~new_n4811_ & new_n4945_;
  assign new_n4947_ = ~new_n4940_ & ~new_n4946_;
  assign new_n4948_ = ~\b[11]  & ~new_n4947_;
  assign new_n4949_ = ~new_n4621_ & ~\quotient[39] ;
  assign new_n4950_ = ~new_n4631_ & new_n4734_;
  assign new_n4951_ = ~new_n4730_ & new_n4950_;
  assign new_n4952_ = ~new_n4731_ & ~new_n4734_;
  assign new_n4953_ = ~new_n4951_ & ~new_n4952_;
  assign new_n4954_ = new_n4813_ & ~new_n4953_;
  assign new_n4955_ = ~new_n4811_ & new_n4954_;
  assign new_n4956_ = ~new_n4949_ & ~new_n4955_;
  assign new_n4957_ = ~\b[10]  & ~new_n4956_;
  assign new_n4958_ = ~new_n4630_ & ~\quotient[39] ;
  assign new_n4959_ = ~new_n4640_ & new_n4729_;
  assign new_n4960_ = ~new_n4725_ & new_n4959_;
  assign new_n4961_ = ~new_n4726_ & ~new_n4729_;
  assign new_n4962_ = ~new_n4960_ & ~new_n4961_;
  assign new_n4963_ = new_n4813_ & ~new_n4962_;
  assign new_n4964_ = ~new_n4811_ & new_n4963_;
  assign new_n4965_ = ~new_n4958_ & ~new_n4964_;
  assign new_n4966_ = ~\b[9]  & ~new_n4965_;
  assign new_n4967_ = ~new_n4639_ & ~\quotient[39] ;
  assign new_n4968_ = ~new_n4649_ & new_n4724_;
  assign new_n4969_ = ~new_n4720_ & new_n4968_;
  assign new_n4970_ = ~new_n4721_ & ~new_n4724_;
  assign new_n4971_ = ~new_n4969_ & ~new_n4970_;
  assign new_n4972_ = new_n4813_ & ~new_n4971_;
  assign new_n4973_ = ~new_n4811_ & new_n4972_;
  assign new_n4974_ = ~new_n4967_ & ~new_n4973_;
  assign new_n4975_ = ~\b[8]  & ~new_n4974_;
  assign new_n4976_ = ~new_n4648_ & ~\quotient[39] ;
  assign new_n4977_ = ~new_n4658_ & new_n4719_;
  assign new_n4978_ = ~new_n4715_ & new_n4977_;
  assign new_n4979_ = ~new_n4716_ & ~new_n4719_;
  assign new_n4980_ = ~new_n4978_ & ~new_n4979_;
  assign new_n4981_ = new_n4813_ & ~new_n4980_;
  assign new_n4982_ = ~new_n4811_ & new_n4981_;
  assign new_n4983_ = ~new_n4976_ & ~new_n4982_;
  assign new_n4984_ = ~\b[7]  & ~new_n4983_;
  assign new_n4985_ = ~new_n4657_ & ~\quotient[39] ;
  assign new_n4986_ = ~new_n4667_ & new_n4714_;
  assign new_n4987_ = ~new_n4710_ & new_n4986_;
  assign new_n4988_ = ~new_n4711_ & ~new_n4714_;
  assign new_n4989_ = ~new_n4987_ & ~new_n4988_;
  assign new_n4990_ = new_n4813_ & ~new_n4989_;
  assign new_n4991_ = ~new_n4811_ & new_n4990_;
  assign new_n4992_ = ~new_n4985_ & ~new_n4991_;
  assign new_n4993_ = ~\b[6]  & ~new_n4992_;
  assign new_n4994_ = ~new_n4666_ & ~\quotient[39] ;
  assign new_n4995_ = ~new_n4676_ & new_n4709_;
  assign new_n4996_ = ~new_n4705_ & new_n4995_;
  assign new_n4997_ = ~new_n4706_ & ~new_n4709_;
  assign new_n4998_ = ~new_n4996_ & ~new_n4997_;
  assign new_n4999_ = new_n4813_ & ~new_n4998_;
  assign new_n5000_ = ~new_n4811_ & new_n4999_;
  assign new_n5001_ = ~new_n4994_ & ~new_n5000_;
  assign new_n5002_ = ~\b[5]  & ~new_n5001_;
  assign new_n5003_ = ~new_n4675_ & ~\quotient[39] ;
  assign new_n5004_ = ~new_n4684_ & new_n4704_;
  assign new_n5005_ = ~new_n4700_ & new_n5004_;
  assign new_n5006_ = ~new_n4701_ & ~new_n4704_;
  assign new_n5007_ = ~new_n5005_ & ~new_n5006_;
  assign new_n5008_ = new_n4813_ & ~new_n5007_;
  assign new_n5009_ = ~new_n4811_ & new_n5008_;
  assign new_n5010_ = ~new_n5003_ & ~new_n5009_;
  assign new_n5011_ = ~\b[4]  & ~new_n5010_;
  assign new_n5012_ = ~new_n4683_ & ~\quotient[39] ;
  assign new_n5013_ = ~new_n4695_ & new_n4699_;
  assign new_n5014_ = ~new_n4694_ & new_n5013_;
  assign new_n5015_ = ~new_n4696_ & ~new_n4699_;
  assign new_n5016_ = ~new_n5014_ & ~new_n5015_;
  assign new_n5017_ = new_n4813_ & ~new_n5016_;
  assign new_n5018_ = ~new_n4811_ & new_n5017_;
  assign new_n5019_ = ~new_n5012_ & ~new_n5018_;
  assign new_n5020_ = ~\b[3]  & ~new_n5019_;
  assign new_n5021_ = ~new_n4688_ & ~\quotient[39] ;
  assign new_n5022_ = ~new_n4691_ & new_n4693_;
  assign new_n5023_ = ~new_n4689_ & new_n5022_;
  assign new_n5024_ = new_n4813_ & ~new_n5023_;
  assign new_n5025_ = ~new_n4694_ & new_n5024_;
  assign new_n5026_ = ~new_n4811_ & new_n5025_;
  assign new_n5027_ = ~new_n5021_ & ~new_n5026_;
  assign new_n5028_ = ~\b[2]  & ~new_n5027_;
  assign new_n5029_ = \b[0]  & ~\b[25] ;
  assign new_n5030_ = new_n305_ & new_n5029_;
  assign new_n5031_ = new_n316_ & new_n5030_;
  assign new_n5032_ = new_n341_ & new_n5031_;
  assign new_n5033_ = new_n338_ & new_n5032_;
  assign new_n5034_ = ~new_n4811_ & new_n5033_;
  assign new_n5035_ = \a[39]  & ~new_n5034_;
  assign new_n5036_ = new_n376_ & new_n4693_;
  assign new_n5037_ = new_n588_ & new_n5036_;
  assign new_n5038_ = new_n598_ & new_n5037_;
  assign new_n5039_ = new_n595_ & new_n5038_;
  assign new_n5040_ = ~new_n4811_ & new_n5039_;
  assign new_n5041_ = ~new_n5035_ & ~new_n5040_;
  assign new_n5042_ = \b[1]  & ~new_n5041_;
  assign new_n5043_ = ~\b[1]  & ~new_n5040_;
  assign new_n5044_ = ~new_n5035_ & new_n5043_;
  assign new_n5045_ = ~new_n5042_ & ~new_n5044_;
  assign new_n5046_ = ~\a[38]  & \b[0] ;
  assign new_n5047_ = ~new_n5045_ & ~new_n5046_;
  assign new_n5048_ = ~\b[1]  & ~new_n5041_;
  assign new_n5049_ = ~new_n5047_ & ~new_n5048_;
  assign new_n5050_ = \b[2]  & ~new_n5026_;
  assign new_n5051_ = ~new_n5021_ & new_n5050_;
  assign new_n5052_ = ~new_n5028_ & ~new_n5051_;
  assign new_n5053_ = ~new_n5049_ & new_n5052_;
  assign new_n5054_ = ~new_n5028_ & ~new_n5053_;
  assign new_n5055_ = \b[3]  & ~new_n5018_;
  assign new_n5056_ = ~new_n5012_ & new_n5055_;
  assign new_n5057_ = ~new_n5020_ & ~new_n5056_;
  assign new_n5058_ = ~new_n5054_ & new_n5057_;
  assign new_n5059_ = ~new_n5020_ & ~new_n5058_;
  assign new_n5060_ = \b[4]  & ~new_n5009_;
  assign new_n5061_ = ~new_n5003_ & new_n5060_;
  assign new_n5062_ = ~new_n5011_ & ~new_n5061_;
  assign new_n5063_ = ~new_n5059_ & new_n5062_;
  assign new_n5064_ = ~new_n5011_ & ~new_n5063_;
  assign new_n5065_ = \b[5]  & ~new_n5000_;
  assign new_n5066_ = ~new_n4994_ & new_n5065_;
  assign new_n5067_ = ~new_n5002_ & ~new_n5066_;
  assign new_n5068_ = ~new_n5064_ & new_n5067_;
  assign new_n5069_ = ~new_n5002_ & ~new_n5068_;
  assign new_n5070_ = \b[6]  & ~new_n4991_;
  assign new_n5071_ = ~new_n4985_ & new_n5070_;
  assign new_n5072_ = ~new_n4993_ & ~new_n5071_;
  assign new_n5073_ = ~new_n5069_ & new_n5072_;
  assign new_n5074_ = ~new_n4993_ & ~new_n5073_;
  assign new_n5075_ = \b[7]  & ~new_n4982_;
  assign new_n5076_ = ~new_n4976_ & new_n5075_;
  assign new_n5077_ = ~new_n4984_ & ~new_n5076_;
  assign new_n5078_ = ~new_n5074_ & new_n5077_;
  assign new_n5079_ = ~new_n4984_ & ~new_n5078_;
  assign new_n5080_ = \b[8]  & ~new_n4973_;
  assign new_n5081_ = ~new_n4967_ & new_n5080_;
  assign new_n5082_ = ~new_n4975_ & ~new_n5081_;
  assign new_n5083_ = ~new_n5079_ & new_n5082_;
  assign new_n5084_ = ~new_n4975_ & ~new_n5083_;
  assign new_n5085_ = \b[9]  & ~new_n4964_;
  assign new_n5086_ = ~new_n4958_ & new_n5085_;
  assign new_n5087_ = ~new_n4966_ & ~new_n5086_;
  assign new_n5088_ = ~new_n5084_ & new_n5087_;
  assign new_n5089_ = ~new_n4966_ & ~new_n5088_;
  assign new_n5090_ = \b[10]  & ~new_n4955_;
  assign new_n5091_ = ~new_n4949_ & new_n5090_;
  assign new_n5092_ = ~new_n4957_ & ~new_n5091_;
  assign new_n5093_ = ~new_n5089_ & new_n5092_;
  assign new_n5094_ = ~new_n4957_ & ~new_n5093_;
  assign new_n5095_ = \b[11]  & ~new_n4946_;
  assign new_n5096_ = ~new_n4940_ & new_n5095_;
  assign new_n5097_ = ~new_n4948_ & ~new_n5096_;
  assign new_n5098_ = ~new_n5094_ & new_n5097_;
  assign new_n5099_ = ~new_n4948_ & ~new_n5098_;
  assign new_n5100_ = \b[12]  & ~new_n4937_;
  assign new_n5101_ = ~new_n4931_ & new_n5100_;
  assign new_n5102_ = ~new_n4939_ & ~new_n5101_;
  assign new_n5103_ = ~new_n5099_ & new_n5102_;
  assign new_n5104_ = ~new_n4939_ & ~new_n5103_;
  assign new_n5105_ = \b[13]  & ~new_n4928_;
  assign new_n5106_ = ~new_n4922_ & new_n5105_;
  assign new_n5107_ = ~new_n4930_ & ~new_n5106_;
  assign new_n5108_ = ~new_n5104_ & new_n5107_;
  assign new_n5109_ = ~new_n4930_ & ~new_n5108_;
  assign new_n5110_ = \b[14]  & ~new_n4919_;
  assign new_n5111_ = ~new_n4913_ & new_n5110_;
  assign new_n5112_ = ~new_n4921_ & ~new_n5111_;
  assign new_n5113_ = ~new_n5109_ & new_n5112_;
  assign new_n5114_ = ~new_n4921_ & ~new_n5113_;
  assign new_n5115_ = \b[15]  & ~new_n4910_;
  assign new_n5116_ = ~new_n4904_ & new_n5115_;
  assign new_n5117_ = ~new_n4912_ & ~new_n5116_;
  assign new_n5118_ = ~new_n5114_ & new_n5117_;
  assign new_n5119_ = ~new_n4912_ & ~new_n5118_;
  assign new_n5120_ = \b[16]  & ~new_n4901_;
  assign new_n5121_ = ~new_n4895_ & new_n5120_;
  assign new_n5122_ = ~new_n4903_ & ~new_n5121_;
  assign new_n5123_ = ~new_n5119_ & new_n5122_;
  assign new_n5124_ = ~new_n4903_ & ~new_n5123_;
  assign new_n5125_ = \b[17]  & ~new_n4892_;
  assign new_n5126_ = ~new_n4886_ & new_n5125_;
  assign new_n5127_ = ~new_n4894_ & ~new_n5126_;
  assign new_n5128_ = ~new_n5124_ & new_n5127_;
  assign new_n5129_ = ~new_n4894_ & ~new_n5128_;
  assign new_n5130_ = \b[18]  & ~new_n4883_;
  assign new_n5131_ = ~new_n4877_ & new_n5130_;
  assign new_n5132_ = ~new_n4885_ & ~new_n5131_;
  assign new_n5133_ = ~new_n5129_ & new_n5132_;
  assign new_n5134_ = ~new_n4885_ & ~new_n5133_;
  assign new_n5135_ = \b[19]  & ~new_n4874_;
  assign new_n5136_ = ~new_n4868_ & new_n5135_;
  assign new_n5137_ = ~new_n4876_ & ~new_n5136_;
  assign new_n5138_ = ~new_n5134_ & new_n5137_;
  assign new_n5139_ = ~new_n4876_ & ~new_n5138_;
  assign new_n5140_ = \b[20]  & ~new_n4865_;
  assign new_n5141_ = ~new_n4859_ & new_n5140_;
  assign new_n5142_ = ~new_n4867_ & ~new_n5141_;
  assign new_n5143_ = ~new_n5139_ & new_n5142_;
  assign new_n5144_ = ~new_n4867_ & ~new_n5143_;
  assign new_n5145_ = \b[21]  & ~new_n4856_;
  assign new_n5146_ = ~new_n4850_ & new_n5145_;
  assign new_n5147_ = ~new_n4858_ & ~new_n5146_;
  assign new_n5148_ = ~new_n5144_ & new_n5147_;
  assign new_n5149_ = ~new_n4858_ & ~new_n5148_;
  assign new_n5150_ = \b[22]  & ~new_n4847_;
  assign new_n5151_ = ~new_n4841_ & new_n5150_;
  assign new_n5152_ = ~new_n4849_ & ~new_n5151_;
  assign new_n5153_ = ~new_n5149_ & new_n5152_;
  assign new_n5154_ = ~new_n4849_ & ~new_n5153_;
  assign new_n5155_ = \b[23]  & ~new_n4838_;
  assign new_n5156_ = ~new_n4832_ & new_n5155_;
  assign new_n5157_ = ~new_n4840_ & ~new_n5156_;
  assign new_n5158_ = ~new_n5154_ & new_n5157_;
  assign new_n5159_ = ~new_n4840_ & ~new_n5158_;
  assign new_n5160_ = \b[24]  & ~new_n4821_;
  assign new_n5161_ = ~new_n4815_ & new_n5160_;
  assign new_n5162_ = ~new_n4831_ & ~new_n5161_;
  assign new_n5163_ = ~new_n5159_ & new_n5162_;
  assign new_n5164_ = ~new_n4831_ & ~new_n5163_;
  assign new_n5165_ = \b[25]  & ~new_n4823_;
  assign new_n5166_ = ~new_n4828_ & new_n5165_;
  assign new_n5167_ = ~new_n4830_ & ~new_n5166_;
  assign new_n5168_ = ~new_n5164_ & new_n5167_;
  assign new_n5169_ = ~new_n4830_ & ~new_n5168_;
  assign new_n5170_ = new_n305_ & new_n316_;
  assign new_n5171_ = new_n341_ & new_n5170_;
  assign new_n5172_ = new_n338_ & new_n5171_;
  assign \quotient[38]  = ~new_n5169_ & new_n5172_;
  assign new_n5174_ = ~new_n4822_ & ~\quotient[38] ;
  assign new_n5175_ = ~new_n4840_ & new_n5162_;
  assign new_n5176_ = ~new_n5158_ & new_n5175_;
  assign new_n5177_ = ~new_n5159_ & ~new_n5162_;
  assign new_n5178_ = ~new_n5176_ & ~new_n5177_;
  assign new_n5179_ = new_n5172_ & ~new_n5178_;
  assign new_n5180_ = ~new_n5169_ & new_n5179_;
  assign new_n5181_ = ~new_n5174_ & ~new_n5180_;
  assign new_n5182_ = ~\b[25]  & ~new_n5181_;
  assign new_n5183_ = ~new_n4839_ & ~\quotient[38] ;
  assign new_n5184_ = ~new_n4849_ & new_n5157_;
  assign new_n5185_ = ~new_n5153_ & new_n5184_;
  assign new_n5186_ = ~new_n5154_ & ~new_n5157_;
  assign new_n5187_ = ~new_n5185_ & ~new_n5186_;
  assign new_n5188_ = new_n5172_ & ~new_n5187_;
  assign new_n5189_ = ~new_n5169_ & new_n5188_;
  assign new_n5190_ = ~new_n5183_ & ~new_n5189_;
  assign new_n5191_ = ~\b[24]  & ~new_n5190_;
  assign new_n5192_ = ~new_n4848_ & ~\quotient[38] ;
  assign new_n5193_ = ~new_n4858_ & new_n5152_;
  assign new_n5194_ = ~new_n5148_ & new_n5193_;
  assign new_n5195_ = ~new_n5149_ & ~new_n5152_;
  assign new_n5196_ = ~new_n5194_ & ~new_n5195_;
  assign new_n5197_ = new_n5172_ & ~new_n5196_;
  assign new_n5198_ = ~new_n5169_ & new_n5197_;
  assign new_n5199_ = ~new_n5192_ & ~new_n5198_;
  assign new_n5200_ = ~\b[23]  & ~new_n5199_;
  assign new_n5201_ = ~new_n4857_ & ~\quotient[38] ;
  assign new_n5202_ = ~new_n4867_ & new_n5147_;
  assign new_n5203_ = ~new_n5143_ & new_n5202_;
  assign new_n5204_ = ~new_n5144_ & ~new_n5147_;
  assign new_n5205_ = ~new_n5203_ & ~new_n5204_;
  assign new_n5206_ = new_n5172_ & ~new_n5205_;
  assign new_n5207_ = ~new_n5169_ & new_n5206_;
  assign new_n5208_ = ~new_n5201_ & ~new_n5207_;
  assign new_n5209_ = ~\b[22]  & ~new_n5208_;
  assign new_n5210_ = ~new_n4866_ & ~\quotient[38] ;
  assign new_n5211_ = ~new_n4876_ & new_n5142_;
  assign new_n5212_ = ~new_n5138_ & new_n5211_;
  assign new_n5213_ = ~new_n5139_ & ~new_n5142_;
  assign new_n5214_ = ~new_n5212_ & ~new_n5213_;
  assign new_n5215_ = new_n5172_ & ~new_n5214_;
  assign new_n5216_ = ~new_n5169_ & new_n5215_;
  assign new_n5217_ = ~new_n5210_ & ~new_n5216_;
  assign new_n5218_ = ~\b[21]  & ~new_n5217_;
  assign new_n5219_ = ~new_n4875_ & ~\quotient[38] ;
  assign new_n5220_ = ~new_n4885_ & new_n5137_;
  assign new_n5221_ = ~new_n5133_ & new_n5220_;
  assign new_n5222_ = ~new_n5134_ & ~new_n5137_;
  assign new_n5223_ = ~new_n5221_ & ~new_n5222_;
  assign new_n5224_ = new_n5172_ & ~new_n5223_;
  assign new_n5225_ = ~new_n5169_ & new_n5224_;
  assign new_n5226_ = ~new_n5219_ & ~new_n5225_;
  assign new_n5227_ = ~\b[20]  & ~new_n5226_;
  assign new_n5228_ = ~new_n4884_ & ~\quotient[38] ;
  assign new_n5229_ = ~new_n4894_ & new_n5132_;
  assign new_n5230_ = ~new_n5128_ & new_n5229_;
  assign new_n5231_ = ~new_n5129_ & ~new_n5132_;
  assign new_n5232_ = ~new_n5230_ & ~new_n5231_;
  assign new_n5233_ = new_n5172_ & ~new_n5232_;
  assign new_n5234_ = ~new_n5169_ & new_n5233_;
  assign new_n5235_ = ~new_n5228_ & ~new_n5234_;
  assign new_n5236_ = ~\b[19]  & ~new_n5235_;
  assign new_n5237_ = ~new_n4893_ & ~\quotient[38] ;
  assign new_n5238_ = ~new_n4903_ & new_n5127_;
  assign new_n5239_ = ~new_n5123_ & new_n5238_;
  assign new_n5240_ = ~new_n5124_ & ~new_n5127_;
  assign new_n5241_ = ~new_n5239_ & ~new_n5240_;
  assign new_n5242_ = new_n5172_ & ~new_n5241_;
  assign new_n5243_ = ~new_n5169_ & new_n5242_;
  assign new_n5244_ = ~new_n5237_ & ~new_n5243_;
  assign new_n5245_ = ~\b[18]  & ~new_n5244_;
  assign new_n5246_ = ~new_n4902_ & ~\quotient[38] ;
  assign new_n5247_ = ~new_n4912_ & new_n5122_;
  assign new_n5248_ = ~new_n5118_ & new_n5247_;
  assign new_n5249_ = ~new_n5119_ & ~new_n5122_;
  assign new_n5250_ = ~new_n5248_ & ~new_n5249_;
  assign new_n5251_ = new_n5172_ & ~new_n5250_;
  assign new_n5252_ = ~new_n5169_ & new_n5251_;
  assign new_n5253_ = ~new_n5246_ & ~new_n5252_;
  assign new_n5254_ = ~\b[17]  & ~new_n5253_;
  assign new_n5255_ = ~new_n4911_ & ~\quotient[38] ;
  assign new_n5256_ = ~new_n4921_ & new_n5117_;
  assign new_n5257_ = ~new_n5113_ & new_n5256_;
  assign new_n5258_ = ~new_n5114_ & ~new_n5117_;
  assign new_n5259_ = ~new_n5257_ & ~new_n5258_;
  assign new_n5260_ = new_n5172_ & ~new_n5259_;
  assign new_n5261_ = ~new_n5169_ & new_n5260_;
  assign new_n5262_ = ~new_n5255_ & ~new_n5261_;
  assign new_n5263_ = ~\b[16]  & ~new_n5262_;
  assign new_n5264_ = ~new_n4920_ & ~\quotient[38] ;
  assign new_n5265_ = ~new_n4930_ & new_n5112_;
  assign new_n5266_ = ~new_n5108_ & new_n5265_;
  assign new_n5267_ = ~new_n5109_ & ~new_n5112_;
  assign new_n5268_ = ~new_n5266_ & ~new_n5267_;
  assign new_n5269_ = new_n5172_ & ~new_n5268_;
  assign new_n5270_ = ~new_n5169_ & new_n5269_;
  assign new_n5271_ = ~new_n5264_ & ~new_n5270_;
  assign new_n5272_ = ~\b[15]  & ~new_n5271_;
  assign new_n5273_ = ~new_n4929_ & ~\quotient[38] ;
  assign new_n5274_ = ~new_n4939_ & new_n5107_;
  assign new_n5275_ = ~new_n5103_ & new_n5274_;
  assign new_n5276_ = ~new_n5104_ & ~new_n5107_;
  assign new_n5277_ = ~new_n5275_ & ~new_n5276_;
  assign new_n5278_ = new_n5172_ & ~new_n5277_;
  assign new_n5279_ = ~new_n5169_ & new_n5278_;
  assign new_n5280_ = ~new_n5273_ & ~new_n5279_;
  assign new_n5281_ = ~\b[14]  & ~new_n5280_;
  assign new_n5282_ = ~new_n4938_ & ~\quotient[38] ;
  assign new_n5283_ = ~new_n4948_ & new_n5102_;
  assign new_n5284_ = ~new_n5098_ & new_n5283_;
  assign new_n5285_ = ~new_n5099_ & ~new_n5102_;
  assign new_n5286_ = ~new_n5284_ & ~new_n5285_;
  assign new_n5287_ = new_n5172_ & ~new_n5286_;
  assign new_n5288_ = ~new_n5169_ & new_n5287_;
  assign new_n5289_ = ~new_n5282_ & ~new_n5288_;
  assign new_n5290_ = ~\b[13]  & ~new_n5289_;
  assign new_n5291_ = ~new_n4947_ & ~\quotient[38] ;
  assign new_n5292_ = ~new_n4957_ & new_n5097_;
  assign new_n5293_ = ~new_n5093_ & new_n5292_;
  assign new_n5294_ = ~new_n5094_ & ~new_n5097_;
  assign new_n5295_ = ~new_n5293_ & ~new_n5294_;
  assign new_n5296_ = new_n5172_ & ~new_n5295_;
  assign new_n5297_ = ~new_n5169_ & new_n5296_;
  assign new_n5298_ = ~new_n5291_ & ~new_n5297_;
  assign new_n5299_ = ~\b[12]  & ~new_n5298_;
  assign new_n5300_ = ~new_n4956_ & ~\quotient[38] ;
  assign new_n5301_ = ~new_n4966_ & new_n5092_;
  assign new_n5302_ = ~new_n5088_ & new_n5301_;
  assign new_n5303_ = ~new_n5089_ & ~new_n5092_;
  assign new_n5304_ = ~new_n5302_ & ~new_n5303_;
  assign new_n5305_ = new_n5172_ & ~new_n5304_;
  assign new_n5306_ = ~new_n5169_ & new_n5305_;
  assign new_n5307_ = ~new_n5300_ & ~new_n5306_;
  assign new_n5308_ = ~\b[11]  & ~new_n5307_;
  assign new_n5309_ = ~new_n4965_ & ~\quotient[38] ;
  assign new_n5310_ = ~new_n4975_ & new_n5087_;
  assign new_n5311_ = ~new_n5083_ & new_n5310_;
  assign new_n5312_ = ~new_n5084_ & ~new_n5087_;
  assign new_n5313_ = ~new_n5311_ & ~new_n5312_;
  assign new_n5314_ = new_n5172_ & ~new_n5313_;
  assign new_n5315_ = ~new_n5169_ & new_n5314_;
  assign new_n5316_ = ~new_n5309_ & ~new_n5315_;
  assign new_n5317_ = ~\b[10]  & ~new_n5316_;
  assign new_n5318_ = ~new_n4974_ & ~\quotient[38] ;
  assign new_n5319_ = ~new_n4984_ & new_n5082_;
  assign new_n5320_ = ~new_n5078_ & new_n5319_;
  assign new_n5321_ = ~new_n5079_ & ~new_n5082_;
  assign new_n5322_ = ~new_n5320_ & ~new_n5321_;
  assign new_n5323_ = new_n5172_ & ~new_n5322_;
  assign new_n5324_ = ~new_n5169_ & new_n5323_;
  assign new_n5325_ = ~new_n5318_ & ~new_n5324_;
  assign new_n5326_ = ~\b[9]  & ~new_n5325_;
  assign new_n5327_ = ~new_n4983_ & ~\quotient[38] ;
  assign new_n5328_ = ~new_n4993_ & new_n5077_;
  assign new_n5329_ = ~new_n5073_ & new_n5328_;
  assign new_n5330_ = ~new_n5074_ & ~new_n5077_;
  assign new_n5331_ = ~new_n5329_ & ~new_n5330_;
  assign new_n5332_ = new_n5172_ & ~new_n5331_;
  assign new_n5333_ = ~new_n5169_ & new_n5332_;
  assign new_n5334_ = ~new_n5327_ & ~new_n5333_;
  assign new_n5335_ = ~\b[8]  & ~new_n5334_;
  assign new_n5336_ = ~new_n4992_ & ~\quotient[38] ;
  assign new_n5337_ = ~new_n5002_ & new_n5072_;
  assign new_n5338_ = ~new_n5068_ & new_n5337_;
  assign new_n5339_ = ~new_n5069_ & ~new_n5072_;
  assign new_n5340_ = ~new_n5338_ & ~new_n5339_;
  assign new_n5341_ = new_n5172_ & ~new_n5340_;
  assign new_n5342_ = ~new_n5169_ & new_n5341_;
  assign new_n5343_ = ~new_n5336_ & ~new_n5342_;
  assign new_n5344_ = ~\b[7]  & ~new_n5343_;
  assign new_n5345_ = ~new_n5001_ & ~\quotient[38] ;
  assign new_n5346_ = ~new_n5011_ & new_n5067_;
  assign new_n5347_ = ~new_n5063_ & new_n5346_;
  assign new_n5348_ = ~new_n5064_ & ~new_n5067_;
  assign new_n5349_ = ~new_n5347_ & ~new_n5348_;
  assign new_n5350_ = new_n5172_ & ~new_n5349_;
  assign new_n5351_ = ~new_n5169_ & new_n5350_;
  assign new_n5352_ = ~new_n5345_ & ~new_n5351_;
  assign new_n5353_ = ~\b[6]  & ~new_n5352_;
  assign new_n5354_ = ~new_n5010_ & ~\quotient[38] ;
  assign new_n5355_ = ~new_n5020_ & new_n5062_;
  assign new_n5356_ = ~new_n5058_ & new_n5355_;
  assign new_n5357_ = ~new_n5059_ & ~new_n5062_;
  assign new_n5358_ = ~new_n5356_ & ~new_n5357_;
  assign new_n5359_ = new_n5172_ & ~new_n5358_;
  assign new_n5360_ = ~new_n5169_ & new_n5359_;
  assign new_n5361_ = ~new_n5354_ & ~new_n5360_;
  assign new_n5362_ = ~\b[5]  & ~new_n5361_;
  assign new_n5363_ = ~new_n5019_ & ~\quotient[38] ;
  assign new_n5364_ = ~new_n5028_ & new_n5057_;
  assign new_n5365_ = ~new_n5053_ & new_n5364_;
  assign new_n5366_ = ~new_n5054_ & ~new_n5057_;
  assign new_n5367_ = ~new_n5365_ & ~new_n5366_;
  assign new_n5368_ = new_n5172_ & ~new_n5367_;
  assign new_n5369_ = ~new_n5169_ & new_n5368_;
  assign new_n5370_ = ~new_n5363_ & ~new_n5369_;
  assign new_n5371_ = ~\b[4]  & ~new_n5370_;
  assign new_n5372_ = ~new_n5027_ & ~\quotient[38] ;
  assign new_n5373_ = ~new_n5048_ & new_n5052_;
  assign new_n5374_ = ~new_n5047_ & new_n5373_;
  assign new_n5375_ = ~new_n5049_ & ~new_n5052_;
  assign new_n5376_ = ~new_n5374_ & ~new_n5375_;
  assign new_n5377_ = new_n5172_ & ~new_n5376_;
  assign new_n5378_ = ~new_n5169_ & new_n5377_;
  assign new_n5379_ = ~new_n5372_ & ~new_n5378_;
  assign new_n5380_ = ~\b[3]  & ~new_n5379_;
  assign new_n5381_ = ~new_n5041_ & ~\quotient[38] ;
  assign new_n5382_ = ~new_n5044_ & new_n5046_;
  assign new_n5383_ = ~new_n5042_ & new_n5382_;
  assign new_n5384_ = new_n5172_ & ~new_n5383_;
  assign new_n5385_ = ~new_n5047_ & new_n5384_;
  assign new_n5386_ = ~new_n5169_ & new_n5385_;
  assign new_n5387_ = ~new_n5381_ & ~new_n5386_;
  assign new_n5388_ = ~\b[2]  & ~new_n5387_;
  assign new_n5389_ = \b[0]  & ~\b[26] ;
  assign new_n5390_ = new_n375_ & new_n5389_;
  assign new_n5391_ = new_n373_ & new_n5390_;
  assign new_n5392_ = new_n423_ & new_n5391_;
  assign new_n5393_ = new_n408_ & new_n5392_;
  assign new_n5394_ = ~new_n5169_ & new_n5393_;
  assign new_n5395_ = \a[38]  & ~new_n5394_;
  assign new_n5396_ = new_n305_ & new_n5046_;
  assign new_n5397_ = new_n316_ & new_n5396_;
  assign new_n5398_ = new_n341_ & new_n5397_;
  assign new_n5399_ = new_n338_ & new_n5398_;
  assign new_n5400_ = ~new_n5169_ & new_n5399_;
  assign new_n5401_ = ~new_n5395_ & ~new_n5400_;
  assign new_n5402_ = \b[1]  & ~new_n5401_;
  assign new_n5403_ = ~\b[1]  & ~new_n5400_;
  assign new_n5404_ = ~new_n5395_ & new_n5403_;
  assign new_n5405_ = ~new_n5402_ & ~new_n5404_;
  assign new_n5406_ = ~\a[37]  & \b[0] ;
  assign new_n5407_ = ~new_n5405_ & ~new_n5406_;
  assign new_n5408_ = ~\b[1]  & ~new_n5401_;
  assign new_n5409_ = ~new_n5407_ & ~new_n5408_;
  assign new_n5410_ = \b[2]  & ~new_n5386_;
  assign new_n5411_ = ~new_n5381_ & new_n5410_;
  assign new_n5412_ = ~new_n5388_ & ~new_n5411_;
  assign new_n5413_ = ~new_n5409_ & new_n5412_;
  assign new_n5414_ = ~new_n5388_ & ~new_n5413_;
  assign new_n5415_ = \b[3]  & ~new_n5378_;
  assign new_n5416_ = ~new_n5372_ & new_n5415_;
  assign new_n5417_ = ~new_n5380_ & ~new_n5416_;
  assign new_n5418_ = ~new_n5414_ & new_n5417_;
  assign new_n5419_ = ~new_n5380_ & ~new_n5418_;
  assign new_n5420_ = \b[4]  & ~new_n5369_;
  assign new_n5421_ = ~new_n5363_ & new_n5420_;
  assign new_n5422_ = ~new_n5371_ & ~new_n5421_;
  assign new_n5423_ = ~new_n5419_ & new_n5422_;
  assign new_n5424_ = ~new_n5371_ & ~new_n5423_;
  assign new_n5425_ = \b[5]  & ~new_n5360_;
  assign new_n5426_ = ~new_n5354_ & new_n5425_;
  assign new_n5427_ = ~new_n5362_ & ~new_n5426_;
  assign new_n5428_ = ~new_n5424_ & new_n5427_;
  assign new_n5429_ = ~new_n5362_ & ~new_n5428_;
  assign new_n5430_ = \b[6]  & ~new_n5351_;
  assign new_n5431_ = ~new_n5345_ & new_n5430_;
  assign new_n5432_ = ~new_n5353_ & ~new_n5431_;
  assign new_n5433_ = ~new_n5429_ & new_n5432_;
  assign new_n5434_ = ~new_n5353_ & ~new_n5433_;
  assign new_n5435_ = \b[7]  & ~new_n5342_;
  assign new_n5436_ = ~new_n5336_ & new_n5435_;
  assign new_n5437_ = ~new_n5344_ & ~new_n5436_;
  assign new_n5438_ = ~new_n5434_ & new_n5437_;
  assign new_n5439_ = ~new_n5344_ & ~new_n5438_;
  assign new_n5440_ = \b[8]  & ~new_n5333_;
  assign new_n5441_ = ~new_n5327_ & new_n5440_;
  assign new_n5442_ = ~new_n5335_ & ~new_n5441_;
  assign new_n5443_ = ~new_n5439_ & new_n5442_;
  assign new_n5444_ = ~new_n5335_ & ~new_n5443_;
  assign new_n5445_ = \b[9]  & ~new_n5324_;
  assign new_n5446_ = ~new_n5318_ & new_n5445_;
  assign new_n5447_ = ~new_n5326_ & ~new_n5446_;
  assign new_n5448_ = ~new_n5444_ & new_n5447_;
  assign new_n5449_ = ~new_n5326_ & ~new_n5448_;
  assign new_n5450_ = \b[10]  & ~new_n5315_;
  assign new_n5451_ = ~new_n5309_ & new_n5450_;
  assign new_n5452_ = ~new_n5317_ & ~new_n5451_;
  assign new_n5453_ = ~new_n5449_ & new_n5452_;
  assign new_n5454_ = ~new_n5317_ & ~new_n5453_;
  assign new_n5455_ = \b[11]  & ~new_n5306_;
  assign new_n5456_ = ~new_n5300_ & new_n5455_;
  assign new_n5457_ = ~new_n5308_ & ~new_n5456_;
  assign new_n5458_ = ~new_n5454_ & new_n5457_;
  assign new_n5459_ = ~new_n5308_ & ~new_n5458_;
  assign new_n5460_ = \b[12]  & ~new_n5297_;
  assign new_n5461_ = ~new_n5291_ & new_n5460_;
  assign new_n5462_ = ~new_n5299_ & ~new_n5461_;
  assign new_n5463_ = ~new_n5459_ & new_n5462_;
  assign new_n5464_ = ~new_n5299_ & ~new_n5463_;
  assign new_n5465_ = \b[13]  & ~new_n5288_;
  assign new_n5466_ = ~new_n5282_ & new_n5465_;
  assign new_n5467_ = ~new_n5290_ & ~new_n5466_;
  assign new_n5468_ = ~new_n5464_ & new_n5467_;
  assign new_n5469_ = ~new_n5290_ & ~new_n5468_;
  assign new_n5470_ = \b[14]  & ~new_n5279_;
  assign new_n5471_ = ~new_n5273_ & new_n5470_;
  assign new_n5472_ = ~new_n5281_ & ~new_n5471_;
  assign new_n5473_ = ~new_n5469_ & new_n5472_;
  assign new_n5474_ = ~new_n5281_ & ~new_n5473_;
  assign new_n5475_ = \b[15]  & ~new_n5270_;
  assign new_n5476_ = ~new_n5264_ & new_n5475_;
  assign new_n5477_ = ~new_n5272_ & ~new_n5476_;
  assign new_n5478_ = ~new_n5474_ & new_n5477_;
  assign new_n5479_ = ~new_n5272_ & ~new_n5478_;
  assign new_n5480_ = \b[16]  & ~new_n5261_;
  assign new_n5481_ = ~new_n5255_ & new_n5480_;
  assign new_n5482_ = ~new_n5263_ & ~new_n5481_;
  assign new_n5483_ = ~new_n5479_ & new_n5482_;
  assign new_n5484_ = ~new_n5263_ & ~new_n5483_;
  assign new_n5485_ = \b[17]  & ~new_n5252_;
  assign new_n5486_ = ~new_n5246_ & new_n5485_;
  assign new_n5487_ = ~new_n5254_ & ~new_n5486_;
  assign new_n5488_ = ~new_n5484_ & new_n5487_;
  assign new_n5489_ = ~new_n5254_ & ~new_n5488_;
  assign new_n5490_ = \b[18]  & ~new_n5243_;
  assign new_n5491_ = ~new_n5237_ & new_n5490_;
  assign new_n5492_ = ~new_n5245_ & ~new_n5491_;
  assign new_n5493_ = ~new_n5489_ & new_n5492_;
  assign new_n5494_ = ~new_n5245_ & ~new_n5493_;
  assign new_n5495_ = \b[19]  & ~new_n5234_;
  assign new_n5496_ = ~new_n5228_ & new_n5495_;
  assign new_n5497_ = ~new_n5236_ & ~new_n5496_;
  assign new_n5498_ = ~new_n5494_ & new_n5497_;
  assign new_n5499_ = ~new_n5236_ & ~new_n5498_;
  assign new_n5500_ = \b[20]  & ~new_n5225_;
  assign new_n5501_ = ~new_n5219_ & new_n5500_;
  assign new_n5502_ = ~new_n5227_ & ~new_n5501_;
  assign new_n5503_ = ~new_n5499_ & new_n5502_;
  assign new_n5504_ = ~new_n5227_ & ~new_n5503_;
  assign new_n5505_ = \b[21]  & ~new_n5216_;
  assign new_n5506_ = ~new_n5210_ & new_n5505_;
  assign new_n5507_ = ~new_n5218_ & ~new_n5506_;
  assign new_n5508_ = ~new_n5504_ & new_n5507_;
  assign new_n5509_ = ~new_n5218_ & ~new_n5508_;
  assign new_n5510_ = \b[22]  & ~new_n5207_;
  assign new_n5511_ = ~new_n5201_ & new_n5510_;
  assign new_n5512_ = ~new_n5209_ & ~new_n5511_;
  assign new_n5513_ = ~new_n5509_ & new_n5512_;
  assign new_n5514_ = ~new_n5209_ & ~new_n5513_;
  assign new_n5515_ = \b[23]  & ~new_n5198_;
  assign new_n5516_ = ~new_n5192_ & new_n5515_;
  assign new_n5517_ = ~new_n5200_ & ~new_n5516_;
  assign new_n5518_ = ~new_n5514_ & new_n5517_;
  assign new_n5519_ = ~new_n5200_ & ~new_n5518_;
  assign new_n5520_ = \b[24]  & ~new_n5189_;
  assign new_n5521_ = ~new_n5183_ & new_n5520_;
  assign new_n5522_ = ~new_n5191_ & ~new_n5521_;
  assign new_n5523_ = ~new_n5519_ & new_n5522_;
  assign new_n5524_ = ~new_n5191_ & ~new_n5523_;
  assign new_n5525_ = \b[25]  & ~new_n5180_;
  assign new_n5526_ = ~new_n5174_ & new_n5525_;
  assign new_n5527_ = ~new_n5182_ & ~new_n5526_;
  assign new_n5528_ = ~new_n5524_ & new_n5527_;
  assign new_n5529_ = ~new_n5182_ & ~new_n5528_;
  assign new_n5530_ = ~new_n4829_ & ~\quotient[38] ;
  assign new_n5531_ = ~new_n4831_ & new_n5167_;
  assign new_n5532_ = ~new_n5163_ & new_n5531_;
  assign new_n5533_ = ~new_n5164_ & ~new_n5167_;
  assign new_n5534_ = ~new_n5532_ & ~new_n5533_;
  assign new_n5535_ = \quotient[38]  & ~new_n5534_;
  assign new_n5536_ = ~new_n5530_ & ~new_n5535_;
  assign new_n5537_ = ~\b[26]  & ~new_n5536_;
  assign new_n5538_ = \b[26]  & ~new_n5530_;
  assign new_n5539_ = ~new_n5535_ & new_n5538_;
  assign new_n5540_ = new_n373_ & new_n375_;
  assign new_n5541_ = new_n423_ & new_n5540_;
  assign new_n5542_ = new_n408_ & new_n5541_;
  assign new_n5543_ = ~new_n5539_ & new_n5542_;
  assign new_n5544_ = ~new_n5537_ & new_n5543_;
  assign new_n5545_ = ~new_n5529_ & new_n5544_;
  assign new_n5546_ = new_n5172_ & ~new_n5536_;
  assign \quotient[37]  = new_n5545_ | new_n5546_;
  assign new_n5548_ = ~new_n5191_ & new_n5527_;
  assign new_n5549_ = ~new_n5523_ & new_n5548_;
  assign new_n5550_ = ~new_n5524_ & ~new_n5527_;
  assign new_n5551_ = ~new_n5549_ & ~new_n5550_;
  assign new_n5552_ = \quotient[37]  & ~new_n5551_;
  assign new_n5553_ = ~new_n5181_ & ~new_n5546_;
  assign new_n5554_ = ~new_n5545_ & new_n5553_;
  assign new_n5555_ = ~new_n5552_ & ~new_n5554_;
  assign new_n5556_ = ~new_n5182_ & ~new_n5539_;
  assign new_n5557_ = ~new_n5537_ & new_n5556_;
  assign new_n5558_ = ~new_n5528_ & new_n5557_;
  assign new_n5559_ = ~new_n5537_ & ~new_n5539_;
  assign new_n5560_ = ~new_n5529_ & ~new_n5559_;
  assign new_n5561_ = ~new_n5558_ & ~new_n5560_;
  assign new_n5562_ = \quotient[37]  & ~new_n5561_;
  assign new_n5563_ = ~new_n5536_ & ~new_n5546_;
  assign new_n5564_ = ~new_n5545_ & new_n5563_;
  assign new_n5565_ = ~new_n5562_ & ~new_n5564_;
  assign new_n5566_ = ~\b[27]  & ~new_n5565_;
  assign new_n5567_ = ~\b[26]  & ~new_n5555_;
  assign new_n5568_ = ~new_n5200_ & new_n5522_;
  assign new_n5569_ = ~new_n5518_ & new_n5568_;
  assign new_n5570_ = ~new_n5519_ & ~new_n5522_;
  assign new_n5571_ = ~new_n5569_ & ~new_n5570_;
  assign new_n5572_ = \quotient[37]  & ~new_n5571_;
  assign new_n5573_ = ~new_n5190_ & ~new_n5546_;
  assign new_n5574_ = ~new_n5545_ & new_n5573_;
  assign new_n5575_ = ~new_n5572_ & ~new_n5574_;
  assign new_n5576_ = ~\b[25]  & ~new_n5575_;
  assign new_n5577_ = ~new_n5209_ & new_n5517_;
  assign new_n5578_ = ~new_n5513_ & new_n5577_;
  assign new_n5579_ = ~new_n5514_ & ~new_n5517_;
  assign new_n5580_ = ~new_n5578_ & ~new_n5579_;
  assign new_n5581_ = \quotient[37]  & ~new_n5580_;
  assign new_n5582_ = ~new_n5199_ & ~new_n5546_;
  assign new_n5583_ = ~new_n5545_ & new_n5582_;
  assign new_n5584_ = ~new_n5581_ & ~new_n5583_;
  assign new_n5585_ = ~\b[24]  & ~new_n5584_;
  assign new_n5586_ = ~new_n5218_ & new_n5512_;
  assign new_n5587_ = ~new_n5508_ & new_n5586_;
  assign new_n5588_ = ~new_n5509_ & ~new_n5512_;
  assign new_n5589_ = ~new_n5587_ & ~new_n5588_;
  assign new_n5590_ = \quotient[37]  & ~new_n5589_;
  assign new_n5591_ = ~new_n5208_ & ~new_n5546_;
  assign new_n5592_ = ~new_n5545_ & new_n5591_;
  assign new_n5593_ = ~new_n5590_ & ~new_n5592_;
  assign new_n5594_ = ~\b[23]  & ~new_n5593_;
  assign new_n5595_ = ~new_n5227_ & new_n5507_;
  assign new_n5596_ = ~new_n5503_ & new_n5595_;
  assign new_n5597_ = ~new_n5504_ & ~new_n5507_;
  assign new_n5598_ = ~new_n5596_ & ~new_n5597_;
  assign new_n5599_ = \quotient[37]  & ~new_n5598_;
  assign new_n5600_ = ~new_n5217_ & ~new_n5546_;
  assign new_n5601_ = ~new_n5545_ & new_n5600_;
  assign new_n5602_ = ~new_n5599_ & ~new_n5601_;
  assign new_n5603_ = ~\b[22]  & ~new_n5602_;
  assign new_n5604_ = ~new_n5236_ & new_n5502_;
  assign new_n5605_ = ~new_n5498_ & new_n5604_;
  assign new_n5606_ = ~new_n5499_ & ~new_n5502_;
  assign new_n5607_ = ~new_n5605_ & ~new_n5606_;
  assign new_n5608_ = \quotient[37]  & ~new_n5607_;
  assign new_n5609_ = ~new_n5226_ & ~new_n5546_;
  assign new_n5610_ = ~new_n5545_ & new_n5609_;
  assign new_n5611_ = ~new_n5608_ & ~new_n5610_;
  assign new_n5612_ = ~\b[21]  & ~new_n5611_;
  assign new_n5613_ = ~new_n5245_ & new_n5497_;
  assign new_n5614_ = ~new_n5493_ & new_n5613_;
  assign new_n5615_ = ~new_n5494_ & ~new_n5497_;
  assign new_n5616_ = ~new_n5614_ & ~new_n5615_;
  assign new_n5617_ = \quotient[37]  & ~new_n5616_;
  assign new_n5618_ = ~new_n5235_ & ~new_n5546_;
  assign new_n5619_ = ~new_n5545_ & new_n5618_;
  assign new_n5620_ = ~new_n5617_ & ~new_n5619_;
  assign new_n5621_ = ~\b[20]  & ~new_n5620_;
  assign new_n5622_ = ~new_n5254_ & new_n5492_;
  assign new_n5623_ = ~new_n5488_ & new_n5622_;
  assign new_n5624_ = ~new_n5489_ & ~new_n5492_;
  assign new_n5625_ = ~new_n5623_ & ~new_n5624_;
  assign new_n5626_ = \quotient[37]  & ~new_n5625_;
  assign new_n5627_ = ~new_n5244_ & ~new_n5546_;
  assign new_n5628_ = ~new_n5545_ & new_n5627_;
  assign new_n5629_ = ~new_n5626_ & ~new_n5628_;
  assign new_n5630_ = ~\b[19]  & ~new_n5629_;
  assign new_n5631_ = ~new_n5263_ & new_n5487_;
  assign new_n5632_ = ~new_n5483_ & new_n5631_;
  assign new_n5633_ = ~new_n5484_ & ~new_n5487_;
  assign new_n5634_ = ~new_n5632_ & ~new_n5633_;
  assign new_n5635_ = \quotient[37]  & ~new_n5634_;
  assign new_n5636_ = ~new_n5253_ & ~new_n5546_;
  assign new_n5637_ = ~new_n5545_ & new_n5636_;
  assign new_n5638_ = ~new_n5635_ & ~new_n5637_;
  assign new_n5639_ = ~\b[18]  & ~new_n5638_;
  assign new_n5640_ = ~new_n5272_ & new_n5482_;
  assign new_n5641_ = ~new_n5478_ & new_n5640_;
  assign new_n5642_ = ~new_n5479_ & ~new_n5482_;
  assign new_n5643_ = ~new_n5641_ & ~new_n5642_;
  assign new_n5644_ = \quotient[37]  & ~new_n5643_;
  assign new_n5645_ = ~new_n5262_ & ~new_n5546_;
  assign new_n5646_ = ~new_n5545_ & new_n5645_;
  assign new_n5647_ = ~new_n5644_ & ~new_n5646_;
  assign new_n5648_ = ~\b[17]  & ~new_n5647_;
  assign new_n5649_ = ~new_n5281_ & new_n5477_;
  assign new_n5650_ = ~new_n5473_ & new_n5649_;
  assign new_n5651_ = ~new_n5474_ & ~new_n5477_;
  assign new_n5652_ = ~new_n5650_ & ~new_n5651_;
  assign new_n5653_ = \quotient[37]  & ~new_n5652_;
  assign new_n5654_ = ~new_n5271_ & ~new_n5546_;
  assign new_n5655_ = ~new_n5545_ & new_n5654_;
  assign new_n5656_ = ~new_n5653_ & ~new_n5655_;
  assign new_n5657_ = ~\b[16]  & ~new_n5656_;
  assign new_n5658_ = ~new_n5290_ & new_n5472_;
  assign new_n5659_ = ~new_n5468_ & new_n5658_;
  assign new_n5660_ = ~new_n5469_ & ~new_n5472_;
  assign new_n5661_ = ~new_n5659_ & ~new_n5660_;
  assign new_n5662_ = \quotient[37]  & ~new_n5661_;
  assign new_n5663_ = ~new_n5280_ & ~new_n5546_;
  assign new_n5664_ = ~new_n5545_ & new_n5663_;
  assign new_n5665_ = ~new_n5662_ & ~new_n5664_;
  assign new_n5666_ = ~\b[15]  & ~new_n5665_;
  assign new_n5667_ = ~new_n5299_ & new_n5467_;
  assign new_n5668_ = ~new_n5463_ & new_n5667_;
  assign new_n5669_ = ~new_n5464_ & ~new_n5467_;
  assign new_n5670_ = ~new_n5668_ & ~new_n5669_;
  assign new_n5671_ = \quotient[37]  & ~new_n5670_;
  assign new_n5672_ = ~new_n5289_ & ~new_n5546_;
  assign new_n5673_ = ~new_n5545_ & new_n5672_;
  assign new_n5674_ = ~new_n5671_ & ~new_n5673_;
  assign new_n5675_ = ~\b[14]  & ~new_n5674_;
  assign new_n5676_ = ~new_n5308_ & new_n5462_;
  assign new_n5677_ = ~new_n5458_ & new_n5676_;
  assign new_n5678_ = ~new_n5459_ & ~new_n5462_;
  assign new_n5679_ = ~new_n5677_ & ~new_n5678_;
  assign new_n5680_ = \quotient[37]  & ~new_n5679_;
  assign new_n5681_ = ~new_n5298_ & ~new_n5546_;
  assign new_n5682_ = ~new_n5545_ & new_n5681_;
  assign new_n5683_ = ~new_n5680_ & ~new_n5682_;
  assign new_n5684_ = ~\b[13]  & ~new_n5683_;
  assign new_n5685_ = ~new_n5317_ & new_n5457_;
  assign new_n5686_ = ~new_n5453_ & new_n5685_;
  assign new_n5687_ = ~new_n5454_ & ~new_n5457_;
  assign new_n5688_ = ~new_n5686_ & ~new_n5687_;
  assign new_n5689_ = \quotient[37]  & ~new_n5688_;
  assign new_n5690_ = ~new_n5307_ & ~new_n5546_;
  assign new_n5691_ = ~new_n5545_ & new_n5690_;
  assign new_n5692_ = ~new_n5689_ & ~new_n5691_;
  assign new_n5693_ = ~\b[12]  & ~new_n5692_;
  assign new_n5694_ = ~new_n5326_ & new_n5452_;
  assign new_n5695_ = ~new_n5448_ & new_n5694_;
  assign new_n5696_ = ~new_n5449_ & ~new_n5452_;
  assign new_n5697_ = ~new_n5695_ & ~new_n5696_;
  assign new_n5698_ = \quotient[37]  & ~new_n5697_;
  assign new_n5699_ = ~new_n5316_ & ~new_n5546_;
  assign new_n5700_ = ~new_n5545_ & new_n5699_;
  assign new_n5701_ = ~new_n5698_ & ~new_n5700_;
  assign new_n5702_ = ~\b[11]  & ~new_n5701_;
  assign new_n5703_ = ~new_n5335_ & new_n5447_;
  assign new_n5704_ = ~new_n5443_ & new_n5703_;
  assign new_n5705_ = ~new_n5444_ & ~new_n5447_;
  assign new_n5706_ = ~new_n5704_ & ~new_n5705_;
  assign new_n5707_ = \quotient[37]  & ~new_n5706_;
  assign new_n5708_ = ~new_n5325_ & ~new_n5546_;
  assign new_n5709_ = ~new_n5545_ & new_n5708_;
  assign new_n5710_ = ~new_n5707_ & ~new_n5709_;
  assign new_n5711_ = ~\b[10]  & ~new_n5710_;
  assign new_n5712_ = ~new_n5344_ & new_n5442_;
  assign new_n5713_ = ~new_n5438_ & new_n5712_;
  assign new_n5714_ = ~new_n5439_ & ~new_n5442_;
  assign new_n5715_ = ~new_n5713_ & ~new_n5714_;
  assign new_n5716_ = \quotient[37]  & ~new_n5715_;
  assign new_n5717_ = ~new_n5334_ & ~new_n5546_;
  assign new_n5718_ = ~new_n5545_ & new_n5717_;
  assign new_n5719_ = ~new_n5716_ & ~new_n5718_;
  assign new_n5720_ = ~\b[9]  & ~new_n5719_;
  assign new_n5721_ = ~new_n5353_ & new_n5437_;
  assign new_n5722_ = ~new_n5433_ & new_n5721_;
  assign new_n5723_ = ~new_n5434_ & ~new_n5437_;
  assign new_n5724_ = ~new_n5722_ & ~new_n5723_;
  assign new_n5725_ = \quotient[37]  & ~new_n5724_;
  assign new_n5726_ = ~new_n5343_ & ~new_n5546_;
  assign new_n5727_ = ~new_n5545_ & new_n5726_;
  assign new_n5728_ = ~new_n5725_ & ~new_n5727_;
  assign new_n5729_ = ~\b[8]  & ~new_n5728_;
  assign new_n5730_ = ~new_n5362_ & new_n5432_;
  assign new_n5731_ = ~new_n5428_ & new_n5730_;
  assign new_n5732_ = ~new_n5429_ & ~new_n5432_;
  assign new_n5733_ = ~new_n5731_ & ~new_n5732_;
  assign new_n5734_ = \quotient[37]  & ~new_n5733_;
  assign new_n5735_ = ~new_n5352_ & ~new_n5546_;
  assign new_n5736_ = ~new_n5545_ & new_n5735_;
  assign new_n5737_ = ~new_n5734_ & ~new_n5736_;
  assign new_n5738_ = ~\b[7]  & ~new_n5737_;
  assign new_n5739_ = ~new_n5371_ & new_n5427_;
  assign new_n5740_ = ~new_n5423_ & new_n5739_;
  assign new_n5741_ = ~new_n5424_ & ~new_n5427_;
  assign new_n5742_ = ~new_n5740_ & ~new_n5741_;
  assign new_n5743_ = \quotient[37]  & ~new_n5742_;
  assign new_n5744_ = ~new_n5361_ & ~new_n5546_;
  assign new_n5745_ = ~new_n5545_ & new_n5744_;
  assign new_n5746_ = ~new_n5743_ & ~new_n5745_;
  assign new_n5747_ = ~\b[6]  & ~new_n5746_;
  assign new_n5748_ = ~new_n5380_ & new_n5422_;
  assign new_n5749_ = ~new_n5418_ & new_n5748_;
  assign new_n5750_ = ~new_n5419_ & ~new_n5422_;
  assign new_n5751_ = ~new_n5749_ & ~new_n5750_;
  assign new_n5752_ = \quotient[37]  & ~new_n5751_;
  assign new_n5753_ = ~new_n5370_ & ~new_n5546_;
  assign new_n5754_ = ~new_n5545_ & new_n5753_;
  assign new_n5755_ = ~new_n5752_ & ~new_n5754_;
  assign new_n5756_ = ~\b[5]  & ~new_n5755_;
  assign new_n5757_ = ~new_n5388_ & new_n5417_;
  assign new_n5758_ = ~new_n5413_ & new_n5757_;
  assign new_n5759_ = ~new_n5414_ & ~new_n5417_;
  assign new_n5760_ = ~new_n5758_ & ~new_n5759_;
  assign new_n5761_ = \quotient[37]  & ~new_n5760_;
  assign new_n5762_ = ~new_n5379_ & ~new_n5546_;
  assign new_n5763_ = ~new_n5545_ & new_n5762_;
  assign new_n5764_ = ~new_n5761_ & ~new_n5763_;
  assign new_n5765_ = ~\b[4]  & ~new_n5764_;
  assign new_n5766_ = ~new_n5408_ & new_n5412_;
  assign new_n5767_ = ~new_n5407_ & new_n5766_;
  assign new_n5768_ = ~new_n5409_ & ~new_n5412_;
  assign new_n5769_ = ~new_n5767_ & ~new_n5768_;
  assign new_n5770_ = \quotient[37]  & ~new_n5769_;
  assign new_n5771_ = ~new_n5387_ & ~new_n5546_;
  assign new_n5772_ = ~new_n5545_ & new_n5771_;
  assign new_n5773_ = ~new_n5770_ & ~new_n5772_;
  assign new_n5774_ = ~\b[3]  & ~new_n5773_;
  assign new_n5775_ = ~new_n5404_ & new_n5406_;
  assign new_n5776_ = ~new_n5402_ & new_n5775_;
  assign new_n5777_ = ~new_n5407_ & ~new_n5776_;
  assign new_n5778_ = \quotient[37]  & new_n5777_;
  assign new_n5779_ = ~new_n5401_ & ~new_n5546_;
  assign new_n5780_ = ~new_n5545_ & new_n5779_;
  assign new_n5781_ = ~new_n5778_ & ~new_n5780_;
  assign new_n5782_ = ~\b[2]  & ~new_n5781_;
  assign new_n5783_ = \b[0]  & \quotient[37] ;
  assign new_n5784_ = \a[37]  & ~new_n5783_;
  assign new_n5785_ = new_n5406_ & \quotient[37] ;
  assign new_n5786_ = ~new_n5784_ & ~new_n5785_;
  assign new_n5787_ = \b[1]  & ~new_n5786_;
  assign new_n5788_ = ~\b[1]  & ~new_n5785_;
  assign new_n5789_ = ~new_n5784_ & new_n5788_;
  assign new_n5790_ = ~new_n5787_ & ~new_n5789_;
  assign new_n5791_ = ~\a[36]  & \b[0] ;
  assign new_n5792_ = ~new_n5790_ & ~new_n5791_;
  assign new_n5793_ = ~\b[1]  & ~new_n5786_;
  assign new_n5794_ = ~new_n5792_ & ~new_n5793_;
  assign new_n5795_ = \b[2]  & ~new_n5780_;
  assign new_n5796_ = ~new_n5778_ & new_n5795_;
  assign new_n5797_ = ~new_n5782_ & ~new_n5796_;
  assign new_n5798_ = ~new_n5794_ & new_n5797_;
  assign new_n5799_ = ~new_n5782_ & ~new_n5798_;
  assign new_n5800_ = \b[3]  & ~new_n5772_;
  assign new_n5801_ = ~new_n5770_ & new_n5800_;
  assign new_n5802_ = ~new_n5774_ & ~new_n5801_;
  assign new_n5803_ = ~new_n5799_ & new_n5802_;
  assign new_n5804_ = ~new_n5774_ & ~new_n5803_;
  assign new_n5805_ = \b[4]  & ~new_n5763_;
  assign new_n5806_ = ~new_n5761_ & new_n5805_;
  assign new_n5807_ = ~new_n5765_ & ~new_n5806_;
  assign new_n5808_ = ~new_n5804_ & new_n5807_;
  assign new_n5809_ = ~new_n5765_ & ~new_n5808_;
  assign new_n5810_ = \b[5]  & ~new_n5754_;
  assign new_n5811_ = ~new_n5752_ & new_n5810_;
  assign new_n5812_ = ~new_n5756_ & ~new_n5811_;
  assign new_n5813_ = ~new_n5809_ & new_n5812_;
  assign new_n5814_ = ~new_n5756_ & ~new_n5813_;
  assign new_n5815_ = \b[6]  & ~new_n5745_;
  assign new_n5816_ = ~new_n5743_ & new_n5815_;
  assign new_n5817_ = ~new_n5747_ & ~new_n5816_;
  assign new_n5818_ = ~new_n5814_ & new_n5817_;
  assign new_n5819_ = ~new_n5747_ & ~new_n5818_;
  assign new_n5820_ = \b[7]  & ~new_n5736_;
  assign new_n5821_ = ~new_n5734_ & new_n5820_;
  assign new_n5822_ = ~new_n5738_ & ~new_n5821_;
  assign new_n5823_ = ~new_n5819_ & new_n5822_;
  assign new_n5824_ = ~new_n5738_ & ~new_n5823_;
  assign new_n5825_ = \b[8]  & ~new_n5727_;
  assign new_n5826_ = ~new_n5725_ & new_n5825_;
  assign new_n5827_ = ~new_n5729_ & ~new_n5826_;
  assign new_n5828_ = ~new_n5824_ & new_n5827_;
  assign new_n5829_ = ~new_n5729_ & ~new_n5828_;
  assign new_n5830_ = \b[9]  & ~new_n5718_;
  assign new_n5831_ = ~new_n5716_ & new_n5830_;
  assign new_n5832_ = ~new_n5720_ & ~new_n5831_;
  assign new_n5833_ = ~new_n5829_ & new_n5832_;
  assign new_n5834_ = ~new_n5720_ & ~new_n5833_;
  assign new_n5835_ = \b[10]  & ~new_n5709_;
  assign new_n5836_ = ~new_n5707_ & new_n5835_;
  assign new_n5837_ = ~new_n5711_ & ~new_n5836_;
  assign new_n5838_ = ~new_n5834_ & new_n5837_;
  assign new_n5839_ = ~new_n5711_ & ~new_n5838_;
  assign new_n5840_ = \b[11]  & ~new_n5700_;
  assign new_n5841_ = ~new_n5698_ & new_n5840_;
  assign new_n5842_ = ~new_n5702_ & ~new_n5841_;
  assign new_n5843_ = ~new_n5839_ & new_n5842_;
  assign new_n5844_ = ~new_n5702_ & ~new_n5843_;
  assign new_n5845_ = \b[12]  & ~new_n5691_;
  assign new_n5846_ = ~new_n5689_ & new_n5845_;
  assign new_n5847_ = ~new_n5693_ & ~new_n5846_;
  assign new_n5848_ = ~new_n5844_ & new_n5847_;
  assign new_n5849_ = ~new_n5693_ & ~new_n5848_;
  assign new_n5850_ = \b[13]  & ~new_n5682_;
  assign new_n5851_ = ~new_n5680_ & new_n5850_;
  assign new_n5852_ = ~new_n5684_ & ~new_n5851_;
  assign new_n5853_ = ~new_n5849_ & new_n5852_;
  assign new_n5854_ = ~new_n5684_ & ~new_n5853_;
  assign new_n5855_ = \b[14]  & ~new_n5673_;
  assign new_n5856_ = ~new_n5671_ & new_n5855_;
  assign new_n5857_ = ~new_n5675_ & ~new_n5856_;
  assign new_n5858_ = ~new_n5854_ & new_n5857_;
  assign new_n5859_ = ~new_n5675_ & ~new_n5858_;
  assign new_n5860_ = \b[15]  & ~new_n5664_;
  assign new_n5861_ = ~new_n5662_ & new_n5860_;
  assign new_n5862_ = ~new_n5666_ & ~new_n5861_;
  assign new_n5863_ = ~new_n5859_ & new_n5862_;
  assign new_n5864_ = ~new_n5666_ & ~new_n5863_;
  assign new_n5865_ = \b[16]  & ~new_n5655_;
  assign new_n5866_ = ~new_n5653_ & new_n5865_;
  assign new_n5867_ = ~new_n5657_ & ~new_n5866_;
  assign new_n5868_ = ~new_n5864_ & new_n5867_;
  assign new_n5869_ = ~new_n5657_ & ~new_n5868_;
  assign new_n5870_ = \b[17]  & ~new_n5646_;
  assign new_n5871_ = ~new_n5644_ & new_n5870_;
  assign new_n5872_ = ~new_n5648_ & ~new_n5871_;
  assign new_n5873_ = ~new_n5869_ & new_n5872_;
  assign new_n5874_ = ~new_n5648_ & ~new_n5873_;
  assign new_n5875_ = \b[18]  & ~new_n5637_;
  assign new_n5876_ = ~new_n5635_ & new_n5875_;
  assign new_n5877_ = ~new_n5639_ & ~new_n5876_;
  assign new_n5878_ = ~new_n5874_ & new_n5877_;
  assign new_n5879_ = ~new_n5639_ & ~new_n5878_;
  assign new_n5880_ = \b[19]  & ~new_n5628_;
  assign new_n5881_ = ~new_n5626_ & new_n5880_;
  assign new_n5882_ = ~new_n5630_ & ~new_n5881_;
  assign new_n5883_ = ~new_n5879_ & new_n5882_;
  assign new_n5884_ = ~new_n5630_ & ~new_n5883_;
  assign new_n5885_ = \b[20]  & ~new_n5619_;
  assign new_n5886_ = ~new_n5617_ & new_n5885_;
  assign new_n5887_ = ~new_n5621_ & ~new_n5886_;
  assign new_n5888_ = ~new_n5884_ & new_n5887_;
  assign new_n5889_ = ~new_n5621_ & ~new_n5888_;
  assign new_n5890_ = \b[21]  & ~new_n5610_;
  assign new_n5891_ = ~new_n5608_ & new_n5890_;
  assign new_n5892_ = ~new_n5612_ & ~new_n5891_;
  assign new_n5893_ = ~new_n5889_ & new_n5892_;
  assign new_n5894_ = ~new_n5612_ & ~new_n5893_;
  assign new_n5895_ = \b[22]  & ~new_n5601_;
  assign new_n5896_ = ~new_n5599_ & new_n5895_;
  assign new_n5897_ = ~new_n5603_ & ~new_n5896_;
  assign new_n5898_ = ~new_n5894_ & new_n5897_;
  assign new_n5899_ = ~new_n5603_ & ~new_n5898_;
  assign new_n5900_ = \b[23]  & ~new_n5592_;
  assign new_n5901_ = ~new_n5590_ & new_n5900_;
  assign new_n5902_ = ~new_n5594_ & ~new_n5901_;
  assign new_n5903_ = ~new_n5899_ & new_n5902_;
  assign new_n5904_ = ~new_n5594_ & ~new_n5903_;
  assign new_n5905_ = \b[24]  & ~new_n5583_;
  assign new_n5906_ = ~new_n5581_ & new_n5905_;
  assign new_n5907_ = ~new_n5585_ & ~new_n5906_;
  assign new_n5908_ = ~new_n5904_ & new_n5907_;
  assign new_n5909_ = ~new_n5585_ & ~new_n5908_;
  assign new_n5910_ = \b[25]  & ~new_n5574_;
  assign new_n5911_ = ~new_n5572_ & new_n5910_;
  assign new_n5912_ = ~new_n5576_ & ~new_n5911_;
  assign new_n5913_ = ~new_n5909_ & new_n5912_;
  assign new_n5914_ = ~new_n5576_ & ~new_n5913_;
  assign new_n5915_ = \b[26]  & ~new_n5554_;
  assign new_n5916_ = ~new_n5552_ & new_n5915_;
  assign new_n5917_ = ~new_n5567_ & ~new_n5916_;
  assign new_n5918_ = ~new_n5914_ & new_n5917_;
  assign new_n5919_ = ~new_n5567_ & ~new_n5918_;
  assign new_n5920_ = \b[27]  & ~new_n5564_;
  assign new_n5921_ = ~new_n5562_ & new_n5920_;
  assign new_n5922_ = ~new_n5566_ & ~new_n5921_;
  assign new_n5923_ = ~new_n5919_ & new_n5922_;
  assign new_n5924_ = ~new_n5566_ & ~new_n5923_;
  assign new_n5925_ = new_n303_ & new_n317_;
  assign new_n5926_ = new_n288_ & new_n5925_;
  assign \quotient[36]  = ~new_n5924_ & new_n5926_;
  assign new_n5928_ = ~new_n5555_ & ~\quotient[36] ;
  assign new_n5929_ = ~new_n5576_ & new_n5917_;
  assign new_n5930_ = ~new_n5913_ & new_n5929_;
  assign new_n5931_ = ~new_n5914_ & ~new_n5917_;
  assign new_n5932_ = ~new_n5930_ & ~new_n5931_;
  assign new_n5933_ = new_n5926_ & ~new_n5932_;
  assign new_n5934_ = ~new_n5924_ & new_n5933_;
  assign new_n5935_ = ~new_n5928_ & ~new_n5934_;
  assign new_n5936_ = ~new_n5565_ & ~\quotient[36] ;
  assign new_n5937_ = ~new_n5567_ & new_n5922_;
  assign new_n5938_ = ~new_n5918_ & new_n5937_;
  assign new_n5939_ = ~new_n5919_ & ~new_n5922_;
  assign new_n5940_ = ~new_n5938_ & ~new_n5939_;
  assign new_n5941_ = \quotient[36]  & ~new_n5940_;
  assign new_n5942_ = ~new_n5936_ & ~new_n5941_;
  assign new_n5943_ = ~\b[28]  & ~new_n5942_;
  assign new_n5944_ = ~\b[27]  & ~new_n5935_;
  assign new_n5945_ = ~new_n5575_ & ~\quotient[36] ;
  assign new_n5946_ = ~new_n5585_ & new_n5912_;
  assign new_n5947_ = ~new_n5908_ & new_n5946_;
  assign new_n5948_ = ~new_n5909_ & ~new_n5912_;
  assign new_n5949_ = ~new_n5947_ & ~new_n5948_;
  assign new_n5950_ = new_n5926_ & ~new_n5949_;
  assign new_n5951_ = ~new_n5924_ & new_n5950_;
  assign new_n5952_ = ~new_n5945_ & ~new_n5951_;
  assign new_n5953_ = ~\b[26]  & ~new_n5952_;
  assign new_n5954_ = ~new_n5584_ & ~\quotient[36] ;
  assign new_n5955_ = ~new_n5594_ & new_n5907_;
  assign new_n5956_ = ~new_n5903_ & new_n5955_;
  assign new_n5957_ = ~new_n5904_ & ~new_n5907_;
  assign new_n5958_ = ~new_n5956_ & ~new_n5957_;
  assign new_n5959_ = new_n5926_ & ~new_n5958_;
  assign new_n5960_ = ~new_n5924_ & new_n5959_;
  assign new_n5961_ = ~new_n5954_ & ~new_n5960_;
  assign new_n5962_ = ~\b[25]  & ~new_n5961_;
  assign new_n5963_ = ~new_n5593_ & ~\quotient[36] ;
  assign new_n5964_ = ~new_n5603_ & new_n5902_;
  assign new_n5965_ = ~new_n5898_ & new_n5964_;
  assign new_n5966_ = ~new_n5899_ & ~new_n5902_;
  assign new_n5967_ = ~new_n5965_ & ~new_n5966_;
  assign new_n5968_ = new_n5926_ & ~new_n5967_;
  assign new_n5969_ = ~new_n5924_ & new_n5968_;
  assign new_n5970_ = ~new_n5963_ & ~new_n5969_;
  assign new_n5971_ = ~\b[24]  & ~new_n5970_;
  assign new_n5972_ = ~new_n5602_ & ~\quotient[36] ;
  assign new_n5973_ = ~new_n5612_ & new_n5897_;
  assign new_n5974_ = ~new_n5893_ & new_n5973_;
  assign new_n5975_ = ~new_n5894_ & ~new_n5897_;
  assign new_n5976_ = ~new_n5974_ & ~new_n5975_;
  assign new_n5977_ = new_n5926_ & ~new_n5976_;
  assign new_n5978_ = ~new_n5924_ & new_n5977_;
  assign new_n5979_ = ~new_n5972_ & ~new_n5978_;
  assign new_n5980_ = ~\b[23]  & ~new_n5979_;
  assign new_n5981_ = ~new_n5611_ & ~\quotient[36] ;
  assign new_n5982_ = ~new_n5621_ & new_n5892_;
  assign new_n5983_ = ~new_n5888_ & new_n5982_;
  assign new_n5984_ = ~new_n5889_ & ~new_n5892_;
  assign new_n5985_ = ~new_n5983_ & ~new_n5984_;
  assign new_n5986_ = new_n5926_ & ~new_n5985_;
  assign new_n5987_ = ~new_n5924_ & new_n5986_;
  assign new_n5988_ = ~new_n5981_ & ~new_n5987_;
  assign new_n5989_ = ~\b[22]  & ~new_n5988_;
  assign new_n5990_ = ~new_n5620_ & ~\quotient[36] ;
  assign new_n5991_ = ~new_n5630_ & new_n5887_;
  assign new_n5992_ = ~new_n5883_ & new_n5991_;
  assign new_n5993_ = ~new_n5884_ & ~new_n5887_;
  assign new_n5994_ = ~new_n5992_ & ~new_n5993_;
  assign new_n5995_ = new_n5926_ & ~new_n5994_;
  assign new_n5996_ = ~new_n5924_ & new_n5995_;
  assign new_n5997_ = ~new_n5990_ & ~new_n5996_;
  assign new_n5998_ = ~\b[21]  & ~new_n5997_;
  assign new_n5999_ = ~new_n5629_ & ~\quotient[36] ;
  assign new_n6000_ = ~new_n5639_ & new_n5882_;
  assign new_n6001_ = ~new_n5878_ & new_n6000_;
  assign new_n6002_ = ~new_n5879_ & ~new_n5882_;
  assign new_n6003_ = ~new_n6001_ & ~new_n6002_;
  assign new_n6004_ = new_n5926_ & ~new_n6003_;
  assign new_n6005_ = ~new_n5924_ & new_n6004_;
  assign new_n6006_ = ~new_n5999_ & ~new_n6005_;
  assign new_n6007_ = ~\b[20]  & ~new_n6006_;
  assign new_n6008_ = ~new_n5638_ & ~\quotient[36] ;
  assign new_n6009_ = ~new_n5648_ & new_n5877_;
  assign new_n6010_ = ~new_n5873_ & new_n6009_;
  assign new_n6011_ = ~new_n5874_ & ~new_n5877_;
  assign new_n6012_ = ~new_n6010_ & ~new_n6011_;
  assign new_n6013_ = new_n5926_ & ~new_n6012_;
  assign new_n6014_ = ~new_n5924_ & new_n6013_;
  assign new_n6015_ = ~new_n6008_ & ~new_n6014_;
  assign new_n6016_ = ~\b[19]  & ~new_n6015_;
  assign new_n6017_ = ~new_n5647_ & ~\quotient[36] ;
  assign new_n6018_ = ~new_n5657_ & new_n5872_;
  assign new_n6019_ = ~new_n5868_ & new_n6018_;
  assign new_n6020_ = ~new_n5869_ & ~new_n5872_;
  assign new_n6021_ = ~new_n6019_ & ~new_n6020_;
  assign new_n6022_ = new_n5926_ & ~new_n6021_;
  assign new_n6023_ = ~new_n5924_ & new_n6022_;
  assign new_n6024_ = ~new_n6017_ & ~new_n6023_;
  assign new_n6025_ = ~\b[18]  & ~new_n6024_;
  assign new_n6026_ = ~new_n5656_ & ~\quotient[36] ;
  assign new_n6027_ = ~new_n5666_ & new_n5867_;
  assign new_n6028_ = ~new_n5863_ & new_n6027_;
  assign new_n6029_ = ~new_n5864_ & ~new_n5867_;
  assign new_n6030_ = ~new_n6028_ & ~new_n6029_;
  assign new_n6031_ = new_n5926_ & ~new_n6030_;
  assign new_n6032_ = ~new_n5924_ & new_n6031_;
  assign new_n6033_ = ~new_n6026_ & ~new_n6032_;
  assign new_n6034_ = ~\b[17]  & ~new_n6033_;
  assign new_n6035_ = ~new_n5665_ & ~\quotient[36] ;
  assign new_n6036_ = ~new_n5675_ & new_n5862_;
  assign new_n6037_ = ~new_n5858_ & new_n6036_;
  assign new_n6038_ = ~new_n5859_ & ~new_n5862_;
  assign new_n6039_ = ~new_n6037_ & ~new_n6038_;
  assign new_n6040_ = new_n5926_ & ~new_n6039_;
  assign new_n6041_ = ~new_n5924_ & new_n6040_;
  assign new_n6042_ = ~new_n6035_ & ~new_n6041_;
  assign new_n6043_ = ~\b[16]  & ~new_n6042_;
  assign new_n6044_ = ~new_n5674_ & ~\quotient[36] ;
  assign new_n6045_ = ~new_n5684_ & new_n5857_;
  assign new_n6046_ = ~new_n5853_ & new_n6045_;
  assign new_n6047_ = ~new_n5854_ & ~new_n5857_;
  assign new_n6048_ = ~new_n6046_ & ~new_n6047_;
  assign new_n6049_ = new_n5926_ & ~new_n6048_;
  assign new_n6050_ = ~new_n5924_ & new_n6049_;
  assign new_n6051_ = ~new_n6044_ & ~new_n6050_;
  assign new_n6052_ = ~\b[15]  & ~new_n6051_;
  assign new_n6053_ = ~new_n5683_ & ~\quotient[36] ;
  assign new_n6054_ = ~new_n5693_ & new_n5852_;
  assign new_n6055_ = ~new_n5848_ & new_n6054_;
  assign new_n6056_ = ~new_n5849_ & ~new_n5852_;
  assign new_n6057_ = ~new_n6055_ & ~new_n6056_;
  assign new_n6058_ = new_n5926_ & ~new_n6057_;
  assign new_n6059_ = ~new_n5924_ & new_n6058_;
  assign new_n6060_ = ~new_n6053_ & ~new_n6059_;
  assign new_n6061_ = ~\b[14]  & ~new_n6060_;
  assign new_n6062_ = ~new_n5692_ & ~\quotient[36] ;
  assign new_n6063_ = ~new_n5702_ & new_n5847_;
  assign new_n6064_ = ~new_n5843_ & new_n6063_;
  assign new_n6065_ = ~new_n5844_ & ~new_n5847_;
  assign new_n6066_ = ~new_n6064_ & ~new_n6065_;
  assign new_n6067_ = new_n5926_ & ~new_n6066_;
  assign new_n6068_ = ~new_n5924_ & new_n6067_;
  assign new_n6069_ = ~new_n6062_ & ~new_n6068_;
  assign new_n6070_ = ~\b[13]  & ~new_n6069_;
  assign new_n6071_ = ~new_n5701_ & ~\quotient[36] ;
  assign new_n6072_ = ~new_n5711_ & new_n5842_;
  assign new_n6073_ = ~new_n5838_ & new_n6072_;
  assign new_n6074_ = ~new_n5839_ & ~new_n5842_;
  assign new_n6075_ = ~new_n6073_ & ~new_n6074_;
  assign new_n6076_ = new_n5926_ & ~new_n6075_;
  assign new_n6077_ = ~new_n5924_ & new_n6076_;
  assign new_n6078_ = ~new_n6071_ & ~new_n6077_;
  assign new_n6079_ = ~\b[12]  & ~new_n6078_;
  assign new_n6080_ = ~new_n5710_ & ~\quotient[36] ;
  assign new_n6081_ = ~new_n5720_ & new_n5837_;
  assign new_n6082_ = ~new_n5833_ & new_n6081_;
  assign new_n6083_ = ~new_n5834_ & ~new_n5837_;
  assign new_n6084_ = ~new_n6082_ & ~new_n6083_;
  assign new_n6085_ = new_n5926_ & ~new_n6084_;
  assign new_n6086_ = ~new_n5924_ & new_n6085_;
  assign new_n6087_ = ~new_n6080_ & ~new_n6086_;
  assign new_n6088_ = ~\b[11]  & ~new_n6087_;
  assign new_n6089_ = ~new_n5719_ & ~\quotient[36] ;
  assign new_n6090_ = ~new_n5729_ & new_n5832_;
  assign new_n6091_ = ~new_n5828_ & new_n6090_;
  assign new_n6092_ = ~new_n5829_ & ~new_n5832_;
  assign new_n6093_ = ~new_n6091_ & ~new_n6092_;
  assign new_n6094_ = new_n5926_ & ~new_n6093_;
  assign new_n6095_ = ~new_n5924_ & new_n6094_;
  assign new_n6096_ = ~new_n6089_ & ~new_n6095_;
  assign new_n6097_ = ~\b[10]  & ~new_n6096_;
  assign new_n6098_ = ~new_n5728_ & ~\quotient[36] ;
  assign new_n6099_ = ~new_n5738_ & new_n5827_;
  assign new_n6100_ = ~new_n5823_ & new_n6099_;
  assign new_n6101_ = ~new_n5824_ & ~new_n5827_;
  assign new_n6102_ = ~new_n6100_ & ~new_n6101_;
  assign new_n6103_ = new_n5926_ & ~new_n6102_;
  assign new_n6104_ = ~new_n5924_ & new_n6103_;
  assign new_n6105_ = ~new_n6098_ & ~new_n6104_;
  assign new_n6106_ = ~\b[9]  & ~new_n6105_;
  assign new_n6107_ = ~new_n5737_ & ~\quotient[36] ;
  assign new_n6108_ = ~new_n5747_ & new_n5822_;
  assign new_n6109_ = ~new_n5818_ & new_n6108_;
  assign new_n6110_ = ~new_n5819_ & ~new_n5822_;
  assign new_n6111_ = ~new_n6109_ & ~new_n6110_;
  assign new_n6112_ = new_n5926_ & ~new_n6111_;
  assign new_n6113_ = ~new_n5924_ & new_n6112_;
  assign new_n6114_ = ~new_n6107_ & ~new_n6113_;
  assign new_n6115_ = ~\b[8]  & ~new_n6114_;
  assign new_n6116_ = ~new_n5746_ & ~\quotient[36] ;
  assign new_n6117_ = ~new_n5756_ & new_n5817_;
  assign new_n6118_ = ~new_n5813_ & new_n6117_;
  assign new_n6119_ = ~new_n5814_ & ~new_n5817_;
  assign new_n6120_ = ~new_n6118_ & ~new_n6119_;
  assign new_n6121_ = new_n5926_ & ~new_n6120_;
  assign new_n6122_ = ~new_n5924_ & new_n6121_;
  assign new_n6123_ = ~new_n6116_ & ~new_n6122_;
  assign new_n6124_ = ~\b[7]  & ~new_n6123_;
  assign new_n6125_ = ~new_n5755_ & ~\quotient[36] ;
  assign new_n6126_ = ~new_n5765_ & new_n5812_;
  assign new_n6127_ = ~new_n5808_ & new_n6126_;
  assign new_n6128_ = ~new_n5809_ & ~new_n5812_;
  assign new_n6129_ = ~new_n6127_ & ~new_n6128_;
  assign new_n6130_ = new_n5926_ & ~new_n6129_;
  assign new_n6131_ = ~new_n5924_ & new_n6130_;
  assign new_n6132_ = ~new_n6125_ & ~new_n6131_;
  assign new_n6133_ = ~\b[6]  & ~new_n6132_;
  assign new_n6134_ = ~new_n5764_ & ~\quotient[36] ;
  assign new_n6135_ = ~new_n5774_ & new_n5807_;
  assign new_n6136_ = ~new_n5803_ & new_n6135_;
  assign new_n6137_ = ~new_n5804_ & ~new_n5807_;
  assign new_n6138_ = ~new_n6136_ & ~new_n6137_;
  assign new_n6139_ = new_n5926_ & ~new_n6138_;
  assign new_n6140_ = ~new_n5924_ & new_n6139_;
  assign new_n6141_ = ~new_n6134_ & ~new_n6140_;
  assign new_n6142_ = ~\b[5]  & ~new_n6141_;
  assign new_n6143_ = ~new_n5773_ & ~\quotient[36] ;
  assign new_n6144_ = ~new_n5782_ & new_n5802_;
  assign new_n6145_ = ~new_n5798_ & new_n6144_;
  assign new_n6146_ = ~new_n5799_ & ~new_n5802_;
  assign new_n6147_ = ~new_n6145_ & ~new_n6146_;
  assign new_n6148_ = new_n5926_ & ~new_n6147_;
  assign new_n6149_ = ~new_n5924_ & new_n6148_;
  assign new_n6150_ = ~new_n6143_ & ~new_n6149_;
  assign new_n6151_ = ~\b[4]  & ~new_n6150_;
  assign new_n6152_ = ~new_n5781_ & ~\quotient[36] ;
  assign new_n6153_ = ~new_n5793_ & new_n5797_;
  assign new_n6154_ = ~new_n5792_ & new_n6153_;
  assign new_n6155_ = ~new_n5794_ & ~new_n5797_;
  assign new_n6156_ = ~new_n6154_ & ~new_n6155_;
  assign new_n6157_ = new_n5926_ & ~new_n6156_;
  assign new_n6158_ = ~new_n5924_ & new_n6157_;
  assign new_n6159_ = ~new_n6152_ & ~new_n6158_;
  assign new_n6160_ = ~\b[3]  & ~new_n6159_;
  assign new_n6161_ = ~new_n5786_ & ~\quotient[36] ;
  assign new_n6162_ = ~new_n5789_ & new_n5791_;
  assign new_n6163_ = ~new_n5787_ & new_n6162_;
  assign new_n6164_ = new_n5926_ & ~new_n6163_;
  assign new_n6165_ = ~new_n5792_ & new_n6164_;
  assign new_n6166_ = ~new_n5924_ & new_n6165_;
  assign new_n6167_ = ~new_n6161_ & ~new_n6166_;
  assign new_n6168_ = ~\b[2]  & ~new_n6167_;
  assign new_n6169_ = \b[0]  & ~\b[28] ;
  assign new_n6170_ = new_n373_ & new_n6169_;
  assign new_n6171_ = new_n423_ & new_n6170_;
  assign new_n6172_ = new_n408_ & new_n6171_;
  assign new_n6173_ = ~new_n5924_ & new_n6172_;
  assign new_n6174_ = \a[36]  & ~new_n6173_;
  assign new_n6175_ = new_n316_ & new_n5791_;
  assign new_n6176_ = new_n341_ & new_n6175_;
  assign new_n6177_ = new_n338_ & new_n6176_;
  assign new_n6178_ = ~new_n5924_ & new_n6177_;
  assign new_n6179_ = ~new_n6174_ & ~new_n6178_;
  assign new_n6180_ = \b[1]  & ~new_n6179_;
  assign new_n6181_ = ~\b[1]  & ~new_n6178_;
  assign new_n6182_ = ~new_n6174_ & new_n6181_;
  assign new_n6183_ = ~new_n6180_ & ~new_n6182_;
  assign new_n6184_ = ~\a[35]  & \b[0] ;
  assign new_n6185_ = ~new_n6183_ & ~new_n6184_;
  assign new_n6186_ = ~\b[1]  & ~new_n6179_;
  assign new_n6187_ = ~new_n6185_ & ~new_n6186_;
  assign new_n6188_ = \b[2]  & ~new_n6166_;
  assign new_n6189_ = ~new_n6161_ & new_n6188_;
  assign new_n6190_ = ~new_n6168_ & ~new_n6189_;
  assign new_n6191_ = ~new_n6187_ & new_n6190_;
  assign new_n6192_ = ~new_n6168_ & ~new_n6191_;
  assign new_n6193_ = \b[3]  & ~new_n6158_;
  assign new_n6194_ = ~new_n6152_ & new_n6193_;
  assign new_n6195_ = ~new_n6160_ & ~new_n6194_;
  assign new_n6196_ = ~new_n6192_ & new_n6195_;
  assign new_n6197_ = ~new_n6160_ & ~new_n6196_;
  assign new_n6198_ = \b[4]  & ~new_n6149_;
  assign new_n6199_ = ~new_n6143_ & new_n6198_;
  assign new_n6200_ = ~new_n6151_ & ~new_n6199_;
  assign new_n6201_ = ~new_n6197_ & new_n6200_;
  assign new_n6202_ = ~new_n6151_ & ~new_n6201_;
  assign new_n6203_ = \b[5]  & ~new_n6140_;
  assign new_n6204_ = ~new_n6134_ & new_n6203_;
  assign new_n6205_ = ~new_n6142_ & ~new_n6204_;
  assign new_n6206_ = ~new_n6202_ & new_n6205_;
  assign new_n6207_ = ~new_n6142_ & ~new_n6206_;
  assign new_n6208_ = \b[6]  & ~new_n6131_;
  assign new_n6209_ = ~new_n6125_ & new_n6208_;
  assign new_n6210_ = ~new_n6133_ & ~new_n6209_;
  assign new_n6211_ = ~new_n6207_ & new_n6210_;
  assign new_n6212_ = ~new_n6133_ & ~new_n6211_;
  assign new_n6213_ = \b[7]  & ~new_n6122_;
  assign new_n6214_ = ~new_n6116_ & new_n6213_;
  assign new_n6215_ = ~new_n6124_ & ~new_n6214_;
  assign new_n6216_ = ~new_n6212_ & new_n6215_;
  assign new_n6217_ = ~new_n6124_ & ~new_n6216_;
  assign new_n6218_ = \b[8]  & ~new_n6113_;
  assign new_n6219_ = ~new_n6107_ & new_n6218_;
  assign new_n6220_ = ~new_n6115_ & ~new_n6219_;
  assign new_n6221_ = ~new_n6217_ & new_n6220_;
  assign new_n6222_ = ~new_n6115_ & ~new_n6221_;
  assign new_n6223_ = \b[9]  & ~new_n6104_;
  assign new_n6224_ = ~new_n6098_ & new_n6223_;
  assign new_n6225_ = ~new_n6106_ & ~new_n6224_;
  assign new_n6226_ = ~new_n6222_ & new_n6225_;
  assign new_n6227_ = ~new_n6106_ & ~new_n6226_;
  assign new_n6228_ = \b[10]  & ~new_n6095_;
  assign new_n6229_ = ~new_n6089_ & new_n6228_;
  assign new_n6230_ = ~new_n6097_ & ~new_n6229_;
  assign new_n6231_ = ~new_n6227_ & new_n6230_;
  assign new_n6232_ = ~new_n6097_ & ~new_n6231_;
  assign new_n6233_ = \b[11]  & ~new_n6086_;
  assign new_n6234_ = ~new_n6080_ & new_n6233_;
  assign new_n6235_ = ~new_n6088_ & ~new_n6234_;
  assign new_n6236_ = ~new_n6232_ & new_n6235_;
  assign new_n6237_ = ~new_n6088_ & ~new_n6236_;
  assign new_n6238_ = \b[12]  & ~new_n6077_;
  assign new_n6239_ = ~new_n6071_ & new_n6238_;
  assign new_n6240_ = ~new_n6079_ & ~new_n6239_;
  assign new_n6241_ = ~new_n6237_ & new_n6240_;
  assign new_n6242_ = ~new_n6079_ & ~new_n6241_;
  assign new_n6243_ = \b[13]  & ~new_n6068_;
  assign new_n6244_ = ~new_n6062_ & new_n6243_;
  assign new_n6245_ = ~new_n6070_ & ~new_n6244_;
  assign new_n6246_ = ~new_n6242_ & new_n6245_;
  assign new_n6247_ = ~new_n6070_ & ~new_n6246_;
  assign new_n6248_ = \b[14]  & ~new_n6059_;
  assign new_n6249_ = ~new_n6053_ & new_n6248_;
  assign new_n6250_ = ~new_n6061_ & ~new_n6249_;
  assign new_n6251_ = ~new_n6247_ & new_n6250_;
  assign new_n6252_ = ~new_n6061_ & ~new_n6251_;
  assign new_n6253_ = \b[15]  & ~new_n6050_;
  assign new_n6254_ = ~new_n6044_ & new_n6253_;
  assign new_n6255_ = ~new_n6052_ & ~new_n6254_;
  assign new_n6256_ = ~new_n6252_ & new_n6255_;
  assign new_n6257_ = ~new_n6052_ & ~new_n6256_;
  assign new_n6258_ = \b[16]  & ~new_n6041_;
  assign new_n6259_ = ~new_n6035_ & new_n6258_;
  assign new_n6260_ = ~new_n6043_ & ~new_n6259_;
  assign new_n6261_ = ~new_n6257_ & new_n6260_;
  assign new_n6262_ = ~new_n6043_ & ~new_n6261_;
  assign new_n6263_ = \b[17]  & ~new_n6032_;
  assign new_n6264_ = ~new_n6026_ & new_n6263_;
  assign new_n6265_ = ~new_n6034_ & ~new_n6264_;
  assign new_n6266_ = ~new_n6262_ & new_n6265_;
  assign new_n6267_ = ~new_n6034_ & ~new_n6266_;
  assign new_n6268_ = \b[18]  & ~new_n6023_;
  assign new_n6269_ = ~new_n6017_ & new_n6268_;
  assign new_n6270_ = ~new_n6025_ & ~new_n6269_;
  assign new_n6271_ = ~new_n6267_ & new_n6270_;
  assign new_n6272_ = ~new_n6025_ & ~new_n6271_;
  assign new_n6273_ = \b[19]  & ~new_n6014_;
  assign new_n6274_ = ~new_n6008_ & new_n6273_;
  assign new_n6275_ = ~new_n6016_ & ~new_n6274_;
  assign new_n6276_ = ~new_n6272_ & new_n6275_;
  assign new_n6277_ = ~new_n6016_ & ~new_n6276_;
  assign new_n6278_ = \b[20]  & ~new_n6005_;
  assign new_n6279_ = ~new_n5999_ & new_n6278_;
  assign new_n6280_ = ~new_n6007_ & ~new_n6279_;
  assign new_n6281_ = ~new_n6277_ & new_n6280_;
  assign new_n6282_ = ~new_n6007_ & ~new_n6281_;
  assign new_n6283_ = \b[21]  & ~new_n5996_;
  assign new_n6284_ = ~new_n5990_ & new_n6283_;
  assign new_n6285_ = ~new_n5998_ & ~new_n6284_;
  assign new_n6286_ = ~new_n6282_ & new_n6285_;
  assign new_n6287_ = ~new_n5998_ & ~new_n6286_;
  assign new_n6288_ = \b[22]  & ~new_n5987_;
  assign new_n6289_ = ~new_n5981_ & new_n6288_;
  assign new_n6290_ = ~new_n5989_ & ~new_n6289_;
  assign new_n6291_ = ~new_n6287_ & new_n6290_;
  assign new_n6292_ = ~new_n5989_ & ~new_n6291_;
  assign new_n6293_ = \b[23]  & ~new_n5978_;
  assign new_n6294_ = ~new_n5972_ & new_n6293_;
  assign new_n6295_ = ~new_n5980_ & ~new_n6294_;
  assign new_n6296_ = ~new_n6292_ & new_n6295_;
  assign new_n6297_ = ~new_n5980_ & ~new_n6296_;
  assign new_n6298_ = \b[24]  & ~new_n5969_;
  assign new_n6299_ = ~new_n5963_ & new_n6298_;
  assign new_n6300_ = ~new_n5971_ & ~new_n6299_;
  assign new_n6301_ = ~new_n6297_ & new_n6300_;
  assign new_n6302_ = ~new_n5971_ & ~new_n6301_;
  assign new_n6303_ = \b[25]  & ~new_n5960_;
  assign new_n6304_ = ~new_n5954_ & new_n6303_;
  assign new_n6305_ = ~new_n5962_ & ~new_n6304_;
  assign new_n6306_ = ~new_n6302_ & new_n6305_;
  assign new_n6307_ = ~new_n5962_ & ~new_n6306_;
  assign new_n6308_ = \b[26]  & ~new_n5951_;
  assign new_n6309_ = ~new_n5945_ & new_n6308_;
  assign new_n6310_ = ~new_n5953_ & ~new_n6309_;
  assign new_n6311_ = ~new_n6307_ & new_n6310_;
  assign new_n6312_ = ~new_n5953_ & ~new_n6311_;
  assign new_n6313_ = \b[27]  & ~new_n5934_;
  assign new_n6314_ = ~new_n5928_ & new_n6313_;
  assign new_n6315_ = ~new_n5944_ & ~new_n6314_;
  assign new_n6316_ = ~new_n6312_ & new_n6315_;
  assign new_n6317_ = ~new_n5944_ & ~new_n6316_;
  assign new_n6318_ = \b[28]  & ~new_n5936_;
  assign new_n6319_ = ~new_n5941_ & new_n6318_;
  assign new_n6320_ = ~new_n5943_ & ~new_n6319_;
  assign new_n6321_ = ~new_n6317_ & new_n6320_;
  assign new_n6322_ = ~new_n5943_ & ~new_n6321_;
  assign new_n6323_ = new_n588_ & new_n598_;
  assign new_n6324_ = new_n595_ & new_n6323_;
  assign \quotient[35]  = ~new_n6322_ & new_n6324_;
  assign new_n6326_ = ~new_n5935_ & ~\quotient[35] ;
  assign new_n6327_ = ~new_n5953_ & new_n6315_;
  assign new_n6328_ = ~new_n6311_ & new_n6327_;
  assign new_n6329_ = ~new_n6312_ & ~new_n6315_;
  assign new_n6330_ = ~new_n6328_ & ~new_n6329_;
  assign new_n6331_ = new_n6324_ & ~new_n6330_;
  assign new_n6332_ = ~new_n6322_ & new_n6331_;
  assign new_n6333_ = ~new_n6326_ & ~new_n6332_;
  assign new_n6334_ = ~\b[28]  & ~new_n6333_;
  assign new_n6335_ = ~new_n5952_ & ~\quotient[35] ;
  assign new_n6336_ = ~new_n5962_ & new_n6310_;
  assign new_n6337_ = ~new_n6306_ & new_n6336_;
  assign new_n6338_ = ~new_n6307_ & ~new_n6310_;
  assign new_n6339_ = ~new_n6337_ & ~new_n6338_;
  assign new_n6340_ = new_n6324_ & ~new_n6339_;
  assign new_n6341_ = ~new_n6322_ & new_n6340_;
  assign new_n6342_ = ~new_n6335_ & ~new_n6341_;
  assign new_n6343_ = ~\b[27]  & ~new_n6342_;
  assign new_n6344_ = ~new_n5961_ & ~\quotient[35] ;
  assign new_n6345_ = ~new_n5971_ & new_n6305_;
  assign new_n6346_ = ~new_n6301_ & new_n6345_;
  assign new_n6347_ = ~new_n6302_ & ~new_n6305_;
  assign new_n6348_ = ~new_n6346_ & ~new_n6347_;
  assign new_n6349_ = new_n6324_ & ~new_n6348_;
  assign new_n6350_ = ~new_n6322_ & new_n6349_;
  assign new_n6351_ = ~new_n6344_ & ~new_n6350_;
  assign new_n6352_ = ~\b[26]  & ~new_n6351_;
  assign new_n6353_ = ~new_n5970_ & ~\quotient[35] ;
  assign new_n6354_ = ~new_n5980_ & new_n6300_;
  assign new_n6355_ = ~new_n6296_ & new_n6354_;
  assign new_n6356_ = ~new_n6297_ & ~new_n6300_;
  assign new_n6357_ = ~new_n6355_ & ~new_n6356_;
  assign new_n6358_ = new_n6324_ & ~new_n6357_;
  assign new_n6359_ = ~new_n6322_ & new_n6358_;
  assign new_n6360_ = ~new_n6353_ & ~new_n6359_;
  assign new_n6361_ = ~\b[25]  & ~new_n6360_;
  assign new_n6362_ = ~new_n5979_ & ~\quotient[35] ;
  assign new_n6363_ = ~new_n5989_ & new_n6295_;
  assign new_n6364_ = ~new_n6291_ & new_n6363_;
  assign new_n6365_ = ~new_n6292_ & ~new_n6295_;
  assign new_n6366_ = ~new_n6364_ & ~new_n6365_;
  assign new_n6367_ = new_n6324_ & ~new_n6366_;
  assign new_n6368_ = ~new_n6322_ & new_n6367_;
  assign new_n6369_ = ~new_n6362_ & ~new_n6368_;
  assign new_n6370_ = ~\b[24]  & ~new_n6369_;
  assign new_n6371_ = ~new_n5988_ & ~\quotient[35] ;
  assign new_n6372_ = ~new_n5998_ & new_n6290_;
  assign new_n6373_ = ~new_n6286_ & new_n6372_;
  assign new_n6374_ = ~new_n6287_ & ~new_n6290_;
  assign new_n6375_ = ~new_n6373_ & ~new_n6374_;
  assign new_n6376_ = new_n6324_ & ~new_n6375_;
  assign new_n6377_ = ~new_n6322_ & new_n6376_;
  assign new_n6378_ = ~new_n6371_ & ~new_n6377_;
  assign new_n6379_ = ~\b[23]  & ~new_n6378_;
  assign new_n6380_ = ~new_n5997_ & ~\quotient[35] ;
  assign new_n6381_ = ~new_n6007_ & new_n6285_;
  assign new_n6382_ = ~new_n6281_ & new_n6381_;
  assign new_n6383_ = ~new_n6282_ & ~new_n6285_;
  assign new_n6384_ = ~new_n6382_ & ~new_n6383_;
  assign new_n6385_ = new_n6324_ & ~new_n6384_;
  assign new_n6386_ = ~new_n6322_ & new_n6385_;
  assign new_n6387_ = ~new_n6380_ & ~new_n6386_;
  assign new_n6388_ = ~\b[22]  & ~new_n6387_;
  assign new_n6389_ = ~new_n6006_ & ~\quotient[35] ;
  assign new_n6390_ = ~new_n6016_ & new_n6280_;
  assign new_n6391_ = ~new_n6276_ & new_n6390_;
  assign new_n6392_ = ~new_n6277_ & ~new_n6280_;
  assign new_n6393_ = ~new_n6391_ & ~new_n6392_;
  assign new_n6394_ = new_n6324_ & ~new_n6393_;
  assign new_n6395_ = ~new_n6322_ & new_n6394_;
  assign new_n6396_ = ~new_n6389_ & ~new_n6395_;
  assign new_n6397_ = ~\b[21]  & ~new_n6396_;
  assign new_n6398_ = ~new_n6015_ & ~\quotient[35] ;
  assign new_n6399_ = ~new_n6025_ & new_n6275_;
  assign new_n6400_ = ~new_n6271_ & new_n6399_;
  assign new_n6401_ = ~new_n6272_ & ~new_n6275_;
  assign new_n6402_ = ~new_n6400_ & ~new_n6401_;
  assign new_n6403_ = new_n6324_ & ~new_n6402_;
  assign new_n6404_ = ~new_n6322_ & new_n6403_;
  assign new_n6405_ = ~new_n6398_ & ~new_n6404_;
  assign new_n6406_ = ~\b[20]  & ~new_n6405_;
  assign new_n6407_ = ~new_n6024_ & ~\quotient[35] ;
  assign new_n6408_ = ~new_n6034_ & new_n6270_;
  assign new_n6409_ = ~new_n6266_ & new_n6408_;
  assign new_n6410_ = ~new_n6267_ & ~new_n6270_;
  assign new_n6411_ = ~new_n6409_ & ~new_n6410_;
  assign new_n6412_ = new_n6324_ & ~new_n6411_;
  assign new_n6413_ = ~new_n6322_ & new_n6412_;
  assign new_n6414_ = ~new_n6407_ & ~new_n6413_;
  assign new_n6415_ = ~\b[19]  & ~new_n6414_;
  assign new_n6416_ = ~new_n6033_ & ~\quotient[35] ;
  assign new_n6417_ = ~new_n6043_ & new_n6265_;
  assign new_n6418_ = ~new_n6261_ & new_n6417_;
  assign new_n6419_ = ~new_n6262_ & ~new_n6265_;
  assign new_n6420_ = ~new_n6418_ & ~new_n6419_;
  assign new_n6421_ = new_n6324_ & ~new_n6420_;
  assign new_n6422_ = ~new_n6322_ & new_n6421_;
  assign new_n6423_ = ~new_n6416_ & ~new_n6422_;
  assign new_n6424_ = ~\b[18]  & ~new_n6423_;
  assign new_n6425_ = ~new_n6042_ & ~\quotient[35] ;
  assign new_n6426_ = ~new_n6052_ & new_n6260_;
  assign new_n6427_ = ~new_n6256_ & new_n6426_;
  assign new_n6428_ = ~new_n6257_ & ~new_n6260_;
  assign new_n6429_ = ~new_n6427_ & ~new_n6428_;
  assign new_n6430_ = new_n6324_ & ~new_n6429_;
  assign new_n6431_ = ~new_n6322_ & new_n6430_;
  assign new_n6432_ = ~new_n6425_ & ~new_n6431_;
  assign new_n6433_ = ~\b[17]  & ~new_n6432_;
  assign new_n6434_ = ~new_n6051_ & ~\quotient[35] ;
  assign new_n6435_ = ~new_n6061_ & new_n6255_;
  assign new_n6436_ = ~new_n6251_ & new_n6435_;
  assign new_n6437_ = ~new_n6252_ & ~new_n6255_;
  assign new_n6438_ = ~new_n6436_ & ~new_n6437_;
  assign new_n6439_ = new_n6324_ & ~new_n6438_;
  assign new_n6440_ = ~new_n6322_ & new_n6439_;
  assign new_n6441_ = ~new_n6434_ & ~new_n6440_;
  assign new_n6442_ = ~\b[16]  & ~new_n6441_;
  assign new_n6443_ = ~new_n6060_ & ~\quotient[35] ;
  assign new_n6444_ = ~new_n6070_ & new_n6250_;
  assign new_n6445_ = ~new_n6246_ & new_n6444_;
  assign new_n6446_ = ~new_n6247_ & ~new_n6250_;
  assign new_n6447_ = ~new_n6445_ & ~new_n6446_;
  assign new_n6448_ = new_n6324_ & ~new_n6447_;
  assign new_n6449_ = ~new_n6322_ & new_n6448_;
  assign new_n6450_ = ~new_n6443_ & ~new_n6449_;
  assign new_n6451_ = ~\b[15]  & ~new_n6450_;
  assign new_n6452_ = ~new_n6069_ & ~\quotient[35] ;
  assign new_n6453_ = ~new_n6079_ & new_n6245_;
  assign new_n6454_ = ~new_n6241_ & new_n6453_;
  assign new_n6455_ = ~new_n6242_ & ~new_n6245_;
  assign new_n6456_ = ~new_n6454_ & ~new_n6455_;
  assign new_n6457_ = new_n6324_ & ~new_n6456_;
  assign new_n6458_ = ~new_n6322_ & new_n6457_;
  assign new_n6459_ = ~new_n6452_ & ~new_n6458_;
  assign new_n6460_ = ~\b[14]  & ~new_n6459_;
  assign new_n6461_ = ~new_n6078_ & ~\quotient[35] ;
  assign new_n6462_ = ~new_n6088_ & new_n6240_;
  assign new_n6463_ = ~new_n6236_ & new_n6462_;
  assign new_n6464_ = ~new_n6237_ & ~new_n6240_;
  assign new_n6465_ = ~new_n6463_ & ~new_n6464_;
  assign new_n6466_ = new_n6324_ & ~new_n6465_;
  assign new_n6467_ = ~new_n6322_ & new_n6466_;
  assign new_n6468_ = ~new_n6461_ & ~new_n6467_;
  assign new_n6469_ = ~\b[13]  & ~new_n6468_;
  assign new_n6470_ = ~new_n6087_ & ~\quotient[35] ;
  assign new_n6471_ = ~new_n6097_ & new_n6235_;
  assign new_n6472_ = ~new_n6231_ & new_n6471_;
  assign new_n6473_ = ~new_n6232_ & ~new_n6235_;
  assign new_n6474_ = ~new_n6472_ & ~new_n6473_;
  assign new_n6475_ = new_n6324_ & ~new_n6474_;
  assign new_n6476_ = ~new_n6322_ & new_n6475_;
  assign new_n6477_ = ~new_n6470_ & ~new_n6476_;
  assign new_n6478_ = ~\b[12]  & ~new_n6477_;
  assign new_n6479_ = ~new_n6096_ & ~\quotient[35] ;
  assign new_n6480_ = ~new_n6106_ & new_n6230_;
  assign new_n6481_ = ~new_n6226_ & new_n6480_;
  assign new_n6482_ = ~new_n6227_ & ~new_n6230_;
  assign new_n6483_ = ~new_n6481_ & ~new_n6482_;
  assign new_n6484_ = new_n6324_ & ~new_n6483_;
  assign new_n6485_ = ~new_n6322_ & new_n6484_;
  assign new_n6486_ = ~new_n6479_ & ~new_n6485_;
  assign new_n6487_ = ~\b[11]  & ~new_n6486_;
  assign new_n6488_ = ~new_n6105_ & ~\quotient[35] ;
  assign new_n6489_ = ~new_n6115_ & new_n6225_;
  assign new_n6490_ = ~new_n6221_ & new_n6489_;
  assign new_n6491_ = ~new_n6222_ & ~new_n6225_;
  assign new_n6492_ = ~new_n6490_ & ~new_n6491_;
  assign new_n6493_ = new_n6324_ & ~new_n6492_;
  assign new_n6494_ = ~new_n6322_ & new_n6493_;
  assign new_n6495_ = ~new_n6488_ & ~new_n6494_;
  assign new_n6496_ = ~\b[10]  & ~new_n6495_;
  assign new_n6497_ = ~new_n6114_ & ~\quotient[35] ;
  assign new_n6498_ = ~new_n6124_ & new_n6220_;
  assign new_n6499_ = ~new_n6216_ & new_n6498_;
  assign new_n6500_ = ~new_n6217_ & ~new_n6220_;
  assign new_n6501_ = ~new_n6499_ & ~new_n6500_;
  assign new_n6502_ = new_n6324_ & ~new_n6501_;
  assign new_n6503_ = ~new_n6322_ & new_n6502_;
  assign new_n6504_ = ~new_n6497_ & ~new_n6503_;
  assign new_n6505_ = ~\b[9]  & ~new_n6504_;
  assign new_n6506_ = ~new_n6123_ & ~\quotient[35] ;
  assign new_n6507_ = ~new_n6133_ & new_n6215_;
  assign new_n6508_ = ~new_n6211_ & new_n6507_;
  assign new_n6509_ = ~new_n6212_ & ~new_n6215_;
  assign new_n6510_ = ~new_n6508_ & ~new_n6509_;
  assign new_n6511_ = new_n6324_ & ~new_n6510_;
  assign new_n6512_ = ~new_n6322_ & new_n6511_;
  assign new_n6513_ = ~new_n6506_ & ~new_n6512_;
  assign new_n6514_ = ~\b[8]  & ~new_n6513_;
  assign new_n6515_ = ~new_n6132_ & ~\quotient[35] ;
  assign new_n6516_ = ~new_n6142_ & new_n6210_;
  assign new_n6517_ = ~new_n6206_ & new_n6516_;
  assign new_n6518_ = ~new_n6207_ & ~new_n6210_;
  assign new_n6519_ = ~new_n6517_ & ~new_n6518_;
  assign new_n6520_ = new_n6324_ & ~new_n6519_;
  assign new_n6521_ = ~new_n6322_ & new_n6520_;
  assign new_n6522_ = ~new_n6515_ & ~new_n6521_;
  assign new_n6523_ = ~\b[7]  & ~new_n6522_;
  assign new_n6524_ = ~new_n6141_ & ~\quotient[35] ;
  assign new_n6525_ = ~new_n6151_ & new_n6205_;
  assign new_n6526_ = ~new_n6201_ & new_n6525_;
  assign new_n6527_ = ~new_n6202_ & ~new_n6205_;
  assign new_n6528_ = ~new_n6526_ & ~new_n6527_;
  assign new_n6529_ = new_n6324_ & ~new_n6528_;
  assign new_n6530_ = ~new_n6322_ & new_n6529_;
  assign new_n6531_ = ~new_n6524_ & ~new_n6530_;
  assign new_n6532_ = ~\b[6]  & ~new_n6531_;
  assign new_n6533_ = ~new_n6150_ & ~\quotient[35] ;
  assign new_n6534_ = ~new_n6160_ & new_n6200_;
  assign new_n6535_ = ~new_n6196_ & new_n6534_;
  assign new_n6536_ = ~new_n6197_ & ~new_n6200_;
  assign new_n6537_ = ~new_n6535_ & ~new_n6536_;
  assign new_n6538_ = new_n6324_ & ~new_n6537_;
  assign new_n6539_ = ~new_n6322_ & new_n6538_;
  assign new_n6540_ = ~new_n6533_ & ~new_n6539_;
  assign new_n6541_ = ~\b[5]  & ~new_n6540_;
  assign new_n6542_ = ~new_n6159_ & ~\quotient[35] ;
  assign new_n6543_ = ~new_n6168_ & new_n6195_;
  assign new_n6544_ = ~new_n6191_ & new_n6543_;
  assign new_n6545_ = ~new_n6192_ & ~new_n6195_;
  assign new_n6546_ = ~new_n6544_ & ~new_n6545_;
  assign new_n6547_ = new_n6324_ & ~new_n6546_;
  assign new_n6548_ = ~new_n6322_ & new_n6547_;
  assign new_n6549_ = ~new_n6542_ & ~new_n6548_;
  assign new_n6550_ = ~\b[4]  & ~new_n6549_;
  assign new_n6551_ = ~new_n6167_ & ~\quotient[35] ;
  assign new_n6552_ = ~new_n6186_ & new_n6190_;
  assign new_n6553_ = ~new_n6185_ & new_n6552_;
  assign new_n6554_ = ~new_n6187_ & ~new_n6190_;
  assign new_n6555_ = ~new_n6553_ & ~new_n6554_;
  assign new_n6556_ = new_n6324_ & ~new_n6555_;
  assign new_n6557_ = ~new_n6322_ & new_n6556_;
  assign new_n6558_ = ~new_n6551_ & ~new_n6557_;
  assign new_n6559_ = ~\b[3]  & ~new_n6558_;
  assign new_n6560_ = ~new_n6179_ & ~\quotient[35] ;
  assign new_n6561_ = ~new_n6182_ & new_n6184_;
  assign new_n6562_ = ~new_n6180_ & new_n6561_;
  assign new_n6563_ = new_n6324_ & ~new_n6562_;
  assign new_n6564_ = ~new_n6185_ & new_n6563_;
  assign new_n6565_ = ~new_n6322_ & new_n6564_;
  assign new_n6566_ = ~new_n6560_ & ~new_n6565_;
  assign new_n6567_ = ~\b[2]  & ~new_n6566_;
  assign new_n6568_ = \b[0]  & ~\b[29] ;
  assign new_n6569_ = new_n315_ & new_n6568_;
  assign new_n6570_ = new_n313_ & new_n6569_;
  assign new_n6571_ = new_n303_ & new_n6570_;
  assign new_n6572_ = new_n288_ & new_n6571_;
  assign new_n6573_ = ~new_n6322_ & new_n6572_;
  assign new_n6574_ = \a[35]  & ~new_n6573_;
  assign new_n6575_ = new_n373_ & new_n6184_;
  assign new_n6576_ = new_n423_ & new_n6575_;
  assign new_n6577_ = new_n408_ & new_n6576_;
  assign new_n6578_ = ~new_n6322_ & new_n6577_;
  assign new_n6579_ = ~new_n6574_ & ~new_n6578_;
  assign new_n6580_ = \b[1]  & ~new_n6579_;
  assign new_n6581_ = ~\b[1]  & ~new_n6578_;
  assign new_n6582_ = ~new_n6574_ & new_n6581_;
  assign new_n6583_ = ~new_n6580_ & ~new_n6582_;
  assign new_n6584_ = ~\a[34]  & \b[0] ;
  assign new_n6585_ = ~new_n6583_ & ~new_n6584_;
  assign new_n6586_ = ~\b[1]  & ~new_n6579_;
  assign new_n6587_ = ~new_n6585_ & ~new_n6586_;
  assign new_n6588_ = \b[2]  & ~new_n6565_;
  assign new_n6589_ = ~new_n6560_ & new_n6588_;
  assign new_n6590_ = ~new_n6567_ & ~new_n6589_;
  assign new_n6591_ = ~new_n6587_ & new_n6590_;
  assign new_n6592_ = ~new_n6567_ & ~new_n6591_;
  assign new_n6593_ = \b[3]  & ~new_n6557_;
  assign new_n6594_ = ~new_n6551_ & new_n6593_;
  assign new_n6595_ = ~new_n6559_ & ~new_n6594_;
  assign new_n6596_ = ~new_n6592_ & new_n6595_;
  assign new_n6597_ = ~new_n6559_ & ~new_n6596_;
  assign new_n6598_ = \b[4]  & ~new_n6548_;
  assign new_n6599_ = ~new_n6542_ & new_n6598_;
  assign new_n6600_ = ~new_n6550_ & ~new_n6599_;
  assign new_n6601_ = ~new_n6597_ & new_n6600_;
  assign new_n6602_ = ~new_n6550_ & ~new_n6601_;
  assign new_n6603_ = \b[5]  & ~new_n6539_;
  assign new_n6604_ = ~new_n6533_ & new_n6603_;
  assign new_n6605_ = ~new_n6541_ & ~new_n6604_;
  assign new_n6606_ = ~new_n6602_ & new_n6605_;
  assign new_n6607_ = ~new_n6541_ & ~new_n6606_;
  assign new_n6608_ = \b[6]  & ~new_n6530_;
  assign new_n6609_ = ~new_n6524_ & new_n6608_;
  assign new_n6610_ = ~new_n6532_ & ~new_n6609_;
  assign new_n6611_ = ~new_n6607_ & new_n6610_;
  assign new_n6612_ = ~new_n6532_ & ~new_n6611_;
  assign new_n6613_ = \b[7]  & ~new_n6521_;
  assign new_n6614_ = ~new_n6515_ & new_n6613_;
  assign new_n6615_ = ~new_n6523_ & ~new_n6614_;
  assign new_n6616_ = ~new_n6612_ & new_n6615_;
  assign new_n6617_ = ~new_n6523_ & ~new_n6616_;
  assign new_n6618_ = \b[8]  & ~new_n6512_;
  assign new_n6619_ = ~new_n6506_ & new_n6618_;
  assign new_n6620_ = ~new_n6514_ & ~new_n6619_;
  assign new_n6621_ = ~new_n6617_ & new_n6620_;
  assign new_n6622_ = ~new_n6514_ & ~new_n6621_;
  assign new_n6623_ = \b[9]  & ~new_n6503_;
  assign new_n6624_ = ~new_n6497_ & new_n6623_;
  assign new_n6625_ = ~new_n6505_ & ~new_n6624_;
  assign new_n6626_ = ~new_n6622_ & new_n6625_;
  assign new_n6627_ = ~new_n6505_ & ~new_n6626_;
  assign new_n6628_ = \b[10]  & ~new_n6494_;
  assign new_n6629_ = ~new_n6488_ & new_n6628_;
  assign new_n6630_ = ~new_n6496_ & ~new_n6629_;
  assign new_n6631_ = ~new_n6627_ & new_n6630_;
  assign new_n6632_ = ~new_n6496_ & ~new_n6631_;
  assign new_n6633_ = \b[11]  & ~new_n6485_;
  assign new_n6634_ = ~new_n6479_ & new_n6633_;
  assign new_n6635_ = ~new_n6487_ & ~new_n6634_;
  assign new_n6636_ = ~new_n6632_ & new_n6635_;
  assign new_n6637_ = ~new_n6487_ & ~new_n6636_;
  assign new_n6638_ = \b[12]  & ~new_n6476_;
  assign new_n6639_ = ~new_n6470_ & new_n6638_;
  assign new_n6640_ = ~new_n6478_ & ~new_n6639_;
  assign new_n6641_ = ~new_n6637_ & new_n6640_;
  assign new_n6642_ = ~new_n6478_ & ~new_n6641_;
  assign new_n6643_ = \b[13]  & ~new_n6467_;
  assign new_n6644_ = ~new_n6461_ & new_n6643_;
  assign new_n6645_ = ~new_n6469_ & ~new_n6644_;
  assign new_n6646_ = ~new_n6642_ & new_n6645_;
  assign new_n6647_ = ~new_n6469_ & ~new_n6646_;
  assign new_n6648_ = \b[14]  & ~new_n6458_;
  assign new_n6649_ = ~new_n6452_ & new_n6648_;
  assign new_n6650_ = ~new_n6460_ & ~new_n6649_;
  assign new_n6651_ = ~new_n6647_ & new_n6650_;
  assign new_n6652_ = ~new_n6460_ & ~new_n6651_;
  assign new_n6653_ = \b[15]  & ~new_n6449_;
  assign new_n6654_ = ~new_n6443_ & new_n6653_;
  assign new_n6655_ = ~new_n6451_ & ~new_n6654_;
  assign new_n6656_ = ~new_n6652_ & new_n6655_;
  assign new_n6657_ = ~new_n6451_ & ~new_n6656_;
  assign new_n6658_ = \b[16]  & ~new_n6440_;
  assign new_n6659_ = ~new_n6434_ & new_n6658_;
  assign new_n6660_ = ~new_n6442_ & ~new_n6659_;
  assign new_n6661_ = ~new_n6657_ & new_n6660_;
  assign new_n6662_ = ~new_n6442_ & ~new_n6661_;
  assign new_n6663_ = \b[17]  & ~new_n6431_;
  assign new_n6664_ = ~new_n6425_ & new_n6663_;
  assign new_n6665_ = ~new_n6433_ & ~new_n6664_;
  assign new_n6666_ = ~new_n6662_ & new_n6665_;
  assign new_n6667_ = ~new_n6433_ & ~new_n6666_;
  assign new_n6668_ = \b[18]  & ~new_n6422_;
  assign new_n6669_ = ~new_n6416_ & new_n6668_;
  assign new_n6670_ = ~new_n6424_ & ~new_n6669_;
  assign new_n6671_ = ~new_n6667_ & new_n6670_;
  assign new_n6672_ = ~new_n6424_ & ~new_n6671_;
  assign new_n6673_ = \b[19]  & ~new_n6413_;
  assign new_n6674_ = ~new_n6407_ & new_n6673_;
  assign new_n6675_ = ~new_n6415_ & ~new_n6674_;
  assign new_n6676_ = ~new_n6672_ & new_n6675_;
  assign new_n6677_ = ~new_n6415_ & ~new_n6676_;
  assign new_n6678_ = \b[20]  & ~new_n6404_;
  assign new_n6679_ = ~new_n6398_ & new_n6678_;
  assign new_n6680_ = ~new_n6406_ & ~new_n6679_;
  assign new_n6681_ = ~new_n6677_ & new_n6680_;
  assign new_n6682_ = ~new_n6406_ & ~new_n6681_;
  assign new_n6683_ = \b[21]  & ~new_n6395_;
  assign new_n6684_ = ~new_n6389_ & new_n6683_;
  assign new_n6685_ = ~new_n6397_ & ~new_n6684_;
  assign new_n6686_ = ~new_n6682_ & new_n6685_;
  assign new_n6687_ = ~new_n6397_ & ~new_n6686_;
  assign new_n6688_ = \b[22]  & ~new_n6386_;
  assign new_n6689_ = ~new_n6380_ & new_n6688_;
  assign new_n6690_ = ~new_n6388_ & ~new_n6689_;
  assign new_n6691_ = ~new_n6687_ & new_n6690_;
  assign new_n6692_ = ~new_n6388_ & ~new_n6691_;
  assign new_n6693_ = \b[23]  & ~new_n6377_;
  assign new_n6694_ = ~new_n6371_ & new_n6693_;
  assign new_n6695_ = ~new_n6379_ & ~new_n6694_;
  assign new_n6696_ = ~new_n6692_ & new_n6695_;
  assign new_n6697_ = ~new_n6379_ & ~new_n6696_;
  assign new_n6698_ = \b[24]  & ~new_n6368_;
  assign new_n6699_ = ~new_n6362_ & new_n6698_;
  assign new_n6700_ = ~new_n6370_ & ~new_n6699_;
  assign new_n6701_ = ~new_n6697_ & new_n6700_;
  assign new_n6702_ = ~new_n6370_ & ~new_n6701_;
  assign new_n6703_ = \b[25]  & ~new_n6359_;
  assign new_n6704_ = ~new_n6353_ & new_n6703_;
  assign new_n6705_ = ~new_n6361_ & ~new_n6704_;
  assign new_n6706_ = ~new_n6702_ & new_n6705_;
  assign new_n6707_ = ~new_n6361_ & ~new_n6706_;
  assign new_n6708_ = \b[26]  & ~new_n6350_;
  assign new_n6709_ = ~new_n6344_ & new_n6708_;
  assign new_n6710_ = ~new_n6352_ & ~new_n6709_;
  assign new_n6711_ = ~new_n6707_ & new_n6710_;
  assign new_n6712_ = ~new_n6352_ & ~new_n6711_;
  assign new_n6713_ = \b[27]  & ~new_n6341_;
  assign new_n6714_ = ~new_n6335_ & new_n6713_;
  assign new_n6715_ = ~new_n6343_ & ~new_n6714_;
  assign new_n6716_ = ~new_n6712_ & new_n6715_;
  assign new_n6717_ = ~new_n6343_ & ~new_n6716_;
  assign new_n6718_ = \b[28]  & ~new_n6332_;
  assign new_n6719_ = ~new_n6326_ & new_n6718_;
  assign new_n6720_ = ~new_n6334_ & ~new_n6719_;
  assign new_n6721_ = ~new_n6717_ & new_n6720_;
  assign new_n6722_ = ~new_n6334_ & ~new_n6721_;
  assign new_n6723_ = ~new_n5942_ & ~\quotient[35] ;
  assign new_n6724_ = ~new_n5944_ & new_n6320_;
  assign new_n6725_ = ~new_n6316_ & new_n6724_;
  assign new_n6726_ = ~new_n6317_ & ~new_n6320_;
  assign new_n6727_ = ~new_n6725_ & ~new_n6726_;
  assign new_n6728_ = \quotient[35]  & ~new_n6727_;
  assign new_n6729_ = ~new_n6723_ & ~new_n6728_;
  assign new_n6730_ = ~\b[29]  & ~new_n6729_;
  assign new_n6731_ = \b[29]  & ~new_n6723_;
  assign new_n6732_ = ~new_n6728_ & new_n6731_;
  assign new_n6733_ = new_n313_ & new_n315_;
  assign new_n6734_ = new_n303_ & new_n6733_;
  assign new_n6735_ = new_n288_ & new_n6734_;
  assign new_n6736_ = ~new_n6732_ & new_n6735_;
  assign new_n6737_ = ~new_n6730_ & new_n6736_;
  assign new_n6738_ = ~new_n6722_ & new_n6737_;
  assign new_n6739_ = new_n6324_ & ~new_n6729_;
  assign \quotient[34]  = new_n6738_ | new_n6739_;
  assign new_n6741_ = ~new_n6343_ & new_n6720_;
  assign new_n6742_ = ~new_n6716_ & new_n6741_;
  assign new_n6743_ = ~new_n6717_ & ~new_n6720_;
  assign new_n6744_ = ~new_n6742_ & ~new_n6743_;
  assign new_n6745_ = \quotient[34]  & ~new_n6744_;
  assign new_n6746_ = ~new_n6333_ & ~new_n6739_;
  assign new_n6747_ = ~new_n6738_ & new_n6746_;
  assign new_n6748_ = ~new_n6745_ & ~new_n6747_;
  assign new_n6749_ = ~new_n6334_ & ~new_n6732_;
  assign new_n6750_ = ~new_n6730_ & new_n6749_;
  assign new_n6751_ = ~new_n6721_ & new_n6750_;
  assign new_n6752_ = ~new_n6730_ & ~new_n6732_;
  assign new_n6753_ = ~new_n6722_ & ~new_n6752_;
  assign new_n6754_ = ~new_n6751_ & ~new_n6753_;
  assign new_n6755_ = \quotient[34]  & ~new_n6754_;
  assign new_n6756_ = ~new_n6729_ & ~new_n6739_;
  assign new_n6757_ = ~new_n6738_ & new_n6756_;
  assign new_n6758_ = ~new_n6755_ & ~new_n6757_;
  assign new_n6759_ = ~\b[30]  & ~new_n6758_;
  assign new_n6760_ = ~\b[29]  & ~new_n6748_;
  assign new_n6761_ = ~new_n6352_ & new_n6715_;
  assign new_n6762_ = ~new_n6711_ & new_n6761_;
  assign new_n6763_ = ~new_n6712_ & ~new_n6715_;
  assign new_n6764_ = ~new_n6762_ & ~new_n6763_;
  assign new_n6765_ = \quotient[34]  & ~new_n6764_;
  assign new_n6766_ = ~new_n6342_ & ~new_n6739_;
  assign new_n6767_ = ~new_n6738_ & new_n6766_;
  assign new_n6768_ = ~new_n6765_ & ~new_n6767_;
  assign new_n6769_ = ~\b[28]  & ~new_n6768_;
  assign new_n6770_ = ~new_n6361_ & new_n6710_;
  assign new_n6771_ = ~new_n6706_ & new_n6770_;
  assign new_n6772_ = ~new_n6707_ & ~new_n6710_;
  assign new_n6773_ = ~new_n6771_ & ~new_n6772_;
  assign new_n6774_ = \quotient[34]  & ~new_n6773_;
  assign new_n6775_ = ~new_n6351_ & ~new_n6739_;
  assign new_n6776_ = ~new_n6738_ & new_n6775_;
  assign new_n6777_ = ~new_n6774_ & ~new_n6776_;
  assign new_n6778_ = ~\b[27]  & ~new_n6777_;
  assign new_n6779_ = ~new_n6370_ & new_n6705_;
  assign new_n6780_ = ~new_n6701_ & new_n6779_;
  assign new_n6781_ = ~new_n6702_ & ~new_n6705_;
  assign new_n6782_ = ~new_n6780_ & ~new_n6781_;
  assign new_n6783_ = \quotient[34]  & ~new_n6782_;
  assign new_n6784_ = ~new_n6360_ & ~new_n6739_;
  assign new_n6785_ = ~new_n6738_ & new_n6784_;
  assign new_n6786_ = ~new_n6783_ & ~new_n6785_;
  assign new_n6787_ = ~\b[26]  & ~new_n6786_;
  assign new_n6788_ = ~new_n6379_ & new_n6700_;
  assign new_n6789_ = ~new_n6696_ & new_n6788_;
  assign new_n6790_ = ~new_n6697_ & ~new_n6700_;
  assign new_n6791_ = ~new_n6789_ & ~new_n6790_;
  assign new_n6792_ = \quotient[34]  & ~new_n6791_;
  assign new_n6793_ = ~new_n6369_ & ~new_n6739_;
  assign new_n6794_ = ~new_n6738_ & new_n6793_;
  assign new_n6795_ = ~new_n6792_ & ~new_n6794_;
  assign new_n6796_ = ~\b[25]  & ~new_n6795_;
  assign new_n6797_ = ~new_n6388_ & new_n6695_;
  assign new_n6798_ = ~new_n6691_ & new_n6797_;
  assign new_n6799_ = ~new_n6692_ & ~new_n6695_;
  assign new_n6800_ = ~new_n6798_ & ~new_n6799_;
  assign new_n6801_ = \quotient[34]  & ~new_n6800_;
  assign new_n6802_ = ~new_n6378_ & ~new_n6739_;
  assign new_n6803_ = ~new_n6738_ & new_n6802_;
  assign new_n6804_ = ~new_n6801_ & ~new_n6803_;
  assign new_n6805_ = ~\b[24]  & ~new_n6804_;
  assign new_n6806_ = ~new_n6397_ & new_n6690_;
  assign new_n6807_ = ~new_n6686_ & new_n6806_;
  assign new_n6808_ = ~new_n6687_ & ~new_n6690_;
  assign new_n6809_ = ~new_n6807_ & ~new_n6808_;
  assign new_n6810_ = \quotient[34]  & ~new_n6809_;
  assign new_n6811_ = ~new_n6387_ & ~new_n6739_;
  assign new_n6812_ = ~new_n6738_ & new_n6811_;
  assign new_n6813_ = ~new_n6810_ & ~new_n6812_;
  assign new_n6814_ = ~\b[23]  & ~new_n6813_;
  assign new_n6815_ = ~new_n6406_ & new_n6685_;
  assign new_n6816_ = ~new_n6681_ & new_n6815_;
  assign new_n6817_ = ~new_n6682_ & ~new_n6685_;
  assign new_n6818_ = ~new_n6816_ & ~new_n6817_;
  assign new_n6819_ = \quotient[34]  & ~new_n6818_;
  assign new_n6820_ = ~new_n6396_ & ~new_n6739_;
  assign new_n6821_ = ~new_n6738_ & new_n6820_;
  assign new_n6822_ = ~new_n6819_ & ~new_n6821_;
  assign new_n6823_ = ~\b[22]  & ~new_n6822_;
  assign new_n6824_ = ~new_n6415_ & new_n6680_;
  assign new_n6825_ = ~new_n6676_ & new_n6824_;
  assign new_n6826_ = ~new_n6677_ & ~new_n6680_;
  assign new_n6827_ = ~new_n6825_ & ~new_n6826_;
  assign new_n6828_ = \quotient[34]  & ~new_n6827_;
  assign new_n6829_ = ~new_n6405_ & ~new_n6739_;
  assign new_n6830_ = ~new_n6738_ & new_n6829_;
  assign new_n6831_ = ~new_n6828_ & ~new_n6830_;
  assign new_n6832_ = ~\b[21]  & ~new_n6831_;
  assign new_n6833_ = ~new_n6424_ & new_n6675_;
  assign new_n6834_ = ~new_n6671_ & new_n6833_;
  assign new_n6835_ = ~new_n6672_ & ~new_n6675_;
  assign new_n6836_ = ~new_n6834_ & ~new_n6835_;
  assign new_n6837_ = \quotient[34]  & ~new_n6836_;
  assign new_n6838_ = ~new_n6414_ & ~new_n6739_;
  assign new_n6839_ = ~new_n6738_ & new_n6838_;
  assign new_n6840_ = ~new_n6837_ & ~new_n6839_;
  assign new_n6841_ = ~\b[20]  & ~new_n6840_;
  assign new_n6842_ = ~new_n6433_ & new_n6670_;
  assign new_n6843_ = ~new_n6666_ & new_n6842_;
  assign new_n6844_ = ~new_n6667_ & ~new_n6670_;
  assign new_n6845_ = ~new_n6843_ & ~new_n6844_;
  assign new_n6846_ = \quotient[34]  & ~new_n6845_;
  assign new_n6847_ = ~new_n6423_ & ~new_n6739_;
  assign new_n6848_ = ~new_n6738_ & new_n6847_;
  assign new_n6849_ = ~new_n6846_ & ~new_n6848_;
  assign new_n6850_ = ~\b[19]  & ~new_n6849_;
  assign new_n6851_ = ~new_n6442_ & new_n6665_;
  assign new_n6852_ = ~new_n6661_ & new_n6851_;
  assign new_n6853_ = ~new_n6662_ & ~new_n6665_;
  assign new_n6854_ = ~new_n6852_ & ~new_n6853_;
  assign new_n6855_ = \quotient[34]  & ~new_n6854_;
  assign new_n6856_ = ~new_n6432_ & ~new_n6739_;
  assign new_n6857_ = ~new_n6738_ & new_n6856_;
  assign new_n6858_ = ~new_n6855_ & ~new_n6857_;
  assign new_n6859_ = ~\b[18]  & ~new_n6858_;
  assign new_n6860_ = ~new_n6451_ & new_n6660_;
  assign new_n6861_ = ~new_n6656_ & new_n6860_;
  assign new_n6862_ = ~new_n6657_ & ~new_n6660_;
  assign new_n6863_ = ~new_n6861_ & ~new_n6862_;
  assign new_n6864_ = \quotient[34]  & ~new_n6863_;
  assign new_n6865_ = ~new_n6441_ & ~new_n6739_;
  assign new_n6866_ = ~new_n6738_ & new_n6865_;
  assign new_n6867_ = ~new_n6864_ & ~new_n6866_;
  assign new_n6868_ = ~\b[17]  & ~new_n6867_;
  assign new_n6869_ = ~new_n6460_ & new_n6655_;
  assign new_n6870_ = ~new_n6651_ & new_n6869_;
  assign new_n6871_ = ~new_n6652_ & ~new_n6655_;
  assign new_n6872_ = ~new_n6870_ & ~new_n6871_;
  assign new_n6873_ = \quotient[34]  & ~new_n6872_;
  assign new_n6874_ = ~new_n6450_ & ~new_n6739_;
  assign new_n6875_ = ~new_n6738_ & new_n6874_;
  assign new_n6876_ = ~new_n6873_ & ~new_n6875_;
  assign new_n6877_ = ~\b[16]  & ~new_n6876_;
  assign new_n6878_ = ~new_n6469_ & new_n6650_;
  assign new_n6879_ = ~new_n6646_ & new_n6878_;
  assign new_n6880_ = ~new_n6647_ & ~new_n6650_;
  assign new_n6881_ = ~new_n6879_ & ~new_n6880_;
  assign new_n6882_ = \quotient[34]  & ~new_n6881_;
  assign new_n6883_ = ~new_n6459_ & ~new_n6739_;
  assign new_n6884_ = ~new_n6738_ & new_n6883_;
  assign new_n6885_ = ~new_n6882_ & ~new_n6884_;
  assign new_n6886_ = ~\b[15]  & ~new_n6885_;
  assign new_n6887_ = ~new_n6478_ & new_n6645_;
  assign new_n6888_ = ~new_n6641_ & new_n6887_;
  assign new_n6889_ = ~new_n6642_ & ~new_n6645_;
  assign new_n6890_ = ~new_n6888_ & ~new_n6889_;
  assign new_n6891_ = \quotient[34]  & ~new_n6890_;
  assign new_n6892_ = ~new_n6468_ & ~new_n6739_;
  assign new_n6893_ = ~new_n6738_ & new_n6892_;
  assign new_n6894_ = ~new_n6891_ & ~new_n6893_;
  assign new_n6895_ = ~\b[14]  & ~new_n6894_;
  assign new_n6896_ = ~new_n6487_ & new_n6640_;
  assign new_n6897_ = ~new_n6636_ & new_n6896_;
  assign new_n6898_ = ~new_n6637_ & ~new_n6640_;
  assign new_n6899_ = ~new_n6897_ & ~new_n6898_;
  assign new_n6900_ = \quotient[34]  & ~new_n6899_;
  assign new_n6901_ = ~new_n6477_ & ~new_n6739_;
  assign new_n6902_ = ~new_n6738_ & new_n6901_;
  assign new_n6903_ = ~new_n6900_ & ~new_n6902_;
  assign new_n6904_ = ~\b[13]  & ~new_n6903_;
  assign new_n6905_ = ~new_n6496_ & new_n6635_;
  assign new_n6906_ = ~new_n6631_ & new_n6905_;
  assign new_n6907_ = ~new_n6632_ & ~new_n6635_;
  assign new_n6908_ = ~new_n6906_ & ~new_n6907_;
  assign new_n6909_ = \quotient[34]  & ~new_n6908_;
  assign new_n6910_ = ~new_n6486_ & ~new_n6739_;
  assign new_n6911_ = ~new_n6738_ & new_n6910_;
  assign new_n6912_ = ~new_n6909_ & ~new_n6911_;
  assign new_n6913_ = ~\b[12]  & ~new_n6912_;
  assign new_n6914_ = ~new_n6505_ & new_n6630_;
  assign new_n6915_ = ~new_n6626_ & new_n6914_;
  assign new_n6916_ = ~new_n6627_ & ~new_n6630_;
  assign new_n6917_ = ~new_n6915_ & ~new_n6916_;
  assign new_n6918_ = \quotient[34]  & ~new_n6917_;
  assign new_n6919_ = ~new_n6495_ & ~new_n6739_;
  assign new_n6920_ = ~new_n6738_ & new_n6919_;
  assign new_n6921_ = ~new_n6918_ & ~new_n6920_;
  assign new_n6922_ = ~\b[11]  & ~new_n6921_;
  assign new_n6923_ = ~new_n6514_ & new_n6625_;
  assign new_n6924_ = ~new_n6621_ & new_n6923_;
  assign new_n6925_ = ~new_n6622_ & ~new_n6625_;
  assign new_n6926_ = ~new_n6924_ & ~new_n6925_;
  assign new_n6927_ = \quotient[34]  & ~new_n6926_;
  assign new_n6928_ = ~new_n6504_ & ~new_n6739_;
  assign new_n6929_ = ~new_n6738_ & new_n6928_;
  assign new_n6930_ = ~new_n6927_ & ~new_n6929_;
  assign new_n6931_ = ~\b[10]  & ~new_n6930_;
  assign new_n6932_ = ~new_n6523_ & new_n6620_;
  assign new_n6933_ = ~new_n6616_ & new_n6932_;
  assign new_n6934_ = ~new_n6617_ & ~new_n6620_;
  assign new_n6935_ = ~new_n6933_ & ~new_n6934_;
  assign new_n6936_ = \quotient[34]  & ~new_n6935_;
  assign new_n6937_ = ~new_n6513_ & ~new_n6739_;
  assign new_n6938_ = ~new_n6738_ & new_n6937_;
  assign new_n6939_ = ~new_n6936_ & ~new_n6938_;
  assign new_n6940_ = ~\b[9]  & ~new_n6939_;
  assign new_n6941_ = ~new_n6532_ & new_n6615_;
  assign new_n6942_ = ~new_n6611_ & new_n6941_;
  assign new_n6943_ = ~new_n6612_ & ~new_n6615_;
  assign new_n6944_ = ~new_n6942_ & ~new_n6943_;
  assign new_n6945_ = \quotient[34]  & ~new_n6944_;
  assign new_n6946_ = ~new_n6522_ & ~new_n6739_;
  assign new_n6947_ = ~new_n6738_ & new_n6946_;
  assign new_n6948_ = ~new_n6945_ & ~new_n6947_;
  assign new_n6949_ = ~\b[8]  & ~new_n6948_;
  assign new_n6950_ = ~new_n6541_ & new_n6610_;
  assign new_n6951_ = ~new_n6606_ & new_n6950_;
  assign new_n6952_ = ~new_n6607_ & ~new_n6610_;
  assign new_n6953_ = ~new_n6951_ & ~new_n6952_;
  assign new_n6954_ = \quotient[34]  & ~new_n6953_;
  assign new_n6955_ = ~new_n6531_ & ~new_n6739_;
  assign new_n6956_ = ~new_n6738_ & new_n6955_;
  assign new_n6957_ = ~new_n6954_ & ~new_n6956_;
  assign new_n6958_ = ~\b[7]  & ~new_n6957_;
  assign new_n6959_ = ~new_n6550_ & new_n6605_;
  assign new_n6960_ = ~new_n6601_ & new_n6959_;
  assign new_n6961_ = ~new_n6602_ & ~new_n6605_;
  assign new_n6962_ = ~new_n6960_ & ~new_n6961_;
  assign new_n6963_ = \quotient[34]  & ~new_n6962_;
  assign new_n6964_ = ~new_n6540_ & ~new_n6739_;
  assign new_n6965_ = ~new_n6738_ & new_n6964_;
  assign new_n6966_ = ~new_n6963_ & ~new_n6965_;
  assign new_n6967_ = ~\b[6]  & ~new_n6966_;
  assign new_n6968_ = ~new_n6559_ & new_n6600_;
  assign new_n6969_ = ~new_n6596_ & new_n6968_;
  assign new_n6970_ = ~new_n6597_ & ~new_n6600_;
  assign new_n6971_ = ~new_n6969_ & ~new_n6970_;
  assign new_n6972_ = \quotient[34]  & ~new_n6971_;
  assign new_n6973_ = ~new_n6549_ & ~new_n6739_;
  assign new_n6974_ = ~new_n6738_ & new_n6973_;
  assign new_n6975_ = ~new_n6972_ & ~new_n6974_;
  assign new_n6976_ = ~\b[5]  & ~new_n6975_;
  assign new_n6977_ = ~new_n6567_ & new_n6595_;
  assign new_n6978_ = ~new_n6591_ & new_n6977_;
  assign new_n6979_ = ~new_n6592_ & ~new_n6595_;
  assign new_n6980_ = ~new_n6978_ & ~new_n6979_;
  assign new_n6981_ = \quotient[34]  & ~new_n6980_;
  assign new_n6982_ = ~new_n6558_ & ~new_n6739_;
  assign new_n6983_ = ~new_n6738_ & new_n6982_;
  assign new_n6984_ = ~new_n6981_ & ~new_n6983_;
  assign new_n6985_ = ~\b[4]  & ~new_n6984_;
  assign new_n6986_ = ~new_n6586_ & new_n6590_;
  assign new_n6987_ = ~new_n6585_ & new_n6986_;
  assign new_n6988_ = ~new_n6587_ & ~new_n6590_;
  assign new_n6989_ = ~new_n6987_ & ~new_n6988_;
  assign new_n6990_ = \quotient[34]  & ~new_n6989_;
  assign new_n6991_ = ~new_n6566_ & ~new_n6739_;
  assign new_n6992_ = ~new_n6738_ & new_n6991_;
  assign new_n6993_ = ~new_n6990_ & ~new_n6992_;
  assign new_n6994_ = ~\b[3]  & ~new_n6993_;
  assign new_n6995_ = ~new_n6582_ & new_n6584_;
  assign new_n6996_ = ~new_n6580_ & new_n6995_;
  assign new_n6997_ = ~new_n6585_ & ~new_n6996_;
  assign new_n6998_ = \quotient[34]  & new_n6997_;
  assign new_n6999_ = ~new_n6579_ & ~new_n6739_;
  assign new_n7000_ = ~new_n6738_ & new_n6999_;
  assign new_n7001_ = ~new_n6998_ & ~new_n7000_;
  assign new_n7002_ = ~\b[2]  & ~new_n7001_;
  assign new_n7003_ = \b[0]  & \quotient[34] ;
  assign new_n7004_ = \a[34]  & ~new_n7003_;
  assign new_n7005_ = new_n6584_ & \quotient[34] ;
  assign new_n7006_ = ~new_n7004_ & ~new_n7005_;
  assign new_n7007_ = \b[1]  & ~new_n7006_;
  assign new_n7008_ = ~\b[1]  & ~new_n7005_;
  assign new_n7009_ = ~new_n7004_ & new_n7008_;
  assign new_n7010_ = ~new_n7007_ & ~new_n7009_;
  assign new_n7011_ = ~\a[33]  & \b[0] ;
  assign new_n7012_ = ~new_n7010_ & ~new_n7011_;
  assign new_n7013_ = ~\b[1]  & ~new_n7006_;
  assign new_n7014_ = ~new_n7012_ & ~new_n7013_;
  assign new_n7015_ = \b[2]  & ~new_n7000_;
  assign new_n7016_ = ~new_n6998_ & new_n7015_;
  assign new_n7017_ = ~new_n7002_ & ~new_n7016_;
  assign new_n7018_ = ~new_n7014_ & new_n7017_;
  assign new_n7019_ = ~new_n7002_ & ~new_n7018_;
  assign new_n7020_ = \b[3]  & ~new_n6992_;
  assign new_n7021_ = ~new_n6990_ & new_n7020_;
  assign new_n7022_ = ~new_n6994_ & ~new_n7021_;
  assign new_n7023_ = ~new_n7019_ & new_n7022_;
  assign new_n7024_ = ~new_n6994_ & ~new_n7023_;
  assign new_n7025_ = \b[4]  & ~new_n6983_;
  assign new_n7026_ = ~new_n6981_ & new_n7025_;
  assign new_n7027_ = ~new_n6985_ & ~new_n7026_;
  assign new_n7028_ = ~new_n7024_ & new_n7027_;
  assign new_n7029_ = ~new_n6985_ & ~new_n7028_;
  assign new_n7030_ = \b[5]  & ~new_n6974_;
  assign new_n7031_ = ~new_n6972_ & new_n7030_;
  assign new_n7032_ = ~new_n6976_ & ~new_n7031_;
  assign new_n7033_ = ~new_n7029_ & new_n7032_;
  assign new_n7034_ = ~new_n6976_ & ~new_n7033_;
  assign new_n7035_ = \b[6]  & ~new_n6965_;
  assign new_n7036_ = ~new_n6963_ & new_n7035_;
  assign new_n7037_ = ~new_n6967_ & ~new_n7036_;
  assign new_n7038_ = ~new_n7034_ & new_n7037_;
  assign new_n7039_ = ~new_n6967_ & ~new_n7038_;
  assign new_n7040_ = \b[7]  & ~new_n6956_;
  assign new_n7041_ = ~new_n6954_ & new_n7040_;
  assign new_n7042_ = ~new_n6958_ & ~new_n7041_;
  assign new_n7043_ = ~new_n7039_ & new_n7042_;
  assign new_n7044_ = ~new_n6958_ & ~new_n7043_;
  assign new_n7045_ = \b[8]  & ~new_n6947_;
  assign new_n7046_ = ~new_n6945_ & new_n7045_;
  assign new_n7047_ = ~new_n6949_ & ~new_n7046_;
  assign new_n7048_ = ~new_n7044_ & new_n7047_;
  assign new_n7049_ = ~new_n6949_ & ~new_n7048_;
  assign new_n7050_ = \b[9]  & ~new_n6938_;
  assign new_n7051_ = ~new_n6936_ & new_n7050_;
  assign new_n7052_ = ~new_n6940_ & ~new_n7051_;
  assign new_n7053_ = ~new_n7049_ & new_n7052_;
  assign new_n7054_ = ~new_n6940_ & ~new_n7053_;
  assign new_n7055_ = \b[10]  & ~new_n6929_;
  assign new_n7056_ = ~new_n6927_ & new_n7055_;
  assign new_n7057_ = ~new_n6931_ & ~new_n7056_;
  assign new_n7058_ = ~new_n7054_ & new_n7057_;
  assign new_n7059_ = ~new_n6931_ & ~new_n7058_;
  assign new_n7060_ = \b[11]  & ~new_n6920_;
  assign new_n7061_ = ~new_n6918_ & new_n7060_;
  assign new_n7062_ = ~new_n6922_ & ~new_n7061_;
  assign new_n7063_ = ~new_n7059_ & new_n7062_;
  assign new_n7064_ = ~new_n6922_ & ~new_n7063_;
  assign new_n7065_ = \b[12]  & ~new_n6911_;
  assign new_n7066_ = ~new_n6909_ & new_n7065_;
  assign new_n7067_ = ~new_n6913_ & ~new_n7066_;
  assign new_n7068_ = ~new_n7064_ & new_n7067_;
  assign new_n7069_ = ~new_n6913_ & ~new_n7068_;
  assign new_n7070_ = \b[13]  & ~new_n6902_;
  assign new_n7071_ = ~new_n6900_ & new_n7070_;
  assign new_n7072_ = ~new_n6904_ & ~new_n7071_;
  assign new_n7073_ = ~new_n7069_ & new_n7072_;
  assign new_n7074_ = ~new_n6904_ & ~new_n7073_;
  assign new_n7075_ = \b[14]  & ~new_n6893_;
  assign new_n7076_ = ~new_n6891_ & new_n7075_;
  assign new_n7077_ = ~new_n6895_ & ~new_n7076_;
  assign new_n7078_ = ~new_n7074_ & new_n7077_;
  assign new_n7079_ = ~new_n6895_ & ~new_n7078_;
  assign new_n7080_ = \b[15]  & ~new_n6884_;
  assign new_n7081_ = ~new_n6882_ & new_n7080_;
  assign new_n7082_ = ~new_n6886_ & ~new_n7081_;
  assign new_n7083_ = ~new_n7079_ & new_n7082_;
  assign new_n7084_ = ~new_n6886_ & ~new_n7083_;
  assign new_n7085_ = \b[16]  & ~new_n6875_;
  assign new_n7086_ = ~new_n6873_ & new_n7085_;
  assign new_n7087_ = ~new_n6877_ & ~new_n7086_;
  assign new_n7088_ = ~new_n7084_ & new_n7087_;
  assign new_n7089_ = ~new_n6877_ & ~new_n7088_;
  assign new_n7090_ = \b[17]  & ~new_n6866_;
  assign new_n7091_ = ~new_n6864_ & new_n7090_;
  assign new_n7092_ = ~new_n6868_ & ~new_n7091_;
  assign new_n7093_ = ~new_n7089_ & new_n7092_;
  assign new_n7094_ = ~new_n6868_ & ~new_n7093_;
  assign new_n7095_ = \b[18]  & ~new_n6857_;
  assign new_n7096_ = ~new_n6855_ & new_n7095_;
  assign new_n7097_ = ~new_n6859_ & ~new_n7096_;
  assign new_n7098_ = ~new_n7094_ & new_n7097_;
  assign new_n7099_ = ~new_n6859_ & ~new_n7098_;
  assign new_n7100_ = \b[19]  & ~new_n6848_;
  assign new_n7101_ = ~new_n6846_ & new_n7100_;
  assign new_n7102_ = ~new_n6850_ & ~new_n7101_;
  assign new_n7103_ = ~new_n7099_ & new_n7102_;
  assign new_n7104_ = ~new_n6850_ & ~new_n7103_;
  assign new_n7105_ = \b[20]  & ~new_n6839_;
  assign new_n7106_ = ~new_n6837_ & new_n7105_;
  assign new_n7107_ = ~new_n6841_ & ~new_n7106_;
  assign new_n7108_ = ~new_n7104_ & new_n7107_;
  assign new_n7109_ = ~new_n6841_ & ~new_n7108_;
  assign new_n7110_ = \b[21]  & ~new_n6830_;
  assign new_n7111_ = ~new_n6828_ & new_n7110_;
  assign new_n7112_ = ~new_n6832_ & ~new_n7111_;
  assign new_n7113_ = ~new_n7109_ & new_n7112_;
  assign new_n7114_ = ~new_n6832_ & ~new_n7113_;
  assign new_n7115_ = \b[22]  & ~new_n6821_;
  assign new_n7116_ = ~new_n6819_ & new_n7115_;
  assign new_n7117_ = ~new_n6823_ & ~new_n7116_;
  assign new_n7118_ = ~new_n7114_ & new_n7117_;
  assign new_n7119_ = ~new_n6823_ & ~new_n7118_;
  assign new_n7120_ = \b[23]  & ~new_n6812_;
  assign new_n7121_ = ~new_n6810_ & new_n7120_;
  assign new_n7122_ = ~new_n6814_ & ~new_n7121_;
  assign new_n7123_ = ~new_n7119_ & new_n7122_;
  assign new_n7124_ = ~new_n6814_ & ~new_n7123_;
  assign new_n7125_ = \b[24]  & ~new_n6803_;
  assign new_n7126_ = ~new_n6801_ & new_n7125_;
  assign new_n7127_ = ~new_n6805_ & ~new_n7126_;
  assign new_n7128_ = ~new_n7124_ & new_n7127_;
  assign new_n7129_ = ~new_n6805_ & ~new_n7128_;
  assign new_n7130_ = \b[25]  & ~new_n6794_;
  assign new_n7131_ = ~new_n6792_ & new_n7130_;
  assign new_n7132_ = ~new_n6796_ & ~new_n7131_;
  assign new_n7133_ = ~new_n7129_ & new_n7132_;
  assign new_n7134_ = ~new_n6796_ & ~new_n7133_;
  assign new_n7135_ = \b[26]  & ~new_n6785_;
  assign new_n7136_ = ~new_n6783_ & new_n7135_;
  assign new_n7137_ = ~new_n6787_ & ~new_n7136_;
  assign new_n7138_ = ~new_n7134_ & new_n7137_;
  assign new_n7139_ = ~new_n6787_ & ~new_n7138_;
  assign new_n7140_ = \b[27]  & ~new_n6776_;
  assign new_n7141_ = ~new_n6774_ & new_n7140_;
  assign new_n7142_ = ~new_n6778_ & ~new_n7141_;
  assign new_n7143_ = ~new_n7139_ & new_n7142_;
  assign new_n7144_ = ~new_n6778_ & ~new_n7143_;
  assign new_n7145_ = \b[28]  & ~new_n6767_;
  assign new_n7146_ = ~new_n6765_ & new_n7145_;
  assign new_n7147_ = ~new_n6769_ & ~new_n7146_;
  assign new_n7148_ = ~new_n7144_ & new_n7147_;
  assign new_n7149_ = ~new_n6769_ & ~new_n7148_;
  assign new_n7150_ = \b[29]  & ~new_n6747_;
  assign new_n7151_ = ~new_n6745_ & new_n7150_;
  assign new_n7152_ = ~new_n6760_ & ~new_n7151_;
  assign new_n7153_ = ~new_n7149_ & new_n7152_;
  assign new_n7154_ = ~new_n6760_ & ~new_n7153_;
  assign new_n7155_ = \b[30]  & ~new_n6757_;
  assign new_n7156_ = ~new_n6755_ & new_n7155_;
  assign new_n7157_ = ~new_n6759_ & ~new_n7156_;
  assign new_n7158_ = ~new_n7154_ & new_n7157_;
  assign new_n7159_ = ~new_n6759_ & ~new_n7158_;
  assign new_n7160_ = new_n372_ & new_n414_;
  assign new_n7161_ = new_n598_ & new_n7160_;
  assign new_n7162_ = new_n595_ & new_n7161_;
  assign \quotient[33]  = ~new_n7159_ & new_n7162_;
  assign new_n7164_ = ~new_n6748_ & ~\quotient[33] ;
  assign new_n7165_ = ~new_n6769_ & new_n7152_;
  assign new_n7166_ = ~new_n7148_ & new_n7165_;
  assign new_n7167_ = ~new_n7149_ & ~new_n7152_;
  assign new_n7168_ = ~new_n7166_ & ~new_n7167_;
  assign new_n7169_ = new_n7162_ & ~new_n7168_;
  assign new_n7170_ = ~new_n7159_ & new_n7169_;
  assign new_n7171_ = ~new_n7164_ & ~new_n7170_;
  assign new_n7172_ = ~new_n6758_ & ~\quotient[33] ;
  assign new_n7173_ = ~new_n6760_ & new_n7157_;
  assign new_n7174_ = ~new_n7153_ & new_n7173_;
  assign new_n7175_ = ~new_n7154_ & ~new_n7157_;
  assign new_n7176_ = ~new_n7174_ & ~new_n7175_;
  assign new_n7177_ = \quotient[33]  & ~new_n7176_;
  assign new_n7178_ = ~new_n7172_ & ~new_n7177_;
  assign new_n7179_ = ~\b[31]  & ~new_n7178_;
  assign new_n7180_ = ~\b[30]  & ~new_n7171_;
  assign new_n7181_ = ~new_n6768_ & ~\quotient[33] ;
  assign new_n7182_ = ~new_n6778_ & new_n7147_;
  assign new_n7183_ = ~new_n7143_ & new_n7182_;
  assign new_n7184_ = ~new_n7144_ & ~new_n7147_;
  assign new_n7185_ = ~new_n7183_ & ~new_n7184_;
  assign new_n7186_ = new_n7162_ & ~new_n7185_;
  assign new_n7187_ = ~new_n7159_ & new_n7186_;
  assign new_n7188_ = ~new_n7181_ & ~new_n7187_;
  assign new_n7189_ = ~\b[29]  & ~new_n7188_;
  assign new_n7190_ = ~new_n6777_ & ~\quotient[33] ;
  assign new_n7191_ = ~new_n6787_ & new_n7142_;
  assign new_n7192_ = ~new_n7138_ & new_n7191_;
  assign new_n7193_ = ~new_n7139_ & ~new_n7142_;
  assign new_n7194_ = ~new_n7192_ & ~new_n7193_;
  assign new_n7195_ = new_n7162_ & ~new_n7194_;
  assign new_n7196_ = ~new_n7159_ & new_n7195_;
  assign new_n7197_ = ~new_n7190_ & ~new_n7196_;
  assign new_n7198_ = ~\b[28]  & ~new_n7197_;
  assign new_n7199_ = ~new_n6786_ & ~\quotient[33] ;
  assign new_n7200_ = ~new_n6796_ & new_n7137_;
  assign new_n7201_ = ~new_n7133_ & new_n7200_;
  assign new_n7202_ = ~new_n7134_ & ~new_n7137_;
  assign new_n7203_ = ~new_n7201_ & ~new_n7202_;
  assign new_n7204_ = new_n7162_ & ~new_n7203_;
  assign new_n7205_ = ~new_n7159_ & new_n7204_;
  assign new_n7206_ = ~new_n7199_ & ~new_n7205_;
  assign new_n7207_ = ~\b[27]  & ~new_n7206_;
  assign new_n7208_ = ~new_n6795_ & ~\quotient[33] ;
  assign new_n7209_ = ~new_n6805_ & new_n7132_;
  assign new_n7210_ = ~new_n7128_ & new_n7209_;
  assign new_n7211_ = ~new_n7129_ & ~new_n7132_;
  assign new_n7212_ = ~new_n7210_ & ~new_n7211_;
  assign new_n7213_ = new_n7162_ & ~new_n7212_;
  assign new_n7214_ = ~new_n7159_ & new_n7213_;
  assign new_n7215_ = ~new_n7208_ & ~new_n7214_;
  assign new_n7216_ = ~\b[26]  & ~new_n7215_;
  assign new_n7217_ = ~new_n6804_ & ~\quotient[33] ;
  assign new_n7218_ = ~new_n6814_ & new_n7127_;
  assign new_n7219_ = ~new_n7123_ & new_n7218_;
  assign new_n7220_ = ~new_n7124_ & ~new_n7127_;
  assign new_n7221_ = ~new_n7219_ & ~new_n7220_;
  assign new_n7222_ = new_n7162_ & ~new_n7221_;
  assign new_n7223_ = ~new_n7159_ & new_n7222_;
  assign new_n7224_ = ~new_n7217_ & ~new_n7223_;
  assign new_n7225_ = ~\b[25]  & ~new_n7224_;
  assign new_n7226_ = ~new_n6813_ & ~\quotient[33] ;
  assign new_n7227_ = ~new_n6823_ & new_n7122_;
  assign new_n7228_ = ~new_n7118_ & new_n7227_;
  assign new_n7229_ = ~new_n7119_ & ~new_n7122_;
  assign new_n7230_ = ~new_n7228_ & ~new_n7229_;
  assign new_n7231_ = new_n7162_ & ~new_n7230_;
  assign new_n7232_ = ~new_n7159_ & new_n7231_;
  assign new_n7233_ = ~new_n7226_ & ~new_n7232_;
  assign new_n7234_ = ~\b[24]  & ~new_n7233_;
  assign new_n7235_ = ~new_n6822_ & ~\quotient[33] ;
  assign new_n7236_ = ~new_n6832_ & new_n7117_;
  assign new_n7237_ = ~new_n7113_ & new_n7236_;
  assign new_n7238_ = ~new_n7114_ & ~new_n7117_;
  assign new_n7239_ = ~new_n7237_ & ~new_n7238_;
  assign new_n7240_ = new_n7162_ & ~new_n7239_;
  assign new_n7241_ = ~new_n7159_ & new_n7240_;
  assign new_n7242_ = ~new_n7235_ & ~new_n7241_;
  assign new_n7243_ = ~\b[23]  & ~new_n7242_;
  assign new_n7244_ = ~new_n6831_ & ~\quotient[33] ;
  assign new_n7245_ = ~new_n6841_ & new_n7112_;
  assign new_n7246_ = ~new_n7108_ & new_n7245_;
  assign new_n7247_ = ~new_n7109_ & ~new_n7112_;
  assign new_n7248_ = ~new_n7246_ & ~new_n7247_;
  assign new_n7249_ = new_n7162_ & ~new_n7248_;
  assign new_n7250_ = ~new_n7159_ & new_n7249_;
  assign new_n7251_ = ~new_n7244_ & ~new_n7250_;
  assign new_n7252_ = ~\b[22]  & ~new_n7251_;
  assign new_n7253_ = ~new_n6840_ & ~\quotient[33] ;
  assign new_n7254_ = ~new_n6850_ & new_n7107_;
  assign new_n7255_ = ~new_n7103_ & new_n7254_;
  assign new_n7256_ = ~new_n7104_ & ~new_n7107_;
  assign new_n7257_ = ~new_n7255_ & ~new_n7256_;
  assign new_n7258_ = new_n7162_ & ~new_n7257_;
  assign new_n7259_ = ~new_n7159_ & new_n7258_;
  assign new_n7260_ = ~new_n7253_ & ~new_n7259_;
  assign new_n7261_ = ~\b[21]  & ~new_n7260_;
  assign new_n7262_ = ~new_n6849_ & ~\quotient[33] ;
  assign new_n7263_ = ~new_n6859_ & new_n7102_;
  assign new_n7264_ = ~new_n7098_ & new_n7263_;
  assign new_n7265_ = ~new_n7099_ & ~new_n7102_;
  assign new_n7266_ = ~new_n7264_ & ~new_n7265_;
  assign new_n7267_ = new_n7162_ & ~new_n7266_;
  assign new_n7268_ = ~new_n7159_ & new_n7267_;
  assign new_n7269_ = ~new_n7262_ & ~new_n7268_;
  assign new_n7270_ = ~\b[20]  & ~new_n7269_;
  assign new_n7271_ = ~new_n6858_ & ~\quotient[33] ;
  assign new_n7272_ = ~new_n6868_ & new_n7097_;
  assign new_n7273_ = ~new_n7093_ & new_n7272_;
  assign new_n7274_ = ~new_n7094_ & ~new_n7097_;
  assign new_n7275_ = ~new_n7273_ & ~new_n7274_;
  assign new_n7276_ = new_n7162_ & ~new_n7275_;
  assign new_n7277_ = ~new_n7159_ & new_n7276_;
  assign new_n7278_ = ~new_n7271_ & ~new_n7277_;
  assign new_n7279_ = ~\b[19]  & ~new_n7278_;
  assign new_n7280_ = ~new_n6867_ & ~\quotient[33] ;
  assign new_n7281_ = ~new_n6877_ & new_n7092_;
  assign new_n7282_ = ~new_n7088_ & new_n7281_;
  assign new_n7283_ = ~new_n7089_ & ~new_n7092_;
  assign new_n7284_ = ~new_n7282_ & ~new_n7283_;
  assign new_n7285_ = new_n7162_ & ~new_n7284_;
  assign new_n7286_ = ~new_n7159_ & new_n7285_;
  assign new_n7287_ = ~new_n7280_ & ~new_n7286_;
  assign new_n7288_ = ~\b[18]  & ~new_n7287_;
  assign new_n7289_ = ~new_n6876_ & ~\quotient[33] ;
  assign new_n7290_ = ~new_n6886_ & new_n7087_;
  assign new_n7291_ = ~new_n7083_ & new_n7290_;
  assign new_n7292_ = ~new_n7084_ & ~new_n7087_;
  assign new_n7293_ = ~new_n7291_ & ~new_n7292_;
  assign new_n7294_ = new_n7162_ & ~new_n7293_;
  assign new_n7295_ = ~new_n7159_ & new_n7294_;
  assign new_n7296_ = ~new_n7289_ & ~new_n7295_;
  assign new_n7297_ = ~\b[17]  & ~new_n7296_;
  assign new_n7298_ = ~new_n6885_ & ~\quotient[33] ;
  assign new_n7299_ = ~new_n6895_ & new_n7082_;
  assign new_n7300_ = ~new_n7078_ & new_n7299_;
  assign new_n7301_ = ~new_n7079_ & ~new_n7082_;
  assign new_n7302_ = ~new_n7300_ & ~new_n7301_;
  assign new_n7303_ = new_n7162_ & ~new_n7302_;
  assign new_n7304_ = ~new_n7159_ & new_n7303_;
  assign new_n7305_ = ~new_n7298_ & ~new_n7304_;
  assign new_n7306_ = ~\b[16]  & ~new_n7305_;
  assign new_n7307_ = ~new_n6894_ & ~\quotient[33] ;
  assign new_n7308_ = ~new_n6904_ & new_n7077_;
  assign new_n7309_ = ~new_n7073_ & new_n7308_;
  assign new_n7310_ = ~new_n7074_ & ~new_n7077_;
  assign new_n7311_ = ~new_n7309_ & ~new_n7310_;
  assign new_n7312_ = new_n7162_ & ~new_n7311_;
  assign new_n7313_ = ~new_n7159_ & new_n7312_;
  assign new_n7314_ = ~new_n7307_ & ~new_n7313_;
  assign new_n7315_ = ~\b[15]  & ~new_n7314_;
  assign new_n7316_ = ~new_n6903_ & ~\quotient[33] ;
  assign new_n7317_ = ~new_n6913_ & new_n7072_;
  assign new_n7318_ = ~new_n7068_ & new_n7317_;
  assign new_n7319_ = ~new_n7069_ & ~new_n7072_;
  assign new_n7320_ = ~new_n7318_ & ~new_n7319_;
  assign new_n7321_ = new_n7162_ & ~new_n7320_;
  assign new_n7322_ = ~new_n7159_ & new_n7321_;
  assign new_n7323_ = ~new_n7316_ & ~new_n7322_;
  assign new_n7324_ = ~\b[14]  & ~new_n7323_;
  assign new_n7325_ = ~new_n6912_ & ~\quotient[33] ;
  assign new_n7326_ = ~new_n6922_ & new_n7067_;
  assign new_n7327_ = ~new_n7063_ & new_n7326_;
  assign new_n7328_ = ~new_n7064_ & ~new_n7067_;
  assign new_n7329_ = ~new_n7327_ & ~new_n7328_;
  assign new_n7330_ = new_n7162_ & ~new_n7329_;
  assign new_n7331_ = ~new_n7159_ & new_n7330_;
  assign new_n7332_ = ~new_n7325_ & ~new_n7331_;
  assign new_n7333_ = ~\b[13]  & ~new_n7332_;
  assign new_n7334_ = ~new_n6921_ & ~\quotient[33] ;
  assign new_n7335_ = ~new_n6931_ & new_n7062_;
  assign new_n7336_ = ~new_n7058_ & new_n7335_;
  assign new_n7337_ = ~new_n7059_ & ~new_n7062_;
  assign new_n7338_ = ~new_n7336_ & ~new_n7337_;
  assign new_n7339_ = new_n7162_ & ~new_n7338_;
  assign new_n7340_ = ~new_n7159_ & new_n7339_;
  assign new_n7341_ = ~new_n7334_ & ~new_n7340_;
  assign new_n7342_ = ~\b[12]  & ~new_n7341_;
  assign new_n7343_ = ~new_n6930_ & ~\quotient[33] ;
  assign new_n7344_ = ~new_n6940_ & new_n7057_;
  assign new_n7345_ = ~new_n7053_ & new_n7344_;
  assign new_n7346_ = ~new_n7054_ & ~new_n7057_;
  assign new_n7347_ = ~new_n7345_ & ~new_n7346_;
  assign new_n7348_ = new_n7162_ & ~new_n7347_;
  assign new_n7349_ = ~new_n7159_ & new_n7348_;
  assign new_n7350_ = ~new_n7343_ & ~new_n7349_;
  assign new_n7351_ = ~\b[11]  & ~new_n7350_;
  assign new_n7352_ = ~new_n6939_ & ~\quotient[33] ;
  assign new_n7353_ = ~new_n6949_ & new_n7052_;
  assign new_n7354_ = ~new_n7048_ & new_n7353_;
  assign new_n7355_ = ~new_n7049_ & ~new_n7052_;
  assign new_n7356_ = ~new_n7354_ & ~new_n7355_;
  assign new_n7357_ = new_n7162_ & ~new_n7356_;
  assign new_n7358_ = ~new_n7159_ & new_n7357_;
  assign new_n7359_ = ~new_n7352_ & ~new_n7358_;
  assign new_n7360_ = ~\b[10]  & ~new_n7359_;
  assign new_n7361_ = ~new_n6948_ & ~\quotient[33] ;
  assign new_n7362_ = ~new_n6958_ & new_n7047_;
  assign new_n7363_ = ~new_n7043_ & new_n7362_;
  assign new_n7364_ = ~new_n7044_ & ~new_n7047_;
  assign new_n7365_ = ~new_n7363_ & ~new_n7364_;
  assign new_n7366_ = new_n7162_ & ~new_n7365_;
  assign new_n7367_ = ~new_n7159_ & new_n7366_;
  assign new_n7368_ = ~new_n7361_ & ~new_n7367_;
  assign new_n7369_ = ~\b[9]  & ~new_n7368_;
  assign new_n7370_ = ~new_n6957_ & ~\quotient[33] ;
  assign new_n7371_ = ~new_n6967_ & new_n7042_;
  assign new_n7372_ = ~new_n7038_ & new_n7371_;
  assign new_n7373_ = ~new_n7039_ & ~new_n7042_;
  assign new_n7374_ = ~new_n7372_ & ~new_n7373_;
  assign new_n7375_ = new_n7162_ & ~new_n7374_;
  assign new_n7376_ = ~new_n7159_ & new_n7375_;
  assign new_n7377_ = ~new_n7370_ & ~new_n7376_;
  assign new_n7378_ = ~\b[8]  & ~new_n7377_;
  assign new_n7379_ = ~new_n6966_ & ~\quotient[33] ;
  assign new_n7380_ = ~new_n6976_ & new_n7037_;
  assign new_n7381_ = ~new_n7033_ & new_n7380_;
  assign new_n7382_ = ~new_n7034_ & ~new_n7037_;
  assign new_n7383_ = ~new_n7381_ & ~new_n7382_;
  assign new_n7384_ = new_n7162_ & ~new_n7383_;
  assign new_n7385_ = ~new_n7159_ & new_n7384_;
  assign new_n7386_ = ~new_n7379_ & ~new_n7385_;
  assign new_n7387_ = ~\b[7]  & ~new_n7386_;
  assign new_n7388_ = ~new_n6975_ & ~\quotient[33] ;
  assign new_n7389_ = ~new_n6985_ & new_n7032_;
  assign new_n7390_ = ~new_n7028_ & new_n7389_;
  assign new_n7391_ = ~new_n7029_ & ~new_n7032_;
  assign new_n7392_ = ~new_n7390_ & ~new_n7391_;
  assign new_n7393_ = new_n7162_ & ~new_n7392_;
  assign new_n7394_ = ~new_n7159_ & new_n7393_;
  assign new_n7395_ = ~new_n7388_ & ~new_n7394_;
  assign new_n7396_ = ~\b[6]  & ~new_n7395_;
  assign new_n7397_ = ~new_n6984_ & ~\quotient[33] ;
  assign new_n7398_ = ~new_n6994_ & new_n7027_;
  assign new_n7399_ = ~new_n7023_ & new_n7398_;
  assign new_n7400_ = ~new_n7024_ & ~new_n7027_;
  assign new_n7401_ = ~new_n7399_ & ~new_n7400_;
  assign new_n7402_ = new_n7162_ & ~new_n7401_;
  assign new_n7403_ = ~new_n7159_ & new_n7402_;
  assign new_n7404_ = ~new_n7397_ & ~new_n7403_;
  assign new_n7405_ = ~\b[5]  & ~new_n7404_;
  assign new_n7406_ = ~new_n6993_ & ~\quotient[33] ;
  assign new_n7407_ = ~new_n7002_ & new_n7022_;
  assign new_n7408_ = ~new_n7018_ & new_n7407_;
  assign new_n7409_ = ~new_n7019_ & ~new_n7022_;
  assign new_n7410_ = ~new_n7408_ & ~new_n7409_;
  assign new_n7411_ = new_n7162_ & ~new_n7410_;
  assign new_n7412_ = ~new_n7159_ & new_n7411_;
  assign new_n7413_ = ~new_n7406_ & ~new_n7412_;
  assign new_n7414_ = ~\b[4]  & ~new_n7413_;
  assign new_n7415_ = ~new_n7001_ & ~\quotient[33] ;
  assign new_n7416_ = ~new_n7013_ & new_n7017_;
  assign new_n7417_ = ~new_n7012_ & new_n7416_;
  assign new_n7418_ = ~new_n7014_ & ~new_n7017_;
  assign new_n7419_ = ~new_n7417_ & ~new_n7418_;
  assign new_n7420_ = new_n7162_ & ~new_n7419_;
  assign new_n7421_ = ~new_n7159_ & new_n7420_;
  assign new_n7422_ = ~new_n7415_ & ~new_n7421_;
  assign new_n7423_ = ~\b[3]  & ~new_n7422_;
  assign new_n7424_ = ~new_n7006_ & ~\quotient[33] ;
  assign new_n7425_ = ~new_n7009_ & new_n7011_;
  assign new_n7426_ = ~new_n7007_ & new_n7425_;
  assign new_n7427_ = new_n7162_ & ~new_n7426_;
  assign new_n7428_ = ~new_n7012_ & new_n7427_;
  assign new_n7429_ = ~new_n7159_ & new_n7428_;
  assign new_n7430_ = ~new_n7424_ & ~new_n7429_;
  assign new_n7431_ = ~\b[2]  & ~new_n7430_;
  assign new_n7432_ = \b[0]  & ~\b[31] ;
  assign new_n7433_ = new_n313_ & new_n7432_;
  assign new_n7434_ = new_n303_ & new_n7433_;
  assign new_n7435_ = new_n288_ & new_n7434_;
  assign new_n7436_ = ~new_n7159_ & new_n7435_;
  assign new_n7437_ = \a[33]  & ~new_n7436_;
  assign new_n7438_ = new_n372_ & new_n7011_;
  assign new_n7439_ = new_n414_ & new_n7438_;
  assign new_n7440_ = new_n598_ & new_n7439_;
  assign new_n7441_ = new_n595_ & new_n7440_;
  assign new_n7442_ = ~new_n7159_ & new_n7441_;
  assign new_n7443_ = ~new_n7437_ & ~new_n7442_;
  assign new_n7444_ = \b[1]  & ~new_n7443_;
  assign new_n7445_ = ~\b[1]  & ~new_n7442_;
  assign new_n7446_ = ~new_n7437_ & new_n7445_;
  assign new_n7447_ = ~new_n7444_ & ~new_n7446_;
  assign new_n7448_ = ~\a[32]  & \b[0] ;
  assign new_n7449_ = ~new_n7447_ & ~new_n7448_;
  assign new_n7450_ = ~\b[1]  & ~new_n7443_;
  assign new_n7451_ = ~new_n7449_ & ~new_n7450_;
  assign new_n7452_ = \b[2]  & ~new_n7429_;
  assign new_n7453_ = ~new_n7424_ & new_n7452_;
  assign new_n7454_ = ~new_n7431_ & ~new_n7453_;
  assign new_n7455_ = ~new_n7451_ & new_n7454_;
  assign new_n7456_ = ~new_n7431_ & ~new_n7455_;
  assign new_n7457_ = \b[3]  & ~new_n7421_;
  assign new_n7458_ = ~new_n7415_ & new_n7457_;
  assign new_n7459_ = ~new_n7423_ & ~new_n7458_;
  assign new_n7460_ = ~new_n7456_ & new_n7459_;
  assign new_n7461_ = ~new_n7423_ & ~new_n7460_;
  assign new_n7462_ = \b[4]  & ~new_n7412_;
  assign new_n7463_ = ~new_n7406_ & new_n7462_;
  assign new_n7464_ = ~new_n7414_ & ~new_n7463_;
  assign new_n7465_ = ~new_n7461_ & new_n7464_;
  assign new_n7466_ = ~new_n7414_ & ~new_n7465_;
  assign new_n7467_ = \b[5]  & ~new_n7403_;
  assign new_n7468_ = ~new_n7397_ & new_n7467_;
  assign new_n7469_ = ~new_n7405_ & ~new_n7468_;
  assign new_n7470_ = ~new_n7466_ & new_n7469_;
  assign new_n7471_ = ~new_n7405_ & ~new_n7470_;
  assign new_n7472_ = \b[6]  & ~new_n7394_;
  assign new_n7473_ = ~new_n7388_ & new_n7472_;
  assign new_n7474_ = ~new_n7396_ & ~new_n7473_;
  assign new_n7475_ = ~new_n7471_ & new_n7474_;
  assign new_n7476_ = ~new_n7396_ & ~new_n7475_;
  assign new_n7477_ = \b[7]  & ~new_n7385_;
  assign new_n7478_ = ~new_n7379_ & new_n7477_;
  assign new_n7479_ = ~new_n7387_ & ~new_n7478_;
  assign new_n7480_ = ~new_n7476_ & new_n7479_;
  assign new_n7481_ = ~new_n7387_ & ~new_n7480_;
  assign new_n7482_ = \b[8]  & ~new_n7376_;
  assign new_n7483_ = ~new_n7370_ & new_n7482_;
  assign new_n7484_ = ~new_n7378_ & ~new_n7483_;
  assign new_n7485_ = ~new_n7481_ & new_n7484_;
  assign new_n7486_ = ~new_n7378_ & ~new_n7485_;
  assign new_n7487_ = \b[9]  & ~new_n7367_;
  assign new_n7488_ = ~new_n7361_ & new_n7487_;
  assign new_n7489_ = ~new_n7369_ & ~new_n7488_;
  assign new_n7490_ = ~new_n7486_ & new_n7489_;
  assign new_n7491_ = ~new_n7369_ & ~new_n7490_;
  assign new_n7492_ = \b[10]  & ~new_n7358_;
  assign new_n7493_ = ~new_n7352_ & new_n7492_;
  assign new_n7494_ = ~new_n7360_ & ~new_n7493_;
  assign new_n7495_ = ~new_n7491_ & new_n7494_;
  assign new_n7496_ = ~new_n7360_ & ~new_n7495_;
  assign new_n7497_ = \b[11]  & ~new_n7349_;
  assign new_n7498_ = ~new_n7343_ & new_n7497_;
  assign new_n7499_ = ~new_n7351_ & ~new_n7498_;
  assign new_n7500_ = ~new_n7496_ & new_n7499_;
  assign new_n7501_ = ~new_n7351_ & ~new_n7500_;
  assign new_n7502_ = \b[12]  & ~new_n7340_;
  assign new_n7503_ = ~new_n7334_ & new_n7502_;
  assign new_n7504_ = ~new_n7342_ & ~new_n7503_;
  assign new_n7505_ = ~new_n7501_ & new_n7504_;
  assign new_n7506_ = ~new_n7342_ & ~new_n7505_;
  assign new_n7507_ = \b[13]  & ~new_n7331_;
  assign new_n7508_ = ~new_n7325_ & new_n7507_;
  assign new_n7509_ = ~new_n7333_ & ~new_n7508_;
  assign new_n7510_ = ~new_n7506_ & new_n7509_;
  assign new_n7511_ = ~new_n7333_ & ~new_n7510_;
  assign new_n7512_ = \b[14]  & ~new_n7322_;
  assign new_n7513_ = ~new_n7316_ & new_n7512_;
  assign new_n7514_ = ~new_n7324_ & ~new_n7513_;
  assign new_n7515_ = ~new_n7511_ & new_n7514_;
  assign new_n7516_ = ~new_n7324_ & ~new_n7515_;
  assign new_n7517_ = \b[15]  & ~new_n7313_;
  assign new_n7518_ = ~new_n7307_ & new_n7517_;
  assign new_n7519_ = ~new_n7315_ & ~new_n7518_;
  assign new_n7520_ = ~new_n7516_ & new_n7519_;
  assign new_n7521_ = ~new_n7315_ & ~new_n7520_;
  assign new_n7522_ = \b[16]  & ~new_n7304_;
  assign new_n7523_ = ~new_n7298_ & new_n7522_;
  assign new_n7524_ = ~new_n7306_ & ~new_n7523_;
  assign new_n7525_ = ~new_n7521_ & new_n7524_;
  assign new_n7526_ = ~new_n7306_ & ~new_n7525_;
  assign new_n7527_ = \b[17]  & ~new_n7295_;
  assign new_n7528_ = ~new_n7289_ & new_n7527_;
  assign new_n7529_ = ~new_n7297_ & ~new_n7528_;
  assign new_n7530_ = ~new_n7526_ & new_n7529_;
  assign new_n7531_ = ~new_n7297_ & ~new_n7530_;
  assign new_n7532_ = \b[18]  & ~new_n7286_;
  assign new_n7533_ = ~new_n7280_ & new_n7532_;
  assign new_n7534_ = ~new_n7288_ & ~new_n7533_;
  assign new_n7535_ = ~new_n7531_ & new_n7534_;
  assign new_n7536_ = ~new_n7288_ & ~new_n7535_;
  assign new_n7537_ = \b[19]  & ~new_n7277_;
  assign new_n7538_ = ~new_n7271_ & new_n7537_;
  assign new_n7539_ = ~new_n7279_ & ~new_n7538_;
  assign new_n7540_ = ~new_n7536_ & new_n7539_;
  assign new_n7541_ = ~new_n7279_ & ~new_n7540_;
  assign new_n7542_ = \b[20]  & ~new_n7268_;
  assign new_n7543_ = ~new_n7262_ & new_n7542_;
  assign new_n7544_ = ~new_n7270_ & ~new_n7543_;
  assign new_n7545_ = ~new_n7541_ & new_n7544_;
  assign new_n7546_ = ~new_n7270_ & ~new_n7545_;
  assign new_n7547_ = \b[21]  & ~new_n7259_;
  assign new_n7548_ = ~new_n7253_ & new_n7547_;
  assign new_n7549_ = ~new_n7261_ & ~new_n7548_;
  assign new_n7550_ = ~new_n7546_ & new_n7549_;
  assign new_n7551_ = ~new_n7261_ & ~new_n7550_;
  assign new_n7552_ = \b[22]  & ~new_n7250_;
  assign new_n7553_ = ~new_n7244_ & new_n7552_;
  assign new_n7554_ = ~new_n7252_ & ~new_n7553_;
  assign new_n7555_ = ~new_n7551_ & new_n7554_;
  assign new_n7556_ = ~new_n7252_ & ~new_n7555_;
  assign new_n7557_ = \b[23]  & ~new_n7241_;
  assign new_n7558_ = ~new_n7235_ & new_n7557_;
  assign new_n7559_ = ~new_n7243_ & ~new_n7558_;
  assign new_n7560_ = ~new_n7556_ & new_n7559_;
  assign new_n7561_ = ~new_n7243_ & ~new_n7560_;
  assign new_n7562_ = \b[24]  & ~new_n7232_;
  assign new_n7563_ = ~new_n7226_ & new_n7562_;
  assign new_n7564_ = ~new_n7234_ & ~new_n7563_;
  assign new_n7565_ = ~new_n7561_ & new_n7564_;
  assign new_n7566_ = ~new_n7234_ & ~new_n7565_;
  assign new_n7567_ = \b[25]  & ~new_n7223_;
  assign new_n7568_ = ~new_n7217_ & new_n7567_;
  assign new_n7569_ = ~new_n7225_ & ~new_n7568_;
  assign new_n7570_ = ~new_n7566_ & new_n7569_;
  assign new_n7571_ = ~new_n7225_ & ~new_n7570_;
  assign new_n7572_ = \b[26]  & ~new_n7214_;
  assign new_n7573_ = ~new_n7208_ & new_n7572_;
  assign new_n7574_ = ~new_n7216_ & ~new_n7573_;
  assign new_n7575_ = ~new_n7571_ & new_n7574_;
  assign new_n7576_ = ~new_n7216_ & ~new_n7575_;
  assign new_n7577_ = \b[27]  & ~new_n7205_;
  assign new_n7578_ = ~new_n7199_ & new_n7577_;
  assign new_n7579_ = ~new_n7207_ & ~new_n7578_;
  assign new_n7580_ = ~new_n7576_ & new_n7579_;
  assign new_n7581_ = ~new_n7207_ & ~new_n7580_;
  assign new_n7582_ = \b[28]  & ~new_n7196_;
  assign new_n7583_ = ~new_n7190_ & new_n7582_;
  assign new_n7584_ = ~new_n7198_ & ~new_n7583_;
  assign new_n7585_ = ~new_n7581_ & new_n7584_;
  assign new_n7586_ = ~new_n7198_ & ~new_n7585_;
  assign new_n7587_ = \b[29]  & ~new_n7187_;
  assign new_n7588_ = ~new_n7181_ & new_n7587_;
  assign new_n7589_ = ~new_n7189_ & ~new_n7588_;
  assign new_n7590_ = ~new_n7586_ & new_n7589_;
  assign new_n7591_ = ~new_n7189_ & ~new_n7590_;
  assign new_n7592_ = \b[30]  & ~new_n7170_;
  assign new_n7593_ = ~new_n7164_ & new_n7592_;
  assign new_n7594_ = ~new_n7180_ & ~new_n7593_;
  assign new_n7595_ = ~new_n7591_ & new_n7594_;
  assign new_n7596_ = ~new_n7180_ & ~new_n7595_;
  assign new_n7597_ = \b[31]  & ~new_n7172_;
  assign new_n7598_ = ~new_n7177_ & new_n7597_;
  assign new_n7599_ = ~new_n7179_ & ~new_n7598_;
  assign new_n7600_ = ~new_n7596_ & new_n7599_;
  assign new_n7601_ = ~new_n7179_ & ~new_n7600_;
  assign \quotient[32]  = new_n432_ & ~new_n7601_;
  assign new_n7603_ = ~new_n7171_ & ~\quotient[32] ;
  assign new_n7604_ = ~new_n7189_ & new_n7594_;
  assign new_n7605_ = ~new_n7590_ & new_n7604_;
  assign new_n7606_ = ~new_n7591_ & ~new_n7594_;
  assign new_n7607_ = ~new_n7605_ & ~new_n7606_;
  assign new_n7608_ = new_n432_ & ~new_n7607_;
  assign new_n7609_ = ~new_n7601_ & new_n7608_;
  assign new_n7610_ = ~new_n7603_ & ~new_n7609_;
  assign new_n7611_ = ~\b[31]  & ~new_n7610_;
  assign new_n7612_ = ~new_n7188_ & ~\quotient[32] ;
  assign new_n7613_ = ~new_n7198_ & new_n7589_;
  assign new_n7614_ = ~new_n7585_ & new_n7613_;
  assign new_n7615_ = ~new_n7586_ & ~new_n7589_;
  assign new_n7616_ = ~new_n7614_ & ~new_n7615_;
  assign new_n7617_ = new_n432_ & ~new_n7616_;
  assign new_n7618_ = ~new_n7601_ & new_n7617_;
  assign new_n7619_ = ~new_n7612_ & ~new_n7618_;
  assign new_n7620_ = ~\b[30]  & ~new_n7619_;
  assign new_n7621_ = ~new_n7197_ & ~\quotient[32] ;
  assign new_n7622_ = ~new_n7207_ & new_n7584_;
  assign new_n7623_ = ~new_n7580_ & new_n7622_;
  assign new_n7624_ = ~new_n7581_ & ~new_n7584_;
  assign new_n7625_ = ~new_n7623_ & ~new_n7624_;
  assign new_n7626_ = new_n432_ & ~new_n7625_;
  assign new_n7627_ = ~new_n7601_ & new_n7626_;
  assign new_n7628_ = ~new_n7621_ & ~new_n7627_;
  assign new_n7629_ = ~\b[29]  & ~new_n7628_;
  assign new_n7630_ = ~new_n7206_ & ~\quotient[32] ;
  assign new_n7631_ = ~new_n7216_ & new_n7579_;
  assign new_n7632_ = ~new_n7575_ & new_n7631_;
  assign new_n7633_ = ~new_n7576_ & ~new_n7579_;
  assign new_n7634_ = ~new_n7632_ & ~new_n7633_;
  assign new_n7635_ = new_n432_ & ~new_n7634_;
  assign new_n7636_ = ~new_n7601_ & new_n7635_;
  assign new_n7637_ = ~new_n7630_ & ~new_n7636_;
  assign new_n7638_ = ~\b[28]  & ~new_n7637_;
  assign new_n7639_ = ~new_n7215_ & ~\quotient[32] ;
  assign new_n7640_ = ~new_n7225_ & new_n7574_;
  assign new_n7641_ = ~new_n7570_ & new_n7640_;
  assign new_n7642_ = ~new_n7571_ & ~new_n7574_;
  assign new_n7643_ = ~new_n7641_ & ~new_n7642_;
  assign new_n7644_ = new_n432_ & ~new_n7643_;
  assign new_n7645_ = ~new_n7601_ & new_n7644_;
  assign new_n7646_ = ~new_n7639_ & ~new_n7645_;
  assign new_n7647_ = ~\b[27]  & ~new_n7646_;
  assign new_n7648_ = ~new_n7224_ & ~\quotient[32] ;
  assign new_n7649_ = ~new_n7234_ & new_n7569_;
  assign new_n7650_ = ~new_n7565_ & new_n7649_;
  assign new_n7651_ = ~new_n7566_ & ~new_n7569_;
  assign new_n7652_ = ~new_n7650_ & ~new_n7651_;
  assign new_n7653_ = new_n432_ & ~new_n7652_;
  assign new_n7654_ = ~new_n7601_ & new_n7653_;
  assign new_n7655_ = ~new_n7648_ & ~new_n7654_;
  assign new_n7656_ = ~\b[26]  & ~new_n7655_;
  assign new_n7657_ = ~new_n7233_ & ~\quotient[32] ;
  assign new_n7658_ = ~new_n7243_ & new_n7564_;
  assign new_n7659_ = ~new_n7560_ & new_n7658_;
  assign new_n7660_ = ~new_n7561_ & ~new_n7564_;
  assign new_n7661_ = ~new_n7659_ & ~new_n7660_;
  assign new_n7662_ = new_n432_ & ~new_n7661_;
  assign new_n7663_ = ~new_n7601_ & new_n7662_;
  assign new_n7664_ = ~new_n7657_ & ~new_n7663_;
  assign new_n7665_ = ~\b[25]  & ~new_n7664_;
  assign new_n7666_ = ~new_n7242_ & ~\quotient[32] ;
  assign new_n7667_ = ~new_n7252_ & new_n7559_;
  assign new_n7668_ = ~new_n7555_ & new_n7667_;
  assign new_n7669_ = ~new_n7556_ & ~new_n7559_;
  assign new_n7670_ = ~new_n7668_ & ~new_n7669_;
  assign new_n7671_ = new_n432_ & ~new_n7670_;
  assign new_n7672_ = ~new_n7601_ & new_n7671_;
  assign new_n7673_ = ~new_n7666_ & ~new_n7672_;
  assign new_n7674_ = ~\b[24]  & ~new_n7673_;
  assign new_n7675_ = ~new_n7251_ & ~\quotient[32] ;
  assign new_n7676_ = ~new_n7261_ & new_n7554_;
  assign new_n7677_ = ~new_n7550_ & new_n7676_;
  assign new_n7678_ = ~new_n7551_ & ~new_n7554_;
  assign new_n7679_ = ~new_n7677_ & ~new_n7678_;
  assign new_n7680_ = new_n432_ & ~new_n7679_;
  assign new_n7681_ = ~new_n7601_ & new_n7680_;
  assign new_n7682_ = ~new_n7675_ & ~new_n7681_;
  assign new_n7683_ = ~\b[23]  & ~new_n7682_;
  assign new_n7684_ = ~new_n7260_ & ~\quotient[32] ;
  assign new_n7685_ = ~new_n7270_ & new_n7549_;
  assign new_n7686_ = ~new_n7545_ & new_n7685_;
  assign new_n7687_ = ~new_n7546_ & ~new_n7549_;
  assign new_n7688_ = ~new_n7686_ & ~new_n7687_;
  assign new_n7689_ = new_n432_ & ~new_n7688_;
  assign new_n7690_ = ~new_n7601_ & new_n7689_;
  assign new_n7691_ = ~new_n7684_ & ~new_n7690_;
  assign new_n7692_ = ~\b[22]  & ~new_n7691_;
  assign new_n7693_ = ~new_n7269_ & ~\quotient[32] ;
  assign new_n7694_ = ~new_n7279_ & new_n7544_;
  assign new_n7695_ = ~new_n7540_ & new_n7694_;
  assign new_n7696_ = ~new_n7541_ & ~new_n7544_;
  assign new_n7697_ = ~new_n7695_ & ~new_n7696_;
  assign new_n7698_ = new_n432_ & ~new_n7697_;
  assign new_n7699_ = ~new_n7601_ & new_n7698_;
  assign new_n7700_ = ~new_n7693_ & ~new_n7699_;
  assign new_n7701_ = ~\b[21]  & ~new_n7700_;
  assign new_n7702_ = ~new_n7278_ & ~\quotient[32] ;
  assign new_n7703_ = ~new_n7288_ & new_n7539_;
  assign new_n7704_ = ~new_n7535_ & new_n7703_;
  assign new_n7705_ = ~new_n7536_ & ~new_n7539_;
  assign new_n7706_ = ~new_n7704_ & ~new_n7705_;
  assign new_n7707_ = new_n432_ & ~new_n7706_;
  assign new_n7708_ = ~new_n7601_ & new_n7707_;
  assign new_n7709_ = ~new_n7702_ & ~new_n7708_;
  assign new_n7710_ = ~\b[20]  & ~new_n7709_;
  assign new_n7711_ = ~new_n7287_ & ~\quotient[32] ;
  assign new_n7712_ = ~new_n7297_ & new_n7534_;
  assign new_n7713_ = ~new_n7530_ & new_n7712_;
  assign new_n7714_ = ~new_n7531_ & ~new_n7534_;
  assign new_n7715_ = ~new_n7713_ & ~new_n7714_;
  assign new_n7716_ = new_n432_ & ~new_n7715_;
  assign new_n7717_ = ~new_n7601_ & new_n7716_;
  assign new_n7718_ = ~new_n7711_ & ~new_n7717_;
  assign new_n7719_ = ~\b[19]  & ~new_n7718_;
  assign new_n7720_ = ~new_n7296_ & ~\quotient[32] ;
  assign new_n7721_ = ~new_n7306_ & new_n7529_;
  assign new_n7722_ = ~new_n7525_ & new_n7721_;
  assign new_n7723_ = ~new_n7526_ & ~new_n7529_;
  assign new_n7724_ = ~new_n7722_ & ~new_n7723_;
  assign new_n7725_ = new_n432_ & ~new_n7724_;
  assign new_n7726_ = ~new_n7601_ & new_n7725_;
  assign new_n7727_ = ~new_n7720_ & ~new_n7726_;
  assign new_n7728_ = ~\b[18]  & ~new_n7727_;
  assign new_n7729_ = ~new_n7305_ & ~\quotient[32] ;
  assign new_n7730_ = ~new_n7315_ & new_n7524_;
  assign new_n7731_ = ~new_n7520_ & new_n7730_;
  assign new_n7732_ = ~new_n7521_ & ~new_n7524_;
  assign new_n7733_ = ~new_n7731_ & ~new_n7732_;
  assign new_n7734_ = new_n432_ & ~new_n7733_;
  assign new_n7735_ = ~new_n7601_ & new_n7734_;
  assign new_n7736_ = ~new_n7729_ & ~new_n7735_;
  assign new_n7737_ = ~\b[17]  & ~new_n7736_;
  assign new_n7738_ = ~new_n7314_ & ~\quotient[32] ;
  assign new_n7739_ = ~new_n7324_ & new_n7519_;
  assign new_n7740_ = ~new_n7515_ & new_n7739_;
  assign new_n7741_ = ~new_n7516_ & ~new_n7519_;
  assign new_n7742_ = ~new_n7740_ & ~new_n7741_;
  assign new_n7743_ = new_n432_ & ~new_n7742_;
  assign new_n7744_ = ~new_n7601_ & new_n7743_;
  assign new_n7745_ = ~new_n7738_ & ~new_n7744_;
  assign new_n7746_ = ~\b[16]  & ~new_n7745_;
  assign new_n7747_ = ~new_n7323_ & ~\quotient[32] ;
  assign new_n7748_ = ~new_n7333_ & new_n7514_;
  assign new_n7749_ = ~new_n7510_ & new_n7748_;
  assign new_n7750_ = ~new_n7511_ & ~new_n7514_;
  assign new_n7751_ = ~new_n7749_ & ~new_n7750_;
  assign new_n7752_ = new_n432_ & ~new_n7751_;
  assign new_n7753_ = ~new_n7601_ & new_n7752_;
  assign new_n7754_ = ~new_n7747_ & ~new_n7753_;
  assign new_n7755_ = ~\b[15]  & ~new_n7754_;
  assign new_n7756_ = ~new_n7332_ & ~\quotient[32] ;
  assign new_n7757_ = ~new_n7342_ & new_n7509_;
  assign new_n7758_ = ~new_n7505_ & new_n7757_;
  assign new_n7759_ = ~new_n7506_ & ~new_n7509_;
  assign new_n7760_ = ~new_n7758_ & ~new_n7759_;
  assign new_n7761_ = new_n432_ & ~new_n7760_;
  assign new_n7762_ = ~new_n7601_ & new_n7761_;
  assign new_n7763_ = ~new_n7756_ & ~new_n7762_;
  assign new_n7764_ = ~\b[14]  & ~new_n7763_;
  assign new_n7765_ = ~new_n7341_ & ~\quotient[32] ;
  assign new_n7766_ = ~new_n7351_ & new_n7504_;
  assign new_n7767_ = ~new_n7500_ & new_n7766_;
  assign new_n7768_ = ~new_n7501_ & ~new_n7504_;
  assign new_n7769_ = ~new_n7767_ & ~new_n7768_;
  assign new_n7770_ = new_n432_ & ~new_n7769_;
  assign new_n7771_ = ~new_n7601_ & new_n7770_;
  assign new_n7772_ = ~new_n7765_ & ~new_n7771_;
  assign new_n7773_ = ~\b[13]  & ~new_n7772_;
  assign new_n7774_ = ~new_n7350_ & ~\quotient[32] ;
  assign new_n7775_ = ~new_n7360_ & new_n7499_;
  assign new_n7776_ = ~new_n7495_ & new_n7775_;
  assign new_n7777_ = ~new_n7496_ & ~new_n7499_;
  assign new_n7778_ = ~new_n7776_ & ~new_n7777_;
  assign new_n7779_ = new_n432_ & ~new_n7778_;
  assign new_n7780_ = ~new_n7601_ & new_n7779_;
  assign new_n7781_ = ~new_n7774_ & ~new_n7780_;
  assign new_n7782_ = ~\b[12]  & ~new_n7781_;
  assign new_n7783_ = ~new_n7359_ & ~\quotient[32] ;
  assign new_n7784_ = ~new_n7369_ & new_n7494_;
  assign new_n7785_ = ~new_n7490_ & new_n7784_;
  assign new_n7786_ = ~new_n7491_ & ~new_n7494_;
  assign new_n7787_ = ~new_n7785_ & ~new_n7786_;
  assign new_n7788_ = new_n432_ & ~new_n7787_;
  assign new_n7789_ = ~new_n7601_ & new_n7788_;
  assign new_n7790_ = ~new_n7783_ & ~new_n7789_;
  assign new_n7791_ = ~\b[11]  & ~new_n7790_;
  assign new_n7792_ = ~new_n7368_ & ~\quotient[32] ;
  assign new_n7793_ = ~new_n7378_ & new_n7489_;
  assign new_n7794_ = ~new_n7485_ & new_n7793_;
  assign new_n7795_ = ~new_n7486_ & ~new_n7489_;
  assign new_n7796_ = ~new_n7794_ & ~new_n7795_;
  assign new_n7797_ = new_n432_ & ~new_n7796_;
  assign new_n7798_ = ~new_n7601_ & new_n7797_;
  assign new_n7799_ = ~new_n7792_ & ~new_n7798_;
  assign new_n7800_ = ~\b[10]  & ~new_n7799_;
  assign new_n7801_ = ~new_n7377_ & ~\quotient[32] ;
  assign new_n7802_ = ~new_n7387_ & new_n7484_;
  assign new_n7803_ = ~new_n7480_ & new_n7802_;
  assign new_n7804_ = ~new_n7481_ & ~new_n7484_;
  assign new_n7805_ = ~new_n7803_ & ~new_n7804_;
  assign new_n7806_ = new_n432_ & ~new_n7805_;
  assign new_n7807_ = ~new_n7601_ & new_n7806_;
  assign new_n7808_ = ~new_n7801_ & ~new_n7807_;
  assign new_n7809_ = ~\b[9]  & ~new_n7808_;
  assign new_n7810_ = ~new_n7386_ & ~\quotient[32] ;
  assign new_n7811_ = ~new_n7396_ & new_n7479_;
  assign new_n7812_ = ~new_n7475_ & new_n7811_;
  assign new_n7813_ = ~new_n7476_ & ~new_n7479_;
  assign new_n7814_ = ~new_n7812_ & ~new_n7813_;
  assign new_n7815_ = new_n432_ & ~new_n7814_;
  assign new_n7816_ = ~new_n7601_ & new_n7815_;
  assign new_n7817_ = ~new_n7810_ & ~new_n7816_;
  assign new_n7818_ = ~\b[8]  & ~new_n7817_;
  assign new_n7819_ = ~new_n7395_ & ~\quotient[32] ;
  assign new_n7820_ = ~new_n7405_ & new_n7474_;
  assign new_n7821_ = ~new_n7470_ & new_n7820_;
  assign new_n7822_ = ~new_n7471_ & ~new_n7474_;
  assign new_n7823_ = ~new_n7821_ & ~new_n7822_;
  assign new_n7824_ = new_n432_ & ~new_n7823_;
  assign new_n7825_ = ~new_n7601_ & new_n7824_;
  assign new_n7826_ = ~new_n7819_ & ~new_n7825_;
  assign new_n7827_ = ~\b[7]  & ~new_n7826_;
  assign new_n7828_ = ~new_n7404_ & ~\quotient[32] ;
  assign new_n7829_ = ~new_n7414_ & new_n7469_;
  assign new_n7830_ = ~new_n7465_ & new_n7829_;
  assign new_n7831_ = ~new_n7466_ & ~new_n7469_;
  assign new_n7832_ = ~new_n7830_ & ~new_n7831_;
  assign new_n7833_ = new_n432_ & ~new_n7832_;
  assign new_n7834_ = ~new_n7601_ & new_n7833_;
  assign new_n7835_ = ~new_n7828_ & ~new_n7834_;
  assign new_n7836_ = ~\b[6]  & ~new_n7835_;
  assign new_n7837_ = ~new_n7413_ & ~\quotient[32] ;
  assign new_n7838_ = ~new_n7423_ & new_n7464_;
  assign new_n7839_ = ~new_n7460_ & new_n7838_;
  assign new_n7840_ = ~new_n7461_ & ~new_n7464_;
  assign new_n7841_ = ~new_n7839_ & ~new_n7840_;
  assign new_n7842_ = new_n432_ & ~new_n7841_;
  assign new_n7843_ = ~new_n7601_ & new_n7842_;
  assign new_n7844_ = ~new_n7837_ & ~new_n7843_;
  assign new_n7845_ = ~\b[5]  & ~new_n7844_;
  assign new_n7846_ = ~new_n7422_ & ~\quotient[32] ;
  assign new_n7847_ = ~new_n7431_ & new_n7459_;
  assign new_n7848_ = ~new_n7455_ & new_n7847_;
  assign new_n7849_ = ~new_n7456_ & ~new_n7459_;
  assign new_n7850_ = ~new_n7848_ & ~new_n7849_;
  assign new_n7851_ = new_n432_ & ~new_n7850_;
  assign new_n7852_ = ~new_n7601_ & new_n7851_;
  assign new_n7853_ = ~new_n7846_ & ~new_n7852_;
  assign new_n7854_ = ~\b[4]  & ~new_n7853_;
  assign new_n7855_ = ~new_n7430_ & ~\quotient[32] ;
  assign new_n7856_ = ~new_n7450_ & new_n7454_;
  assign new_n7857_ = ~new_n7449_ & new_n7856_;
  assign new_n7858_ = ~new_n7451_ & ~new_n7454_;
  assign new_n7859_ = ~new_n7857_ & ~new_n7858_;
  assign new_n7860_ = new_n432_ & ~new_n7859_;
  assign new_n7861_ = ~new_n7601_ & new_n7860_;
  assign new_n7862_ = ~new_n7855_ & ~new_n7861_;
  assign new_n7863_ = ~\b[3]  & ~new_n7862_;
  assign new_n7864_ = ~new_n7443_ & ~\quotient[32] ;
  assign new_n7865_ = ~new_n7446_ & new_n7448_;
  assign new_n7866_ = ~new_n7444_ & new_n7865_;
  assign new_n7867_ = new_n432_ & ~new_n7866_;
  assign new_n7868_ = ~new_n7449_ & new_n7867_;
  assign new_n7869_ = ~new_n7601_ & new_n7868_;
  assign new_n7870_ = ~new_n7864_ & ~new_n7869_;
  assign new_n7871_ = ~\b[2]  & ~new_n7870_;
  assign new_n7872_ = \b[0]  & ~\b[32] ;
  assign new_n7873_ = new_n414_ & new_n7872_;
  assign new_n7874_ = new_n598_ & new_n7873_;
  assign new_n7875_ = new_n595_ & new_n7874_;
  assign new_n7876_ = ~new_n7601_ & new_n7875_;
  assign new_n7877_ = \a[32]  & ~new_n7876_;
  assign new_n7878_ = new_n313_ & new_n7448_;
  assign new_n7879_ = new_n303_ & new_n7878_;
  assign new_n7880_ = new_n288_ & new_n7879_;
  assign new_n7881_ = ~new_n7601_ & new_n7880_;
  assign new_n7882_ = ~new_n7877_ & ~new_n7881_;
  assign new_n7883_ = \b[1]  & ~new_n7882_;
  assign new_n7884_ = ~\b[1]  & ~new_n7881_;
  assign new_n7885_ = ~new_n7877_ & new_n7884_;
  assign new_n7886_ = ~new_n7883_ & ~new_n7885_;
  assign new_n7887_ = ~\a[31]  & \b[0] ;
  assign new_n7888_ = ~new_n7886_ & ~new_n7887_;
  assign new_n7889_ = ~\b[1]  & ~new_n7882_;
  assign new_n7890_ = ~new_n7888_ & ~new_n7889_;
  assign new_n7891_ = \b[2]  & ~new_n7869_;
  assign new_n7892_ = ~new_n7864_ & new_n7891_;
  assign new_n7893_ = ~new_n7871_ & ~new_n7892_;
  assign new_n7894_ = ~new_n7890_ & new_n7893_;
  assign new_n7895_ = ~new_n7871_ & ~new_n7894_;
  assign new_n7896_ = \b[3]  & ~new_n7861_;
  assign new_n7897_ = ~new_n7855_ & new_n7896_;
  assign new_n7898_ = ~new_n7863_ & ~new_n7897_;
  assign new_n7899_ = ~new_n7895_ & new_n7898_;
  assign new_n7900_ = ~new_n7863_ & ~new_n7899_;
  assign new_n7901_ = \b[4]  & ~new_n7852_;
  assign new_n7902_ = ~new_n7846_ & new_n7901_;
  assign new_n7903_ = ~new_n7854_ & ~new_n7902_;
  assign new_n7904_ = ~new_n7900_ & new_n7903_;
  assign new_n7905_ = ~new_n7854_ & ~new_n7904_;
  assign new_n7906_ = \b[5]  & ~new_n7843_;
  assign new_n7907_ = ~new_n7837_ & new_n7906_;
  assign new_n7908_ = ~new_n7845_ & ~new_n7907_;
  assign new_n7909_ = ~new_n7905_ & new_n7908_;
  assign new_n7910_ = ~new_n7845_ & ~new_n7909_;
  assign new_n7911_ = \b[6]  & ~new_n7834_;
  assign new_n7912_ = ~new_n7828_ & new_n7911_;
  assign new_n7913_ = ~new_n7836_ & ~new_n7912_;
  assign new_n7914_ = ~new_n7910_ & new_n7913_;
  assign new_n7915_ = ~new_n7836_ & ~new_n7914_;
  assign new_n7916_ = \b[7]  & ~new_n7825_;
  assign new_n7917_ = ~new_n7819_ & new_n7916_;
  assign new_n7918_ = ~new_n7827_ & ~new_n7917_;
  assign new_n7919_ = ~new_n7915_ & new_n7918_;
  assign new_n7920_ = ~new_n7827_ & ~new_n7919_;
  assign new_n7921_ = \b[8]  & ~new_n7816_;
  assign new_n7922_ = ~new_n7810_ & new_n7921_;
  assign new_n7923_ = ~new_n7818_ & ~new_n7922_;
  assign new_n7924_ = ~new_n7920_ & new_n7923_;
  assign new_n7925_ = ~new_n7818_ & ~new_n7924_;
  assign new_n7926_ = \b[9]  & ~new_n7807_;
  assign new_n7927_ = ~new_n7801_ & new_n7926_;
  assign new_n7928_ = ~new_n7809_ & ~new_n7927_;
  assign new_n7929_ = ~new_n7925_ & new_n7928_;
  assign new_n7930_ = ~new_n7809_ & ~new_n7929_;
  assign new_n7931_ = \b[10]  & ~new_n7798_;
  assign new_n7932_ = ~new_n7792_ & new_n7931_;
  assign new_n7933_ = ~new_n7800_ & ~new_n7932_;
  assign new_n7934_ = ~new_n7930_ & new_n7933_;
  assign new_n7935_ = ~new_n7800_ & ~new_n7934_;
  assign new_n7936_ = \b[11]  & ~new_n7789_;
  assign new_n7937_ = ~new_n7783_ & new_n7936_;
  assign new_n7938_ = ~new_n7791_ & ~new_n7937_;
  assign new_n7939_ = ~new_n7935_ & new_n7938_;
  assign new_n7940_ = ~new_n7791_ & ~new_n7939_;
  assign new_n7941_ = \b[12]  & ~new_n7780_;
  assign new_n7942_ = ~new_n7774_ & new_n7941_;
  assign new_n7943_ = ~new_n7782_ & ~new_n7942_;
  assign new_n7944_ = ~new_n7940_ & new_n7943_;
  assign new_n7945_ = ~new_n7782_ & ~new_n7944_;
  assign new_n7946_ = \b[13]  & ~new_n7771_;
  assign new_n7947_ = ~new_n7765_ & new_n7946_;
  assign new_n7948_ = ~new_n7773_ & ~new_n7947_;
  assign new_n7949_ = ~new_n7945_ & new_n7948_;
  assign new_n7950_ = ~new_n7773_ & ~new_n7949_;
  assign new_n7951_ = \b[14]  & ~new_n7762_;
  assign new_n7952_ = ~new_n7756_ & new_n7951_;
  assign new_n7953_ = ~new_n7764_ & ~new_n7952_;
  assign new_n7954_ = ~new_n7950_ & new_n7953_;
  assign new_n7955_ = ~new_n7764_ & ~new_n7954_;
  assign new_n7956_ = \b[15]  & ~new_n7753_;
  assign new_n7957_ = ~new_n7747_ & new_n7956_;
  assign new_n7958_ = ~new_n7755_ & ~new_n7957_;
  assign new_n7959_ = ~new_n7955_ & new_n7958_;
  assign new_n7960_ = ~new_n7755_ & ~new_n7959_;
  assign new_n7961_ = \b[16]  & ~new_n7744_;
  assign new_n7962_ = ~new_n7738_ & new_n7961_;
  assign new_n7963_ = ~new_n7746_ & ~new_n7962_;
  assign new_n7964_ = ~new_n7960_ & new_n7963_;
  assign new_n7965_ = ~new_n7746_ & ~new_n7964_;
  assign new_n7966_ = \b[17]  & ~new_n7735_;
  assign new_n7967_ = ~new_n7729_ & new_n7966_;
  assign new_n7968_ = ~new_n7737_ & ~new_n7967_;
  assign new_n7969_ = ~new_n7965_ & new_n7968_;
  assign new_n7970_ = ~new_n7737_ & ~new_n7969_;
  assign new_n7971_ = \b[18]  & ~new_n7726_;
  assign new_n7972_ = ~new_n7720_ & new_n7971_;
  assign new_n7973_ = ~new_n7728_ & ~new_n7972_;
  assign new_n7974_ = ~new_n7970_ & new_n7973_;
  assign new_n7975_ = ~new_n7728_ & ~new_n7974_;
  assign new_n7976_ = \b[19]  & ~new_n7717_;
  assign new_n7977_ = ~new_n7711_ & new_n7976_;
  assign new_n7978_ = ~new_n7719_ & ~new_n7977_;
  assign new_n7979_ = ~new_n7975_ & new_n7978_;
  assign new_n7980_ = ~new_n7719_ & ~new_n7979_;
  assign new_n7981_ = \b[20]  & ~new_n7708_;
  assign new_n7982_ = ~new_n7702_ & new_n7981_;
  assign new_n7983_ = ~new_n7710_ & ~new_n7982_;
  assign new_n7984_ = ~new_n7980_ & new_n7983_;
  assign new_n7985_ = ~new_n7710_ & ~new_n7984_;
  assign new_n7986_ = \b[21]  & ~new_n7699_;
  assign new_n7987_ = ~new_n7693_ & new_n7986_;
  assign new_n7988_ = ~new_n7701_ & ~new_n7987_;
  assign new_n7989_ = ~new_n7985_ & new_n7988_;
  assign new_n7990_ = ~new_n7701_ & ~new_n7989_;
  assign new_n7991_ = \b[22]  & ~new_n7690_;
  assign new_n7992_ = ~new_n7684_ & new_n7991_;
  assign new_n7993_ = ~new_n7692_ & ~new_n7992_;
  assign new_n7994_ = ~new_n7990_ & new_n7993_;
  assign new_n7995_ = ~new_n7692_ & ~new_n7994_;
  assign new_n7996_ = \b[23]  & ~new_n7681_;
  assign new_n7997_ = ~new_n7675_ & new_n7996_;
  assign new_n7998_ = ~new_n7683_ & ~new_n7997_;
  assign new_n7999_ = ~new_n7995_ & new_n7998_;
  assign new_n8000_ = ~new_n7683_ & ~new_n7999_;
  assign new_n8001_ = \b[24]  & ~new_n7672_;
  assign new_n8002_ = ~new_n7666_ & new_n8001_;
  assign new_n8003_ = ~new_n7674_ & ~new_n8002_;
  assign new_n8004_ = ~new_n8000_ & new_n8003_;
  assign new_n8005_ = ~new_n7674_ & ~new_n8004_;
  assign new_n8006_ = \b[25]  & ~new_n7663_;
  assign new_n8007_ = ~new_n7657_ & new_n8006_;
  assign new_n8008_ = ~new_n7665_ & ~new_n8007_;
  assign new_n8009_ = ~new_n8005_ & new_n8008_;
  assign new_n8010_ = ~new_n7665_ & ~new_n8009_;
  assign new_n8011_ = \b[26]  & ~new_n7654_;
  assign new_n8012_ = ~new_n7648_ & new_n8011_;
  assign new_n8013_ = ~new_n7656_ & ~new_n8012_;
  assign new_n8014_ = ~new_n8010_ & new_n8013_;
  assign new_n8015_ = ~new_n7656_ & ~new_n8014_;
  assign new_n8016_ = \b[27]  & ~new_n7645_;
  assign new_n8017_ = ~new_n7639_ & new_n8016_;
  assign new_n8018_ = ~new_n7647_ & ~new_n8017_;
  assign new_n8019_ = ~new_n8015_ & new_n8018_;
  assign new_n8020_ = ~new_n7647_ & ~new_n8019_;
  assign new_n8021_ = \b[28]  & ~new_n7636_;
  assign new_n8022_ = ~new_n7630_ & new_n8021_;
  assign new_n8023_ = ~new_n7638_ & ~new_n8022_;
  assign new_n8024_ = ~new_n8020_ & new_n8023_;
  assign new_n8025_ = ~new_n7638_ & ~new_n8024_;
  assign new_n8026_ = \b[29]  & ~new_n7627_;
  assign new_n8027_ = ~new_n7621_ & new_n8026_;
  assign new_n8028_ = ~new_n7629_ & ~new_n8027_;
  assign new_n8029_ = ~new_n8025_ & new_n8028_;
  assign new_n8030_ = ~new_n7629_ & ~new_n8029_;
  assign new_n8031_ = \b[30]  & ~new_n7618_;
  assign new_n8032_ = ~new_n7612_ & new_n8031_;
  assign new_n8033_ = ~new_n7620_ & ~new_n8032_;
  assign new_n8034_ = ~new_n8030_ & new_n8033_;
  assign new_n8035_ = ~new_n7620_ & ~new_n8034_;
  assign new_n8036_ = \b[31]  & ~new_n7609_;
  assign new_n8037_ = ~new_n7603_ & new_n8036_;
  assign new_n8038_ = ~new_n7611_ & ~new_n8037_;
  assign new_n8039_ = ~new_n8035_ & new_n8038_;
  assign new_n8040_ = ~new_n7611_ & ~new_n8039_;
  assign new_n8041_ = ~new_n7178_ & ~\quotient[32] ;
  assign new_n8042_ = ~new_n7180_ & new_n7599_;
  assign new_n8043_ = ~new_n7595_ & new_n8042_;
  assign new_n8044_ = ~new_n7596_ & ~new_n7599_;
  assign new_n8045_ = ~new_n8043_ & ~new_n8044_;
  assign new_n8046_ = \quotient[32]  & ~new_n8045_;
  assign new_n8047_ = ~new_n8041_ & ~new_n8046_;
  assign new_n8048_ = ~\b[32]  & ~new_n8047_;
  assign new_n8049_ = \b[32]  & ~new_n8041_;
  assign new_n8050_ = ~new_n8046_ & new_n8049_;
  assign new_n8051_ = new_n424_ & ~new_n8050_;
  assign new_n8052_ = ~new_n8048_ & new_n8051_;
  assign new_n8053_ = ~new_n8040_ & new_n8052_;
  assign new_n8054_ = new_n432_ & ~new_n8047_;
  assign \quotient[31]  = new_n8053_ | new_n8054_;
  assign new_n8056_ = ~new_n7620_ & new_n8038_;
  assign new_n8057_ = ~new_n8034_ & new_n8056_;
  assign new_n8058_ = ~new_n8035_ & ~new_n8038_;
  assign new_n8059_ = ~new_n8057_ & ~new_n8058_;
  assign new_n8060_ = \quotient[31]  & ~new_n8059_;
  assign new_n8061_ = ~new_n7610_ & ~new_n8054_;
  assign new_n8062_ = ~new_n8053_ & new_n8061_;
  assign new_n8063_ = ~new_n8060_ & ~new_n8062_;
  assign new_n8064_ = ~new_n7611_ & ~new_n8050_;
  assign new_n8065_ = ~new_n8048_ & new_n8064_;
  assign new_n8066_ = ~new_n8039_ & new_n8065_;
  assign new_n8067_ = ~new_n8048_ & ~new_n8050_;
  assign new_n8068_ = ~new_n8040_ & ~new_n8067_;
  assign new_n8069_ = ~new_n8066_ & ~new_n8068_;
  assign new_n8070_ = \quotient[31]  & ~new_n8069_;
  assign new_n8071_ = ~new_n8047_ & ~new_n8054_;
  assign new_n8072_ = ~new_n8053_ & new_n8071_;
  assign new_n8073_ = ~new_n8070_ & ~new_n8072_;
  assign new_n8074_ = ~\b[33]  & ~new_n8073_;
  assign new_n8075_ = ~\b[32]  & ~new_n8063_;
  assign new_n8076_ = ~new_n7629_ & new_n8033_;
  assign new_n8077_ = ~new_n8029_ & new_n8076_;
  assign new_n8078_ = ~new_n8030_ & ~new_n8033_;
  assign new_n8079_ = ~new_n8077_ & ~new_n8078_;
  assign new_n8080_ = \quotient[31]  & ~new_n8079_;
  assign new_n8081_ = ~new_n7619_ & ~new_n8054_;
  assign new_n8082_ = ~new_n8053_ & new_n8081_;
  assign new_n8083_ = ~new_n8080_ & ~new_n8082_;
  assign new_n8084_ = ~\b[31]  & ~new_n8083_;
  assign new_n8085_ = ~new_n7638_ & new_n8028_;
  assign new_n8086_ = ~new_n8024_ & new_n8085_;
  assign new_n8087_ = ~new_n8025_ & ~new_n8028_;
  assign new_n8088_ = ~new_n8086_ & ~new_n8087_;
  assign new_n8089_ = \quotient[31]  & ~new_n8088_;
  assign new_n8090_ = ~new_n7628_ & ~new_n8054_;
  assign new_n8091_ = ~new_n8053_ & new_n8090_;
  assign new_n8092_ = ~new_n8089_ & ~new_n8091_;
  assign new_n8093_ = ~\b[30]  & ~new_n8092_;
  assign new_n8094_ = ~new_n7647_ & new_n8023_;
  assign new_n8095_ = ~new_n8019_ & new_n8094_;
  assign new_n8096_ = ~new_n8020_ & ~new_n8023_;
  assign new_n8097_ = ~new_n8095_ & ~new_n8096_;
  assign new_n8098_ = \quotient[31]  & ~new_n8097_;
  assign new_n8099_ = ~new_n7637_ & ~new_n8054_;
  assign new_n8100_ = ~new_n8053_ & new_n8099_;
  assign new_n8101_ = ~new_n8098_ & ~new_n8100_;
  assign new_n8102_ = ~\b[29]  & ~new_n8101_;
  assign new_n8103_ = ~new_n7656_ & new_n8018_;
  assign new_n8104_ = ~new_n8014_ & new_n8103_;
  assign new_n8105_ = ~new_n8015_ & ~new_n8018_;
  assign new_n8106_ = ~new_n8104_ & ~new_n8105_;
  assign new_n8107_ = \quotient[31]  & ~new_n8106_;
  assign new_n8108_ = ~new_n7646_ & ~new_n8054_;
  assign new_n8109_ = ~new_n8053_ & new_n8108_;
  assign new_n8110_ = ~new_n8107_ & ~new_n8109_;
  assign new_n8111_ = ~\b[28]  & ~new_n8110_;
  assign new_n8112_ = ~new_n7665_ & new_n8013_;
  assign new_n8113_ = ~new_n8009_ & new_n8112_;
  assign new_n8114_ = ~new_n8010_ & ~new_n8013_;
  assign new_n8115_ = ~new_n8113_ & ~new_n8114_;
  assign new_n8116_ = \quotient[31]  & ~new_n8115_;
  assign new_n8117_ = ~new_n7655_ & ~new_n8054_;
  assign new_n8118_ = ~new_n8053_ & new_n8117_;
  assign new_n8119_ = ~new_n8116_ & ~new_n8118_;
  assign new_n8120_ = ~\b[27]  & ~new_n8119_;
  assign new_n8121_ = ~new_n7674_ & new_n8008_;
  assign new_n8122_ = ~new_n8004_ & new_n8121_;
  assign new_n8123_ = ~new_n8005_ & ~new_n8008_;
  assign new_n8124_ = ~new_n8122_ & ~new_n8123_;
  assign new_n8125_ = \quotient[31]  & ~new_n8124_;
  assign new_n8126_ = ~new_n7664_ & ~new_n8054_;
  assign new_n8127_ = ~new_n8053_ & new_n8126_;
  assign new_n8128_ = ~new_n8125_ & ~new_n8127_;
  assign new_n8129_ = ~\b[26]  & ~new_n8128_;
  assign new_n8130_ = ~new_n7683_ & new_n8003_;
  assign new_n8131_ = ~new_n7999_ & new_n8130_;
  assign new_n8132_ = ~new_n8000_ & ~new_n8003_;
  assign new_n8133_ = ~new_n8131_ & ~new_n8132_;
  assign new_n8134_ = \quotient[31]  & ~new_n8133_;
  assign new_n8135_ = ~new_n7673_ & ~new_n8054_;
  assign new_n8136_ = ~new_n8053_ & new_n8135_;
  assign new_n8137_ = ~new_n8134_ & ~new_n8136_;
  assign new_n8138_ = ~\b[25]  & ~new_n8137_;
  assign new_n8139_ = ~new_n7692_ & new_n7998_;
  assign new_n8140_ = ~new_n7994_ & new_n8139_;
  assign new_n8141_ = ~new_n7995_ & ~new_n7998_;
  assign new_n8142_ = ~new_n8140_ & ~new_n8141_;
  assign new_n8143_ = \quotient[31]  & ~new_n8142_;
  assign new_n8144_ = ~new_n7682_ & ~new_n8054_;
  assign new_n8145_ = ~new_n8053_ & new_n8144_;
  assign new_n8146_ = ~new_n8143_ & ~new_n8145_;
  assign new_n8147_ = ~\b[24]  & ~new_n8146_;
  assign new_n8148_ = ~new_n7701_ & new_n7993_;
  assign new_n8149_ = ~new_n7989_ & new_n8148_;
  assign new_n8150_ = ~new_n7990_ & ~new_n7993_;
  assign new_n8151_ = ~new_n8149_ & ~new_n8150_;
  assign new_n8152_ = \quotient[31]  & ~new_n8151_;
  assign new_n8153_ = ~new_n7691_ & ~new_n8054_;
  assign new_n8154_ = ~new_n8053_ & new_n8153_;
  assign new_n8155_ = ~new_n8152_ & ~new_n8154_;
  assign new_n8156_ = ~\b[23]  & ~new_n8155_;
  assign new_n8157_ = ~new_n7710_ & new_n7988_;
  assign new_n8158_ = ~new_n7984_ & new_n8157_;
  assign new_n8159_ = ~new_n7985_ & ~new_n7988_;
  assign new_n8160_ = ~new_n8158_ & ~new_n8159_;
  assign new_n8161_ = \quotient[31]  & ~new_n8160_;
  assign new_n8162_ = ~new_n7700_ & ~new_n8054_;
  assign new_n8163_ = ~new_n8053_ & new_n8162_;
  assign new_n8164_ = ~new_n8161_ & ~new_n8163_;
  assign new_n8165_ = ~\b[22]  & ~new_n8164_;
  assign new_n8166_ = ~new_n7719_ & new_n7983_;
  assign new_n8167_ = ~new_n7979_ & new_n8166_;
  assign new_n8168_ = ~new_n7980_ & ~new_n7983_;
  assign new_n8169_ = ~new_n8167_ & ~new_n8168_;
  assign new_n8170_ = \quotient[31]  & ~new_n8169_;
  assign new_n8171_ = ~new_n7709_ & ~new_n8054_;
  assign new_n8172_ = ~new_n8053_ & new_n8171_;
  assign new_n8173_ = ~new_n8170_ & ~new_n8172_;
  assign new_n8174_ = ~\b[21]  & ~new_n8173_;
  assign new_n8175_ = ~new_n7728_ & new_n7978_;
  assign new_n8176_ = ~new_n7974_ & new_n8175_;
  assign new_n8177_ = ~new_n7975_ & ~new_n7978_;
  assign new_n8178_ = ~new_n8176_ & ~new_n8177_;
  assign new_n8179_ = \quotient[31]  & ~new_n8178_;
  assign new_n8180_ = ~new_n7718_ & ~new_n8054_;
  assign new_n8181_ = ~new_n8053_ & new_n8180_;
  assign new_n8182_ = ~new_n8179_ & ~new_n8181_;
  assign new_n8183_ = ~\b[20]  & ~new_n8182_;
  assign new_n8184_ = ~new_n7737_ & new_n7973_;
  assign new_n8185_ = ~new_n7969_ & new_n8184_;
  assign new_n8186_ = ~new_n7970_ & ~new_n7973_;
  assign new_n8187_ = ~new_n8185_ & ~new_n8186_;
  assign new_n8188_ = \quotient[31]  & ~new_n8187_;
  assign new_n8189_ = ~new_n7727_ & ~new_n8054_;
  assign new_n8190_ = ~new_n8053_ & new_n8189_;
  assign new_n8191_ = ~new_n8188_ & ~new_n8190_;
  assign new_n8192_ = ~\b[19]  & ~new_n8191_;
  assign new_n8193_ = ~new_n7746_ & new_n7968_;
  assign new_n8194_ = ~new_n7964_ & new_n8193_;
  assign new_n8195_ = ~new_n7965_ & ~new_n7968_;
  assign new_n8196_ = ~new_n8194_ & ~new_n8195_;
  assign new_n8197_ = \quotient[31]  & ~new_n8196_;
  assign new_n8198_ = ~new_n7736_ & ~new_n8054_;
  assign new_n8199_ = ~new_n8053_ & new_n8198_;
  assign new_n8200_ = ~new_n8197_ & ~new_n8199_;
  assign new_n8201_ = ~\b[18]  & ~new_n8200_;
  assign new_n8202_ = ~new_n7755_ & new_n7963_;
  assign new_n8203_ = ~new_n7959_ & new_n8202_;
  assign new_n8204_ = ~new_n7960_ & ~new_n7963_;
  assign new_n8205_ = ~new_n8203_ & ~new_n8204_;
  assign new_n8206_ = \quotient[31]  & ~new_n8205_;
  assign new_n8207_ = ~new_n7745_ & ~new_n8054_;
  assign new_n8208_ = ~new_n8053_ & new_n8207_;
  assign new_n8209_ = ~new_n8206_ & ~new_n8208_;
  assign new_n8210_ = ~\b[17]  & ~new_n8209_;
  assign new_n8211_ = ~new_n7764_ & new_n7958_;
  assign new_n8212_ = ~new_n7954_ & new_n8211_;
  assign new_n8213_ = ~new_n7955_ & ~new_n7958_;
  assign new_n8214_ = ~new_n8212_ & ~new_n8213_;
  assign new_n8215_ = \quotient[31]  & ~new_n8214_;
  assign new_n8216_ = ~new_n7754_ & ~new_n8054_;
  assign new_n8217_ = ~new_n8053_ & new_n8216_;
  assign new_n8218_ = ~new_n8215_ & ~new_n8217_;
  assign new_n8219_ = ~\b[16]  & ~new_n8218_;
  assign new_n8220_ = ~new_n7773_ & new_n7953_;
  assign new_n8221_ = ~new_n7949_ & new_n8220_;
  assign new_n8222_ = ~new_n7950_ & ~new_n7953_;
  assign new_n8223_ = ~new_n8221_ & ~new_n8222_;
  assign new_n8224_ = \quotient[31]  & ~new_n8223_;
  assign new_n8225_ = ~new_n7763_ & ~new_n8054_;
  assign new_n8226_ = ~new_n8053_ & new_n8225_;
  assign new_n8227_ = ~new_n8224_ & ~new_n8226_;
  assign new_n8228_ = ~\b[15]  & ~new_n8227_;
  assign new_n8229_ = ~new_n7782_ & new_n7948_;
  assign new_n8230_ = ~new_n7944_ & new_n8229_;
  assign new_n8231_ = ~new_n7945_ & ~new_n7948_;
  assign new_n8232_ = ~new_n8230_ & ~new_n8231_;
  assign new_n8233_ = \quotient[31]  & ~new_n8232_;
  assign new_n8234_ = ~new_n7772_ & ~new_n8054_;
  assign new_n8235_ = ~new_n8053_ & new_n8234_;
  assign new_n8236_ = ~new_n8233_ & ~new_n8235_;
  assign new_n8237_ = ~\b[14]  & ~new_n8236_;
  assign new_n8238_ = ~new_n7791_ & new_n7943_;
  assign new_n8239_ = ~new_n7939_ & new_n8238_;
  assign new_n8240_ = ~new_n7940_ & ~new_n7943_;
  assign new_n8241_ = ~new_n8239_ & ~new_n8240_;
  assign new_n8242_ = \quotient[31]  & ~new_n8241_;
  assign new_n8243_ = ~new_n7781_ & ~new_n8054_;
  assign new_n8244_ = ~new_n8053_ & new_n8243_;
  assign new_n8245_ = ~new_n8242_ & ~new_n8244_;
  assign new_n8246_ = ~\b[13]  & ~new_n8245_;
  assign new_n8247_ = ~new_n7800_ & new_n7938_;
  assign new_n8248_ = ~new_n7934_ & new_n8247_;
  assign new_n8249_ = ~new_n7935_ & ~new_n7938_;
  assign new_n8250_ = ~new_n8248_ & ~new_n8249_;
  assign new_n8251_ = \quotient[31]  & ~new_n8250_;
  assign new_n8252_ = ~new_n7790_ & ~new_n8054_;
  assign new_n8253_ = ~new_n8053_ & new_n8252_;
  assign new_n8254_ = ~new_n8251_ & ~new_n8253_;
  assign new_n8255_ = ~\b[12]  & ~new_n8254_;
  assign new_n8256_ = ~new_n7809_ & new_n7933_;
  assign new_n8257_ = ~new_n7929_ & new_n8256_;
  assign new_n8258_ = ~new_n7930_ & ~new_n7933_;
  assign new_n8259_ = ~new_n8257_ & ~new_n8258_;
  assign new_n8260_ = \quotient[31]  & ~new_n8259_;
  assign new_n8261_ = ~new_n7799_ & ~new_n8054_;
  assign new_n8262_ = ~new_n8053_ & new_n8261_;
  assign new_n8263_ = ~new_n8260_ & ~new_n8262_;
  assign new_n8264_ = ~\b[11]  & ~new_n8263_;
  assign new_n8265_ = ~new_n7818_ & new_n7928_;
  assign new_n8266_ = ~new_n7924_ & new_n8265_;
  assign new_n8267_ = ~new_n7925_ & ~new_n7928_;
  assign new_n8268_ = ~new_n8266_ & ~new_n8267_;
  assign new_n8269_ = \quotient[31]  & ~new_n8268_;
  assign new_n8270_ = ~new_n7808_ & ~new_n8054_;
  assign new_n8271_ = ~new_n8053_ & new_n8270_;
  assign new_n8272_ = ~new_n8269_ & ~new_n8271_;
  assign new_n8273_ = ~\b[10]  & ~new_n8272_;
  assign new_n8274_ = ~new_n7827_ & new_n7923_;
  assign new_n8275_ = ~new_n7919_ & new_n8274_;
  assign new_n8276_ = ~new_n7920_ & ~new_n7923_;
  assign new_n8277_ = ~new_n8275_ & ~new_n8276_;
  assign new_n8278_ = \quotient[31]  & ~new_n8277_;
  assign new_n8279_ = ~new_n7817_ & ~new_n8054_;
  assign new_n8280_ = ~new_n8053_ & new_n8279_;
  assign new_n8281_ = ~new_n8278_ & ~new_n8280_;
  assign new_n8282_ = ~\b[9]  & ~new_n8281_;
  assign new_n8283_ = ~new_n7836_ & new_n7918_;
  assign new_n8284_ = ~new_n7914_ & new_n8283_;
  assign new_n8285_ = ~new_n7915_ & ~new_n7918_;
  assign new_n8286_ = ~new_n8284_ & ~new_n8285_;
  assign new_n8287_ = \quotient[31]  & ~new_n8286_;
  assign new_n8288_ = ~new_n7826_ & ~new_n8054_;
  assign new_n8289_ = ~new_n8053_ & new_n8288_;
  assign new_n8290_ = ~new_n8287_ & ~new_n8289_;
  assign new_n8291_ = ~\b[8]  & ~new_n8290_;
  assign new_n8292_ = ~new_n7845_ & new_n7913_;
  assign new_n8293_ = ~new_n7909_ & new_n8292_;
  assign new_n8294_ = ~new_n7910_ & ~new_n7913_;
  assign new_n8295_ = ~new_n8293_ & ~new_n8294_;
  assign new_n8296_ = \quotient[31]  & ~new_n8295_;
  assign new_n8297_ = ~new_n7835_ & ~new_n8054_;
  assign new_n8298_ = ~new_n8053_ & new_n8297_;
  assign new_n8299_ = ~new_n8296_ & ~new_n8298_;
  assign new_n8300_ = ~\b[7]  & ~new_n8299_;
  assign new_n8301_ = ~new_n7854_ & new_n7908_;
  assign new_n8302_ = ~new_n7904_ & new_n8301_;
  assign new_n8303_ = ~new_n7905_ & ~new_n7908_;
  assign new_n8304_ = ~new_n8302_ & ~new_n8303_;
  assign new_n8305_ = \quotient[31]  & ~new_n8304_;
  assign new_n8306_ = ~new_n7844_ & ~new_n8054_;
  assign new_n8307_ = ~new_n8053_ & new_n8306_;
  assign new_n8308_ = ~new_n8305_ & ~new_n8307_;
  assign new_n8309_ = ~\b[6]  & ~new_n8308_;
  assign new_n8310_ = ~new_n7863_ & new_n7903_;
  assign new_n8311_ = ~new_n7899_ & new_n8310_;
  assign new_n8312_ = ~new_n7900_ & ~new_n7903_;
  assign new_n8313_ = ~new_n8311_ & ~new_n8312_;
  assign new_n8314_ = \quotient[31]  & ~new_n8313_;
  assign new_n8315_ = ~new_n7853_ & ~new_n8054_;
  assign new_n8316_ = ~new_n8053_ & new_n8315_;
  assign new_n8317_ = ~new_n8314_ & ~new_n8316_;
  assign new_n8318_ = ~\b[5]  & ~new_n8317_;
  assign new_n8319_ = ~new_n7871_ & new_n7898_;
  assign new_n8320_ = ~new_n7894_ & new_n8319_;
  assign new_n8321_ = ~new_n7895_ & ~new_n7898_;
  assign new_n8322_ = ~new_n8320_ & ~new_n8321_;
  assign new_n8323_ = \quotient[31]  & ~new_n8322_;
  assign new_n8324_ = ~new_n7862_ & ~new_n8054_;
  assign new_n8325_ = ~new_n8053_ & new_n8324_;
  assign new_n8326_ = ~new_n8323_ & ~new_n8325_;
  assign new_n8327_ = ~\b[4]  & ~new_n8326_;
  assign new_n8328_ = ~new_n7889_ & new_n7893_;
  assign new_n8329_ = ~new_n7888_ & new_n8328_;
  assign new_n8330_ = ~new_n7890_ & ~new_n7893_;
  assign new_n8331_ = ~new_n8329_ & ~new_n8330_;
  assign new_n8332_ = \quotient[31]  & ~new_n8331_;
  assign new_n8333_ = ~new_n7870_ & ~new_n8054_;
  assign new_n8334_ = ~new_n8053_ & new_n8333_;
  assign new_n8335_ = ~new_n8332_ & ~new_n8334_;
  assign new_n8336_ = ~\b[3]  & ~new_n8335_;
  assign new_n8337_ = ~new_n7885_ & new_n7887_;
  assign new_n8338_ = ~new_n7883_ & new_n8337_;
  assign new_n8339_ = ~new_n7888_ & ~new_n8338_;
  assign new_n8340_ = \quotient[31]  & new_n8339_;
  assign new_n8341_ = ~new_n7882_ & ~new_n8054_;
  assign new_n8342_ = ~new_n8053_ & new_n8341_;
  assign new_n8343_ = ~new_n8340_ & ~new_n8342_;
  assign new_n8344_ = ~\b[2]  & ~new_n8343_;
  assign new_n8345_ = \b[0]  & \quotient[31] ;
  assign new_n8346_ = \a[31]  & ~new_n8345_;
  assign new_n8347_ = new_n7887_ & \quotient[31] ;
  assign new_n8348_ = ~new_n8346_ & ~new_n8347_;
  assign new_n8349_ = \b[1]  & ~new_n8348_;
  assign new_n8350_ = ~\b[1]  & ~new_n8347_;
  assign new_n8351_ = ~new_n8346_ & new_n8350_;
  assign new_n8352_ = ~new_n8349_ & ~new_n8351_;
  assign new_n8353_ = ~\a[30]  & \b[0] ;
  assign new_n8354_ = ~new_n8352_ & ~new_n8353_;
  assign new_n8355_ = ~\b[1]  & ~new_n8348_;
  assign new_n8356_ = ~new_n8354_ & ~new_n8355_;
  assign new_n8357_ = \b[2]  & ~new_n8342_;
  assign new_n8358_ = ~new_n8340_ & new_n8357_;
  assign new_n8359_ = ~new_n8344_ & ~new_n8358_;
  assign new_n8360_ = ~new_n8356_ & new_n8359_;
  assign new_n8361_ = ~new_n8344_ & ~new_n8360_;
  assign new_n8362_ = \b[3]  & ~new_n8334_;
  assign new_n8363_ = ~new_n8332_ & new_n8362_;
  assign new_n8364_ = ~new_n8336_ & ~new_n8363_;
  assign new_n8365_ = ~new_n8361_ & new_n8364_;
  assign new_n8366_ = ~new_n8336_ & ~new_n8365_;
  assign new_n8367_ = \b[4]  & ~new_n8325_;
  assign new_n8368_ = ~new_n8323_ & new_n8367_;
  assign new_n8369_ = ~new_n8327_ & ~new_n8368_;
  assign new_n8370_ = ~new_n8366_ & new_n8369_;
  assign new_n8371_ = ~new_n8327_ & ~new_n8370_;
  assign new_n8372_ = \b[5]  & ~new_n8316_;
  assign new_n8373_ = ~new_n8314_ & new_n8372_;
  assign new_n8374_ = ~new_n8318_ & ~new_n8373_;
  assign new_n8375_ = ~new_n8371_ & new_n8374_;
  assign new_n8376_ = ~new_n8318_ & ~new_n8375_;
  assign new_n8377_ = \b[6]  & ~new_n8307_;
  assign new_n8378_ = ~new_n8305_ & new_n8377_;
  assign new_n8379_ = ~new_n8309_ & ~new_n8378_;
  assign new_n8380_ = ~new_n8376_ & new_n8379_;
  assign new_n8381_ = ~new_n8309_ & ~new_n8380_;
  assign new_n8382_ = \b[7]  & ~new_n8298_;
  assign new_n8383_ = ~new_n8296_ & new_n8382_;
  assign new_n8384_ = ~new_n8300_ & ~new_n8383_;
  assign new_n8385_ = ~new_n8381_ & new_n8384_;
  assign new_n8386_ = ~new_n8300_ & ~new_n8385_;
  assign new_n8387_ = \b[8]  & ~new_n8289_;
  assign new_n8388_ = ~new_n8287_ & new_n8387_;
  assign new_n8389_ = ~new_n8291_ & ~new_n8388_;
  assign new_n8390_ = ~new_n8386_ & new_n8389_;
  assign new_n8391_ = ~new_n8291_ & ~new_n8390_;
  assign new_n8392_ = \b[9]  & ~new_n8280_;
  assign new_n8393_ = ~new_n8278_ & new_n8392_;
  assign new_n8394_ = ~new_n8282_ & ~new_n8393_;
  assign new_n8395_ = ~new_n8391_ & new_n8394_;
  assign new_n8396_ = ~new_n8282_ & ~new_n8395_;
  assign new_n8397_ = \b[10]  & ~new_n8271_;
  assign new_n8398_ = ~new_n8269_ & new_n8397_;
  assign new_n8399_ = ~new_n8273_ & ~new_n8398_;
  assign new_n8400_ = ~new_n8396_ & new_n8399_;
  assign new_n8401_ = ~new_n8273_ & ~new_n8400_;
  assign new_n8402_ = \b[11]  & ~new_n8262_;
  assign new_n8403_ = ~new_n8260_ & new_n8402_;
  assign new_n8404_ = ~new_n8264_ & ~new_n8403_;
  assign new_n8405_ = ~new_n8401_ & new_n8404_;
  assign new_n8406_ = ~new_n8264_ & ~new_n8405_;
  assign new_n8407_ = \b[12]  & ~new_n8253_;
  assign new_n8408_ = ~new_n8251_ & new_n8407_;
  assign new_n8409_ = ~new_n8255_ & ~new_n8408_;
  assign new_n8410_ = ~new_n8406_ & new_n8409_;
  assign new_n8411_ = ~new_n8255_ & ~new_n8410_;
  assign new_n8412_ = \b[13]  & ~new_n8244_;
  assign new_n8413_ = ~new_n8242_ & new_n8412_;
  assign new_n8414_ = ~new_n8246_ & ~new_n8413_;
  assign new_n8415_ = ~new_n8411_ & new_n8414_;
  assign new_n8416_ = ~new_n8246_ & ~new_n8415_;
  assign new_n8417_ = \b[14]  & ~new_n8235_;
  assign new_n8418_ = ~new_n8233_ & new_n8417_;
  assign new_n8419_ = ~new_n8237_ & ~new_n8418_;
  assign new_n8420_ = ~new_n8416_ & new_n8419_;
  assign new_n8421_ = ~new_n8237_ & ~new_n8420_;
  assign new_n8422_ = \b[15]  & ~new_n8226_;
  assign new_n8423_ = ~new_n8224_ & new_n8422_;
  assign new_n8424_ = ~new_n8228_ & ~new_n8423_;
  assign new_n8425_ = ~new_n8421_ & new_n8424_;
  assign new_n8426_ = ~new_n8228_ & ~new_n8425_;
  assign new_n8427_ = \b[16]  & ~new_n8217_;
  assign new_n8428_ = ~new_n8215_ & new_n8427_;
  assign new_n8429_ = ~new_n8219_ & ~new_n8428_;
  assign new_n8430_ = ~new_n8426_ & new_n8429_;
  assign new_n8431_ = ~new_n8219_ & ~new_n8430_;
  assign new_n8432_ = \b[17]  & ~new_n8208_;
  assign new_n8433_ = ~new_n8206_ & new_n8432_;
  assign new_n8434_ = ~new_n8210_ & ~new_n8433_;
  assign new_n8435_ = ~new_n8431_ & new_n8434_;
  assign new_n8436_ = ~new_n8210_ & ~new_n8435_;
  assign new_n8437_ = \b[18]  & ~new_n8199_;
  assign new_n8438_ = ~new_n8197_ & new_n8437_;
  assign new_n8439_ = ~new_n8201_ & ~new_n8438_;
  assign new_n8440_ = ~new_n8436_ & new_n8439_;
  assign new_n8441_ = ~new_n8201_ & ~new_n8440_;
  assign new_n8442_ = \b[19]  & ~new_n8190_;
  assign new_n8443_ = ~new_n8188_ & new_n8442_;
  assign new_n8444_ = ~new_n8192_ & ~new_n8443_;
  assign new_n8445_ = ~new_n8441_ & new_n8444_;
  assign new_n8446_ = ~new_n8192_ & ~new_n8445_;
  assign new_n8447_ = \b[20]  & ~new_n8181_;
  assign new_n8448_ = ~new_n8179_ & new_n8447_;
  assign new_n8449_ = ~new_n8183_ & ~new_n8448_;
  assign new_n8450_ = ~new_n8446_ & new_n8449_;
  assign new_n8451_ = ~new_n8183_ & ~new_n8450_;
  assign new_n8452_ = \b[21]  & ~new_n8172_;
  assign new_n8453_ = ~new_n8170_ & new_n8452_;
  assign new_n8454_ = ~new_n8174_ & ~new_n8453_;
  assign new_n8455_ = ~new_n8451_ & new_n8454_;
  assign new_n8456_ = ~new_n8174_ & ~new_n8455_;
  assign new_n8457_ = \b[22]  & ~new_n8163_;
  assign new_n8458_ = ~new_n8161_ & new_n8457_;
  assign new_n8459_ = ~new_n8165_ & ~new_n8458_;
  assign new_n8460_ = ~new_n8456_ & new_n8459_;
  assign new_n8461_ = ~new_n8165_ & ~new_n8460_;
  assign new_n8462_ = \b[23]  & ~new_n8154_;
  assign new_n8463_ = ~new_n8152_ & new_n8462_;
  assign new_n8464_ = ~new_n8156_ & ~new_n8463_;
  assign new_n8465_ = ~new_n8461_ & new_n8464_;
  assign new_n8466_ = ~new_n8156_ & ~new_n8465_;
  assign new_n8467_ = \b[24]  & ~new_n8145_;
  assign new_n8468_ = ~new_n8143_ & new_n8467_;
  assign new_n8469_ = ~new_n8147_ & ~new_n8468_;
  assign new_n8470_ = ~new_n8466_ & new_n8469_;
  assign new_n8471_ = ~new_n8147_ & ~new_n8470_;
  assign new_n8472_ = \b[25]  & ~new_n8136_;
  assign new_n8473_ = ~new_n8134_ & new_n8472_;
  assign new_n8474_ = ~new_n8138_ & ~new_n8473_;
  assign new_n8475_ = ~new_n8471_ & new_n8474_;
  assign new_n8476_ = ~new_n8138_ & ~new_n8475_;
  assign new_n8477_ = \b[26]  & ~new_n8127_;
  assign new_n8478_ = ~new_n8125_ & new_n8477_;
  assign new_n8479_ = ~new_n8129_ & ~new_n8478_;
  assign new_n8480_ = ~new_n8476_ & new_n8479_;
  assign new_n8481_ = ~new_n8129_ & ~new_n8480_;
  assign new_n8482_ = \b[27]  & ~new_n8118_;
  assign new_n8483_ = ~new_n8116_ & new_n8482_;
  assign new_n8484_ = ~new_n8120_ & ~new_n8483_;
  assign new_n8485_ = ~new_n8481_ & new_n8484_;
  assign new_n8486_ = ~new_n8120_ & ~new_n8485_;
  assign new_n8487_ = \b[28]  & ~new_n8109_;
  assign new_n8488_ = ~new_n8107_ & new_n8487_;
  assign new_n8489_ = ~new_n8111_ & ~new_n8488_;
  assign new_n8490_ = ~new_n8486_ & new_n8489_;
  assign new_n8491_ = ~new_n8111_ & ~new_n8490_;
  assign new_n8492_ = \b[29]  & ~new_n8100_;
  assign new_n8493_ = ~new_n8098_ & new_n8492_;
  assign new_n8494_ = ~new_n8102_ & ~new_n8493_;
  assign new_n8495_ = ~new_n8491_ & new_n8494_;
  assign new_n8496_ = ~new_n8102_ & ~new_n8495_;
  assign new_n8497_ = \b[30]  & ~new_n8091_;
  assign new_n8498_ = ~new_n8089_ & new_n8497_;
  assign new_n8499_ = ~new_n8093_ & ~new_n8498_;
  assign new_n8500_ = ~new_n8496_ & new_n8499_;
  assign new_n8501_ = ~new_n8093_ & ~new_n8500_;
  assign new_n8502_ = \b[31]  & ~new_n8082_;
  assign new_n8503_ = ~new_n8080_ & new_n8502_;
  assign new_n8504_ = ~new_n8084_ & ~new_n8503_;
  assign new_n8505_ = ~new_n8501_ & new_n8504_;
  assign new_n8506_ = ~new_n8084_ & ~new_n8505_;
  assign new_n8507_ = \b[32]  & ~new_n8062_;
  assign new_n8508_ = ~new_n8060_ & new_n8507_;
  assign new_n8509_ = ~new_n8075_ & ~new_n8508_;
  assign new_n8510_ = ~new_n8506_ & new_n8509_;
  assign new_n8511_ = ~new_n8075_ & ~new_n8510_;
  assign new_n8512_ = \b[33]  & ~new_n8072_;
  assign new_n8513_ = ~new_n8070_ & new_n8512_;
  assign new_n8514_ = ~new_n8074_ & ~new_n8513_;
  assign new_n8515_ = ~new_n8511_ & new_n8514_;
  assign new_n8516_ = ~new_n8074_ & ~new_n8515_;
  assign new_n8517_ = new_n294_ & new_n312_;
  assign new_n8518_ = new_n340_ & new_n8517_;
  assign new_n8519_ = new_n338_ & new_n8518_;
  assign \quotient[30]  = ~new_n8516_ & new_n8519_;
  assign new_n8521_ = ~new_n8063_ & ~\quotient[30] ;
  assign new_n8522_ = ~new_n8084_ & new_n8509_;
  assign new_n8523_ = ~new_n8505_ & new_n8522_;
  assign new_n8524_ = ~new_n8506_ & ~new_n8509_;
  assign new_n8525_ = ~new_n8523_ & ~new_n8524_;
  assign new_n8526_ = new_n8519_ & ~new_n8525_;
  assign new_n8527_ = ~new_n8516_ & new_n8526_;
  assign new_n8528_ = ~new_n8521_ & ~new_n8527_;
  assign new_n8529_ = ~new_n8073_ & ~\quotient[30] ;
  assign new_n8530_ = ~new_n8075_ & new_n8514_;
  assign new_n8531_ = ~new_n8510_ & new_n8530_;
  assign new_n8532_ = ~new_n8511_ & ~new_n8514_;
  assign new_n8533_ = ~new_n8531_ & ~new_n8532_;
  assign new_n8534_ = \quotient[30]  & ~new_n8533_;
  assign new_n8535_ = ~new_n8529_ & ~new_n8534_;
  assign new_n8536_ = ~\b[34]  & ~new_n8535_;
  assign new_n8537_ = ~\b[33]  & ~new_n8528_;
  assign new_n8538_ = ~new_n8083_ & ~\quotient[30] ;
  assign new_n8539_ = ~new_n8093_ & new_n8504_;
  assign new_n8540_ = ~new_n8500_ & new_n8539_;
  assign new_n8541_ = ~new_n8501_ & ~new_n8504_;
  assign new_n8542_ = ~new_n8540_ & ~new_n8541_;
  assign new_n8543_ = new_n8519_ & ~new_n8542_;
  assign new_n8544_ = ~new_n8516_ & new_n8543_;
  assign new_n8545_ = ~new_n8538_ & ~new_n8544_;
  assign new_n8546_ = ~\b[32]  & ~new_n8545_;
  assign new_n8547_ = ~new_n8092_ & ~\quotient[30] ;
  assign new_n8548_ = ~new_n8102_ & new_n8499_;
  assign new_n8549_ = ~new_n8495_ & new_n8548_;
  assign new_n8550_ = ~new_n8496_ & ~new_n8499_;
  assign new_n8551_ = ~new_n8549_ & ~new_n8550_;
  assign new_n8552_ = new_n8519_ & ~new_n8551_;
  assign new_n8553_ = ~new_n8516_ & new_n8552_;
  assign new_n8554_ = ~new_n8547_ & ~new_n8553_;
  assign new_n8555_ = ~\b[31]  & ~new_n8554_;
  assign new_n8556_ = ~new_n8101_ & ~\quotient[30] ;
  assign new_n8557_ = ~new_n8111_ & new_n8494_;
  assign new_n8558_ = ~new_n8490_ & new_n8557_;
  assign new_n8559_ = ~new_n8491_ & ~new_n8494_;
  assign new_n8560_ = ~new_n8558_ & ~new_n8559_;
  assign new_n8561_ = new_n8519_ & ~new_n8560_;
  assign new_n8562_ = ~new_n8516_ & new_n8561_;
  assign new_n8563_ = ~new_n8556_ & ~new_n8562_;
  assign new_n8564_ = ~\b[30]  & ~new_n8563_;
  assign new_n8565_ = ~new_n8110_ & ~\quotient[30] ;
  assign new_n8566_ = ~new_n8120_ & new_n8489_;
  assign new_n8567_ = ~new_n8485_ & new_n8566_;
  assign new_n8568_ = ~new_n8486_ & ~new_n8489_;
  assign new_n8569_ = ~new_n8567_ & ~new_n8568_;
  assign new_n8570_ = new_n8519_ & ~new_n8569_;
  assign new_n8571_ = ~new_n8516_ & new_n8570_;
  assign new_n8572_ = ~new_n8565_ & ~new_n8571_;
  assign new_n8573_ = ~\b[29]  & ~new_n8572_;
  assign new_n8574_ = ~new_n8119_ & ~\quotient[30] ;
  assign new_n8575_ = ~new_n8129_ & new_n8484_;
  assign new_n8576_ = ~new_n8480_ & new_n8575_;
  assign new_n8577_ = ~new_n8481_ & ~new_n8484_;
  assign new_n8578_ = ~new_n8576_ & ~new_n8577_;
  assign new_n8579_ = new_n8519_ & ~new_n8578_;
  assign new_n8580_ = ~new_n8516_ & new_n8579_;
  assign new_n8581_ = ~new_n8574_ & ~new_n8580_;
  assign new_n8582_ = ~\b[28]  & ~new_n8581_;
  assign new_n8583_ = ~new_n8128_ & ~\quotient[30] ;
  assign new_n8584_ = ~new_n8138_ & new_n8479_;
  assign new_n8585_ = ~new_n8475_ & new_n8584_;
  assign new_n8586_ = ~new_n8476_ & ~new_n8479_;
  assign new_n8587_ = ~new_n8585_ & ~new_n8586_;
  assign new_n8588_ = new_n8519_ & ~new_n8587_;
  assign new_n8589_ = ~new_n8516_ & new_n8588_;
  assign new_n8590_ = ~new_n8583_ & ~new_n8589_;
  assign new_n8591_ = ~\b[27]  & ~new_n8590_;
  assign new_n8592_ = ~new_n8137_ & ~\quotient[30] ;
  assign new_n8593_ = ~new_n8147_ & new_n8474_;
  assign new_n8594_ = ~new_n8470_ & new_n8593_;
  assign new_n8595_ = ~new_n8471_ & ~new_n8474_;
  assign new_n8596_ = ~new_n8594_ & ~new_n8595_;
  assign new_n8597_ = new_n8519_ & ~new_n8596_;
  assign new_n8598_ = ~new_n8516_ & new_n8597_;
  assign new_n8599_ = ~new_n8592_ & ~new_n8598_;
  assign new_n8600_ = ~\b[26]  & ~new_n8599_;
  assign new_n8601_ = ~new_n8146_ & ~\quotient[30] ;
  assign new_n8602_ = ~new_n8156_ & new_n8469_;
  assign new_n8603_ = ~new_n8465_ & new_n8602_;
  assign new_n8604_ = ~new_n8466_ & ~new_n8469_;
  assign new_n8605_ = ~new_n8603_ & ~new_n8604_;
  assign new_n8606_ = new_n8519_ & ~new_n8605_;
  assign new_n8607_ = ~new_n8516_ & new_n8606_;
  assign new_n8608_ = ~new_n8601_ & ~new_n8607_;
  assign new_n8609_ = ~\b[25]  & ~new_n8608_;
  assign new_n8610_ = ~new_n8155_ & ~\quotient[30] ;
  assign new_n8611_ = ~new_n8165_ & new_n8464_;
  assign new_n8612_ = ~new_n8460_ & new_n8611_;
  assign new_n8613_ = ~new_n8461_ & ~new_n8464_;
  assign new_n8614_ = ~new_n8612_ & ~new_n8613_;
  assign new_n8615_ = new_n8519_ & ~new_n8614_;
  assign new_n8616_ = ~new_n8516_ & new_n8615_;
  assign new_n8617_ = ~new_n8610_ & ~new_n8616_;
  assign new_n8618_ = ~\b[24]  & ~new_n8617_;
  assign new_n8619_ = ~new_n8164_ & ~\quotient[30] ;
  assign new_n8620_ = ~new_n8174_ & new_n8459_;
  assign new_n8621_ = ~new_n8455_ & new_n8620_;
  assign new_n8622_ = ~new_n8456_ & ~new_n8459_;
  assign new_n8623_ = ~new_n8621_ & ~new_n8622_;
  assign new_n8624_ = new_n8519_ & ~new_n8623_;
  assign new_n8625_ = ~new_n8516_ & new_n8624_;
  assign new_n8626_ = ~new_n8619_ & ~new_n8625_;
  assign new_n8627_ = ~\b[23]  & ~new_n8626_;
  assign new_n8628_ = ~new_n8173_ & ~\quotient[30] ;
  assign new_n8629_ = ~new_n8183_ & new_n8454_;
  assign new_n8630_ = ~new_n8450_ & new_n8629_;
  assign new_n8631_ = ~new_n8451_ & ~new_n8454_;
  assign new_n8632_ = ~new_n8630_ & ~new_n8631_;
  assign new_n8633_ = new_n8519_ & ~new_n8632_;
  assign new_n8634_ = ~new_n8516_ & new_n8633_;
  assign new_n8635_ = ~new_n8628_ & ~new_n8634_;
  assign new_n8636_ = ~\b[22]  & ~new_n8635_;
  assign new_n8637_ = ~new_n8182_ & ~\quotient[30] ;
  assign new_n8638_ = ~new_n8192_ & new_n8449_;
  assign new_n8639_ = ~new_n8445_ & new_n8638_;
  assign new_n8640_ = ~new_n8446_ & ~new_n8449_;
  assign new_n8641_ = ~new_n8639_ & ~new_n8640_;
  assign new_n8642_ = new_n8519_ & ~new_n8641_;
  assign new_n8643_ = ~new_n8516_ & new_n8642_;
  assign new_n8644_ = ~new_n8637_ & ~new_n8643_;
  assign new_n8645_ = ~\b[21]  & ~new_n8644_;
  assign new_n8646_ = ~new_n8191_ & ~\quotient[30] ;
  assign new_n8647_ = ~new_n8201_ & new_n8444_;
  assign new_n8648_ = ~new_n8440_ & new_n8647_;
  assign new_n8649_ = ~new_n8441_ & ~new_n8444_;
  assign new_n8650_ = ~new_n8648_ & ~new_n8649_;
  assign new_n8651_ = new_n8519_ & ~new_n8650_;
  assign new_n8652_ = ~new_n8516_ & new_n8651_;
  assign new_n8653_ = ~new_n8646_ & ~new_n8652_;
  assign new_n8654_ = ~\b[20]  & ~new_n8653_;
  assign new_n8655_ = ~new_n8200_ & ~\quotient[30] ;
  assign new_n8656_ = ~new_n8210_ & new_n8439_;
  assign new_n8657_ = ~new_n8435_ & new_n8656_;
  assign new_n8658_ = ~new_n8436_ & ~new_n8439_;
  assign new_n8659_ = ~new_n8657_ & ~new_n8658_;
  assign new_n8660_ = new_n8519_ & ~new_n8659_;
  assign new_n8661_ = ~new_n8516_ & new_n8660_;
  assign new_n8662_ = ~new_n8655_ & ~new_n8661_;
  assign new_n8663_ = ~\b[19]  & ~new_n8662_;
  assign new_n8664_ = ~new_n8209_ & ~\quotient[30] ;
  assign new_n8665_ = ~new_n8219_ & new_n8434_;
  assign new_n8666_ = ~new_n8430_ & new_n8665_;
  assign new_n8667_ = ~new_n8431_ & ~new_n8434_;
  assign new_n8668_ = ~new_n8666_ & ~new_n8667_;
  assign new_n8669_ = new_n8519_ & ~new_n8668_;
  assign new_n8670_ = ~new_n8516_ & new_n8669_;
  assign new_n8671_ = ~new_n8664_ & ~new_n8670_;
  assign new_n8672_ = ~\b[18]  & ~new_n8671_;
  assign new_n8673_ = ~new_n8218_ & ~\quotient[30] ;
  assign new_n8674_ = ~new_n8228_ & new_n8429_;
  assign new_n8675_ = ~new_n8425_ & new_n8674_;
  assign new_n8676_ = ~new_n8426_ & ~new_n8429_;
  assign new_n8677_ = ~new_n8675_ & ~new_n8676_;
  assign new_n8678_ = new_n8519_ & ~new_n8677_;
  assign new_n8679_ = ~new_n8516_ & new_n8678_;
  assign new_n8680_ = ~new_n8673_ & ~new_n8679_;
  assign new_n8681_ = ~\b[17]  & ~new_n8680_;
  assign new_n8682_ = ~new_n8227_ & ~\quotient[30] ;
  assign new_n8683_ = ~new_n8237_ & new_n8424_;
  assign new_n8684_ = ~new_n8420_ & new_n8683_;
  assign new_n8685_ = ~new_n8421_ & ~new_n8424_;
  assign new_n8686_ = ~new_n8684_ & ~new_n8685_;
  assign new_n8687_ = new_n8519_ & ~new_n8686_;
  assign new_n8688_ = ~new_n8516_ & new_n8687_;
  assign new_n8689_ = ~new_n8682_ & ~new_n8688_;
  assign new_n8690_ = ~\b[16]  & ~new_n8689_;
  assign new_n8691_ = ~new_n8236_ & ~\quotient[30] ;
  assign new_n8692_ = ~new_n8246_ & new_n8419_;
  assign new_n8693_ = ~new_n8415_ & new_n8692_;
  assign new_n8694_ = ~new_n8416_ & ~new_n8419_;
  assign new_n8695_ = ~new_n8693_ & ~new_n8694_;
  assign new_n8696_ = new_n8519_ & ~new_n8695_;
  assign new_n8697_ = ~new_n8516_ & new_n8696_;
  assign new_n8698_ = ~new_n8691_ & ~new_n8697_;
  assign new_n8699_ = ~\b[15]  & ~new_n8698_;
  assign new_n8700_ = ~new_n8245_ & ~\quotient[30] ;
  assign new_n8701_ = ~new_n8255_ & new_n8414_;
  assign new_n8702_ = ~new_n8410_ & new_n8701_;
  assign new_n8703_ = ~new_n8411_ & ~new_n8414_;
  assign new_n8704_ = ~new_n8702_ & ~new_n8703_;
  assign new_n8705_ = new_n8519_ & ~new_n8704_;
  assign new_n8706_ = ~new_n8516_ & new_n8705_;
  assign new_n8707_ = ~new_n8700_ & ~new_n8706_;
  assign new_n8708_ = ~\b[14]  & ~new_n8707_;
  assign new_n8709_ = ~new_n8254_ & ~\quotient[30] ;
  assign new_n8710_ = ~new_n8264_ & new_n8409_;
  assign new_n8711_ = ~new_n8405_ & new_n8710_;
  assign new_n8712_ = ~new_n8406_ & ~new_n8409_;
  assign new_n8713_ = ~new_n8711_ & ~new_n8712_;
  assign new_n8714_ = new_n8519_ & ~new_n8713_;
  assign new_n8715_ = ~new_n8516_ & new_n8714_;
  assign new_n8716_ = ~new_n8709_ & ~new_n8715_;
  assign new_n8717_ = ~\b[13]  & ~new_n8716_;
  assign new_n8718_ = ~new_n8263_ & ~\quotient[30] ;
  assign new_n8719_ = ~new_n8273_ & new_n8404_;
  assign new_n8720_ = ~new_n8400_ & new_n8719_;
  assign new_n8721_ = ~new_n8401_ & ~new_n8404_;
  assign new_n8722_ = ~new_n8720_ & ~new_n8721_;
  assign new_n8723_ = new_n8519_ & ~new_n8722_;
  assign new_n8724_ = ~new_n8516_ & new_n8723_;
  assign new_n8725_ = ~new_n8718_ & ~new_n8724_;
  assign new_n8726_ = ~\b[12]  & ~new_n8725_;
  assign new_n8727_ = ~new_n8272_ & ~\quotient[30] ;
  assign new_n8728_ = ~new_n8282_ & new_n8399_;
  assign new_n8729_ = ~new_n8395_ & new_n8728_;
  assign new_n8730_ = ~new_n8396_ & ~new_n8399_;
  assign new_n8731_ = ~new_n8729_ & ~new_n8730_;
  assign new_n8732_ = new_n8519_ & ~new_n8731_;
  assign new_n8733_ = ~new_n8516_ & new_n8732_;
  assign new_n8734_ = ~new_n8727_ & ~new_n8733_;
  assign new_n8735_ = ~\b[11]  & ~new_n8734_;
  assign new_n8736_ = ~new_n8281_ & ~\quotient[30] ;
  assign new_n8737_ = ~new_n8291_ & new_n8394_;
  assign new_n8738_ = ~new_n8390_ & new_n8737_;
  assign new_n8739_ = ~new_n8391_ & ~new_n8394_;
  assign new_n8740_ = ~new_n8738_ & ~new_n8739_;
  assign new_n8741_ = new_n8519_ & ~new_n8740_;
  assign new_n8742_ = ~new_n8516_ & new_n8741_;
  assign new_n8743_ = ~new_n8736_ & ~new_n8742_;
  assign new_n8744_ = ~\b[10]  & ~new_n8743_;
  assign new_n8745_ = ~new_n8290_ & ~\quotient[30] ;
  assign new_n8746_ = ~new_n8300_ & new_n8389_;
  assign new_n8747_ = ~new_n8385_ & new_n8746_;
  assign new_n8748_ = ~new_n8386_ & ~new_n8389_;
  assign new_n8749_ = ~new_n8747_ & ~new_n8748_;
  assign new_n8750_ = new_n8519_ & ~new_n8749_;
  assign new_n8751_ = ~new_n8516_ & new_n8750_;
  assign new_n8752_ = ~new_n8745_ & ~new_n8751_;
  assign new_n8753_ = ~\b[9]  & ~new_n8752_;
  assign new_n8754_ = ~new_n8299_ & ~\quotient[30] ;
  assign new_n8755_ = ~new_n8309_ & new_n8384_;
  assign new_n8756_ = ~new_n8380_ & new_n8755_;
  assign new_n8757_ = ~new_n8381_ & ~new_n8384_;
  assign new_n8758_ = ~new_n8756_ & ~new_n8757_;
  assign new_n8759_ = new_n8519_ & ~new_n8758_;
  assign new_n8760_ = ~new_n8516_ & new_n8759_;
  assign new_n8761_ = ~new_n8754_ & ~new_n8760_;
  assign new_n8762_ = ~\b[8]  & ~new_n8761_;
  assign new_n8763_ = ~new_n8308_ & ~\quotient[30] ;
  assign new_n8764_ = ~new_n8318_ & new_n8379_;
  assign new_n8765_ = ~new_n8375_ & new_n8764_;
  assign new_n8766_ = ~new_n8376_ & ~new_n8379_;
  assign new_n8767_ = ~new_n8765_ & ~new_n8766_;
  assign new_n8768_ = new_n8519_ & ~new_n8767_;
  assign new_n8769_ = ~new_n8516_ & new_n8768_;
  assign new_n8770_ = ~new_n8763_ & ~new_n8769_;
  assign new_n8771_ = ~\b[7]  & ~new_n8770_;
  assign new_n8772_ = ~new_n8317_ & ~\quotient[30] ;
  assign new_n8773_ = ~new_n8327_ & new_n8374_;
  assign new_n8774_ = ~new_n8370_ & new_n8773_;
  assign new_n8775_ = ~new_n8371_ & ~new_n8374_;
  assign new_n8776_ = ~new_n8774_ & ~new_n8775_;
  assign new_n8777_ = new_n8519_ & ~new_n8776_;
  assign new_n8778_ = ~new_n8516_ & new_n8777_;
  assign new_n8779_ = ~new_n8772_ & ~new_n8778_;
  assign new_n8780_ = ~\b[6]  & ~new_n8779_;
  assign new_n8781_ = ~new_n8326_ & ~\quotient[30] ;
  assign new_n8782_ = ~new_n8336_ & new_n8369_;
  assign new_n8783_ = ~new_n8365_ & new_n8782_;
  assign new_n8784_ = ~new_n8366_ & ~new_n8369_;
  assign new_n8785_ = ~new_n8783_ & ~new_n8784_;
  assign new_n8786_ = new_n8519_ & ~new_n8785_;
  assign new_n8787_ = ~new_n8516_ & new_n8786_;
  assign new_n8788_ = ~new_n8781_ & ~new_n8787_;
  assign new_n8789_ = ~\b[5]  & ~new_n8788_;
  assign new_n8790_ = ~new_n8335_ & ~\quotient[30] ;
  assign new_n8791_ = ~new_n8344_ & new_n8364_;
  assign new_n8792_ = ~new_n8360_ & new_n8791_;
  assign new_n8793_ = ~new_n8361_ & ~new_n8364_;
  assign new_n8794_ = ~new_n8792_ & ~new_n8793_;
  assign new_n8795_ = new_n8519_ & ~new_n8794_;
  assign new_n8796_ = ~new_n8516_ & new_n8795_;
  assign new_n8797_ = ~new_n8790_ & ~new_n8796_;
  assign new_n8798_ = ~\b[4]  & ~new_n8797_;
  assign new_n8799_ = ~new_n8343_ & ~\quotient[30] ;
  assign new_n8800_ = ~new_n8355_ & new_n8359_;
  assign new_n8801_ = ~new_n8354_ & new_n8800_;
  assign new_n8802_ = ~new_n8356_ & ~new_n8359_;
  assign new_n8803_ = ~new_n8801_ & ~new_n8802_;
  assign new_n8804_ = new_n8519_ & ~new_n8803_;
  assign new_n8805_ = ~new_n8516_ & new_n8804_;
  assign new_n8806_ = ~new_n8799_ & ~new_n8805_;
  assign new_n8807_ = ~\b[3]  & ~new_n8806_;
  assign new_n8808_ = ~new_n8348_ & ~\quotient[30] ;
  assign new_n8809_ = ~new_n8351_ & new_n8353_;
  assign new_n8810_ = ~new_n8349_ & new_n8809_;
  assign new_n8811_ = new_n8519_ & ~new_n8810_;
  assign new_n8812_ = ~new_n8354_ & new_n8811_;
  assign new_n8813_ = ~new_n8516_ & new_n8812_;
  assign new_n8814_ = ~new_n8808_ & ~new_n8813_;
  assign new_n8815_ = ~\b[2]  & ~new_n8814_;
  assign new_n8816_ = \b[0]  & ~\b[34] ;
  assign new_n8817_ = new_n413_ & new_n8816_;
  assign new_n8818_ = new_n411_ & new_n8817_;
  assign new_n8819_ = new_n422_ & new_n8818_;
  assign new_n8820_ = new_n408_ & new_n8819_;
  assign new_n8821_ = ~new_n8516_ & new_n8820_;
  assign new_n8822_ = \a[30]  & ~new_n8821_;
  assign new_n8823_ = new_n312_ & new_n8353_;
  assign new_n8824_ = new_n294_ & new_n8823_;
  assign new_n8825_ = new_n340_ & new_n8824_;
  assign new_n8826_ = new_n338_ & new_n8825_;
  assign new_n8827_ = ~new_n8516_ & new_n8826_;
  assign new_n8828_ = ~new_n8822_ & ~new_n8827_;
  assign new_n8829_ = \b[1]  & ~new_n8828_;
  assign new_n8830_ = ~\b[1]  & ~new_n8827_;
  assign new_n8831_ = ~new_n8822_ & new_n8830_;
  assign new_n8832_ = ~new_n8829_ & ~new_n8831_;
  assign new_n8833_ = ~\a[29]  & \b[0] ;
  assign new_n8834_ = ~new_n8832_ & ~new_n8833_;
  assign new_n8835_ = ~\b[1]  & ~new_n8828_;
  assign new_n8836_ = ~new_n8834_ & ~new_n8835_;
  assign new_n8837_ = \b[2]  & ~new_n8813_;
  assign new_n8838_ = ~new_n8808_ & new_n8837_;
  assign new_n8839_ = ~new_n8815_ & ~new_n8838_;
  assign new_n8840_ = ~new_n8836_ & new_n8839_;
  assign new_n8841_ = ~new_n8815_ & ~new_n8840_;
  assign new_n8842_ = \b[3]  & ~new_n8805_;
  assign new_n8843_ = ~new_n8799_ & new_n8842_;
  assign new_n8844_ = ~new_n8807_ & ~new_n8843_;
  assign new_n8845_ = ~new_n8841_ & new_n8844_;
  assign new_n8846_ = ~new_n8807_ & ~new_n8845_;
  assign new_n8847_ = \b[4]  & ~new_n8796_;
  assign new_n8848_ = ~new_n8790_ & new_n8847_;
  assign new_n8849_ = ~new_n8798_ & ~new_n8848_;
  assign new_n8850_ = ~new_n8846_ & new_n8849_;
  assign new_n8851_ = ~new_n8798_ & ~new_n8850_;
  assign new_n8852_ = \b[5]  & ~new_n8787_;
  assign new_n8853_ = ~new_n8781_ & new_n8852_;
  assign new_n8854_ = ~new_n8789_ & ~new_n8853_;
  assign new_n8855_ = ~new_n8851_ & new_n8854_;
  assign new_n8856_ = ~new_n8789_ & ~new_n8855_;
  assign new_n8857_ = \b[6]  & ~new_n8778_;
  assign new_n8858_ = ~new_n8772_ & new_n8857_;
  assign new_n8859_ = ~new_n8780_ & ~new_n8858_;
  assign new_n8860_ = ~new_n8856_ & new_n8859_;
  assign new_n8861_ = ~new_n8780_ & ~new_n8860_;
  assign new_n8862_ = \b[7]  & ~new_n8769_;
  assign new_n8863_ = ~new_n8763_ & new_n8862_;
  assign new_n8864_ = ~new_n8771_ & ~new_n8863_;
  assign new_n8865_ = ~new_n8861_ & new_n8864_;
  assign new_n8866_ = ~new_n8771_ & ~new_n8865_;
  assign new_n8867_ = \b[8]  & ~new_n8760_;
  assign new_n8868_ = ~new_n8754_ & new_n8867_;
  assign new_n8869_ = ~new_n8762_ & ~new_n8868_;
  assign new_n8870_ = ~new_n8866_ & new_n8869_;
  assign new_n8871_ = ~new_n8762_ & ~new_n8870_;
  assign new_n8872_ = \b[9]  & ~new_n8751_;
  assign new_n8873_ = ~new_n8745_ & new_n8872_;
  assign new_n8874_ = ~new_n8753_ & ~new_n8873_;
  assign new_n8875_ = ~new_n8871_ & new_n8874_;
  assign new_n8876_ = ~new_n8753_ & ~new_n8875_;
  assign new_n8877_ = \b[10]  & ~new_n8742_;
  assign new_n8878_ = ~new_n8736_ & new_n8877_;
  assign new_n8879_ = ~new_n8744_ & ~new_n8878_;
  assign new_n8880_ = ~new_n8876_ & new_n8879_;
  assign new_n8881_ = ~new_n8744_ & ~new_n8880_;
  assign new_n8882_ = \b[11]  & ~new_n8733_;
  assign new_n8883_ = ~new_n8727_ & new_n8882_;
  assign new_n8884_ = ~new_n8735_ & ~new_n8883_;
  assign new_n8885_ = ~new_n8881_ & new_n8884_;
  assign new_n8886_ = ~new_n8735_ & ~new_n8885_;
  assign new_n8887_ = \b[12]  & ~new_n8724_;
  assign new_n8888_ = ~new_n8718_ & new_n8887_;
  assign new_n8889_ = ~new_n8726_ & ~new_n8888_;
  assign new_n8890_ = ~new_n8886_ & new_n8889_;
  assign new_n8891_ = ~new_n8726_ & ~new_n8890_;
  assign new_n8892_ = \b[13]  & ~new_n8715_;
  assign new_n8893_ = ~new_n8709_ & new_n8892_;
  assign new_n8894_ = ~new_n8717_ & ~new_n8893_;
  assign new_n8895_ = ~new_n8891_ & new_n8894_;
  assign new_n8896_ = ~new_n8717_ & ~new_n8895_;
  assign new_n8897_ = \b[14]  & ~new_n8706_;
  assign new_n8898_ = ~new_n8700_ & new_n8897_;
  assign new_n8899_ = ~new_n8708_ & ~new_n8898_;
  assign new_n8900_ = ~new_n8896_ & new_n8899_;
  assign new_n8901_ = ~new_n8708_ & ~new_n8900_;
  assign new_n8902_ = \b[15]  & ~new_n8697_;
  assign new_n8903_ = ~new_n8691_ & new_n8902_;
  assign new_n8904_ = ~new_n8699_ & ~new_n8903_;
  assign new_n8905_ = ~new_n8901_ & new_n8904_;
  assign new_n8906_ = ~new_n8699_ & ~new_n8905_;
  assign new_n8907_ = \b[16]  & ~new_n8688_;
  assign new_n8908_ = ~new_n8682_ & new_n8907_;
  assign new_n8909_ = ~new_n8690_ & ~new_n8908_;
  assign new_n8910_ = ~new_n8906_ & new_n8909_;
  assign new_n8911_ = ~new_n8690_ & ~new_n8910_;
  assign new_n8912_ = \b[17]  & ~new_n8679_;
  assign new_n8913_ = ~new_n8673_ & new_n8912_;
  assign new_n8914_ = ~new_n8681_ & ~new_n8913_;
  assign new_n8915_ = ~new_n8911_ & new_n8914_;
  assign new_n8916_ = ~new_n8681_ & ~new_n8915_;
  assign new_n8917_ = \b[18]  & ~new_n8670_;
  assign new_n8918_ = ~new_n8664_ & new_n8917_;
  assign new_n8919_ = ~new_n8672_ & ~new_n8918_;
  assign new_n8920_ = ~new_n8916_ & new_n8919_;
  assign new_n8921_ = ~new_n8672_ & ~new_n8920_;
  assign new_n8922_ = \b[19]  & ~new_n8661_;
  assign new_n8923_ = ~new_n8655_ & new_n8922_;
  assign new_n8924_ = ~new_n8663_ & ~new_n8923_;
  assign new_n8925_ = ~new_n8921_ & new_n8924_;
  assign new_n8926_ = ~new_n8663_ & ~new_n8925_;
  assign new_n8927_ = \b[20]  & ~new_n8652_;
  assign new_n8928_ = ~new_n8646_ & new_n8927_;
  assign new_n8929_ = ~new_n8654_ & ~new_n8928_;
  assign new_n8930_ = ~new_n8926_ & new_n8929_;
  assign new_n8931_ = ~new_n8654_ & ~new_n8930_;
  assign new_n8932_ = \b[21]  & ~new_n8643_;
  assign new_n8933_ = ~new_n8637_ & new_n8932_;
  assign new_n8934_ = ~new_n8645_ & ~new_n8933_;
  assign new_n8935_ = ~new_n8931_ & new_n8934_;
  assign new_n8936_ = ~new_n8645_ & ~new_n8935_;
  assign new_n8937_ = \b[22]  & ~new_n8634_;
  assign new_n8938_ = ~new_n8628_ & new_n8937_;
  assign new_n8939_ = ~new_n8636_ & ~new_n8938_;
  assign new_n8940_ = ~new_n8936_ & new_n8939_;
  assign new_n8941_ = ~new_n8636_ & ~new_n8940_;
  assign new_n8942_ = \b[23]  & ~new_n8625_;
  assign new_n8943_ = ~new_n8619_ & new_n8942_;
  assign new_n8944_ = ~new_n8627_ & ~new_n8943_;
  assign new_n8945_ = ~new_n8941_ & new_n8944_;
  assign new_n8946_ = ~new_n8627_ & ~new_n8945_;
  assign new_n8947_ = \b[24]  & ~new_n8616_;
  assign new_n8948_ = ~new_n8610_ & new_n8947_;
  assign new_n8949_ = ~new_n8618_ & ~new_n8948_;
  assign new_n8950_ = ~new_n8946_ & new_n8949_;
  assign new_n8951_ = ~new_n8618_ & ~new_n8950_;
  assign new_n8952_ = \b[25]  & ~new_n8607_;
  assign new_n8953_ = ~new_n8601_ & new_n8952_;
  assign new_n8954_ = ~new_n8609_ & ~new_n8953_;
  assign new_n8955_ = ~new_n8951_ & new_n8954_;
  assign new_n8956_ = ~new_n8609_ & ~new_n8955_;
  assign new_n8957_ = \b[26]  & ~new_n8598_;
  assign new_n8958_ = ~new_n8592_ & new_n8957_;
  assign new_n8959_ = ~new_n8600_ & ~new_n8958_;
  assign new_n8960_ = ~new_n8956_ & new_n8959_;
  assign new_n8961_ = ~new_n8600_ & ~new_n8960_;
  assign new_n8962_ = \b[27]  & ~new_n8589_;
  assign new_n8963_ = ~new_n8583_ & new_n8962_;
  assign new_n8964_ = ~new_n8591_ & ~new_n8963_;
  assign new_n8965_ = ~new_n8961_ & new_n8964_;
  assign new_n8966_ = ~new_n8591_ & ~new_n8965_;
  assign new_n8967_ = \b[28]  & ~new_n8580_;
  assign new_n8968_ = ~new_n8574_ & new_n8967_;
  assign new_n8969_ = ~new_n8582_ & ~new_n8968_;
  assign new_n8970_ = ~new_n8966_ & new_n8969_;
  assign new_n8971_ = ~new_n8582_ & ~new_n8970_;
  assign new_n8972_ = \b[29]  & ~new_n8571_;
  assign new_n8973_ = ~new_n8565_ & new_n8972_;
  assign new_n8974_ = ~new_n8573_ & ~new_n8973_;
  assign new_n8975_ = ~new_n8971_ & new_n8974_;
  assign new_n8976_ = ~new_n8573_ & ~new_n8975_;
  assign new_n8977_ = \b[30]  & ~new_n8562_;
  assign new_n8978_ = ~new_n8556_ & new_n8977_;
  assign new_n8979_ = ~new_n8564_ & ~new_n8978_;
  assign new_n8980_ = ~new_n8976_ & new_n8979_;
  assign new_n8981_ = ~new_n8564_ & ~new_n8980_;
  assign new_n8982_ = \b[31]  & ~new_n8553_;
  assign new_n8983_ = ~new_n8547_ & new_n8982_;
  assign new_n8984_ = ~new_n8555_ & ~new_n8983_;
  assign new_n8985_ = ~new_n8981_ & new_n8984_;
  assign new_n8986_ = ~new_n8555_ & ~new_n8985_;
  assign new_n8987_ = \b[32]  & ~new_n8544_;
  assign new_n8988_ = ~new_n8538_ & new_n8987_;
  assign new_n8989_ = ~new_n8546_ & ~new_n8988_;
  assign new_n8990_ = ~new_n8986_ & new_n8989_;
  assign new_n8991_ = ~new_n8546_ & ~new_n8990_;
  assign new_n8992_ = \b[33]  & ~new_n8527_;
  assign new_n8993_ = ~new_n8521_ & new_n8992_;
  assign new_n8994_ = ~new_n8537_ & ~new_n8993_;
  assign new_n8995_ = ~new_n8991_ & new_n8994_;
  assign new_n8996_ = ~new_n8537_ & ~new_n8995_;
  assign new_n8997_ = \b[34]  & ~new_n8529_;
  assign new_n8998_ = ~new_n8534_ & new_n8997_;
  assign new_n8999_ = ~new_n8536_ & ~new_n8998_;
  assign new_n9000_ = ~new_n8996_ & new_n8999_;
  assign new_n9001_ = ~new_n8536_ & ~new_n9000_;
  assign new_n9002_ = new_n411_ & new_n413_;
  assign new_n9003_ = new_n422_ & new_n9002_;
  assign new_n9004_ = new_n408_ & new_n9003_;
  assign \quotient[29]  = ~new_n9001_ & new_n9004_;
  assign new_n9006_ = ~new_n8528_ & ~\quotient[29] ;
  assign new_n9007_ = ~new_n8546_ & new_n8994_;
  assign new_n9008_ = ~new_n8990_ & new_n9007_;
  assign new_n9009_ = ~new_n8991_ & ~new_n8994_;
  assign new_n9010_ = ~new_n9008_ & ~new_n9009_;
  assign new_n9011_ = new_n9004_ & ~new_n9010_;
  assign new_n9012_ = ~new_n9001_ & new_n9011_;
  assign new_n9013_ = ~new_n9006_ & ~new_n9012_;
  assign new_n9014_ = ~\b[34]  & ~new_n9013_;
  assign new_n9015_ = ~new_n8545_ & ~\quotient[29] ;
  assign new_n9016_ = ~new_n8555_ & new_n8989_;
  assign new_n9017_ = ~new_n8985_ & new_n9016_;
  assign new_n9018_ = ~new_n8986_ & ~new_n8989_;
  assign new_n9019_ = ~new_n9017_ & ~new_n9018_;
  assign new_n9020_ = new_n9004_ & ~new_n9019_;
  assign new_n9021_ = ~new_n9001_ & new_n9020_;
  assign new_n9022_ = ~new_n9015_ & ~new_n9021_;
  assign new_n9023_ = ~\b[33]  & ~new_n9022_;
  assign new_n9024_ = ~new_n8554_ & ~\quotient[29] ;
  assign new_n9025_ = ~new_n8564_ & new_n8984_;
  assign new_n9026_ = ~new_n8980_ & new_n9025_;
  assign new_n9027_ = ~new_n8981_ & ~new_n8984_;
  assign new_n9028_ = ~new_n9026_ & ~new_n9027_;
  assign new_n9029_ = new_n9004_ & ~new_n9028_;
  assign new_n9030_ = ~new_n9001_ & new_n9029_;
  assign new_n9031_ = ~new_n9024_ & ~new_n9030_;
  assign new_n9032_ = ~\b[32]  & ~new_n9031_;
  assign new_n9033_ = ~new_n8563_ & ~\quotient[29] ;
  assign new_n9034_ = ~new_n8573_ & new_n8979_;
  assign new_n9035_ = ~new_n8975_ & new_n9034_;
  assign new_n9036_ = ~new_n8976_ & ~new_n8979_;
  assign new_n9037_ = ~new_n9035_ & ~new_n9036_;
  assign new_n9038_ = new_n9004_ & ~new_n9037_;
  assign new_n9039_ = ~new_n9001_ & new_n9038_;
  assign new_n9040_ = ~new_n9033_ & ~new_n9039_;
  assign new_n9041_ = ~\b[31]  & ~new_n9040_;
  assign new_n9042_ = ~new_n8572_ & ~\quotient[29] ;
  assign new_n9043_ = ~new_n8582_ & new_n8974_;
  assign new_n9044_ = ~new_n8970_ & new_n9043_;
  assign new_n9045_ = ~new_n8971_ & ~new_n8974_;
  assign new_n9046_ = ~new_n9044_ & ~new_n9045_;
  assign new_n9047_ = new_n9004_ & ~new_n9046_;
  assign new_n9048_ = ~new_n9001_ & new_n9047_;
  assign new_n9049_ = ~new_n9042_ & ~new_n9048_;
  assign new_n9050_ = ~\b[30]  & ~new_n9049_;
  assign new_n9051_ = ~new_n8581_ & ~\quotient[29] ;
  assign new_n9052_ = ~new_n8591_ & new_n8969_;
  assign new_n9053_ = ~new_n8965_ & new_n9052_;
  assign new_n9054_ = ~new_n8966_ & ~new_n8969_;
  assign new_n9055_ = ~new_n9053_ & ~new_n9054_;
  assign new_n9056_ = new_n9004_ & ~new_n9055_;
  assign new_n9057_ = ~new_n9001_ & new_n9056_;
  assign new_n9058_ = ~new_n9051_ & ~new_n9057_;
  assign new_n9059_ = ~\b[29]  & ~new_n9058_;
  assign new_n9060_ = ~new_n8590_ & ~\quotient[29] ;
  assign new_n9061_ = ~new_n8600_ & new_n8964_;
  assign new_n9062_ = ~new_n8960_ & new_n9061_;
  assign new_n9063_ = ~new_n8961_ & ~new_n8964_;
  assign new_n9064_ = ~new_n9062_ & ~new_n9063_;
  assign new_n9065_ = new_n9004_ & ~new_n9064_;
  assign new_n9066_ = ~new_n9001_ & new_n9065_;
  assign new_n9067_ = ~new_n9060_ & ~new_n9066_;
  assign new_n9068_ = ~\b[28]  & ~new_n9067_;
  assign new_n9069_ = ~new_n8599_ & ~\quotient[29] ;
  assign new_n9070_ = ~new_n8609_ & new_n8959_;
  assign new_n9071_ = ~new_n8955_ & new_n9070_;
  assign new_n9072_ = ~new_n8956_ & ~new_n8959_;
  assign new_n9073_ = ~new_n9071_ & ~new_n9072_;
  assign new_n9074_ = new_n9004_ & ~new_n9073_;
  assign new_n9075_ = ~new_n9001_ & new_n9074_;
  assign new_n9076_ = ~new_n9069_ & ~new_n9075_;
  assign new_n9077_ = ~\b[27]  & ~new_n9076_;
  assign new_n9078_ = ~new_n8608_ & ~\quotient[29] ;
  assign new_n9079_ = ~new_n8618_ & new_n8954_;
  assign new_n9080_ = ~new_n8950_ & new_n9079_;
  assign new_n9081_ = ~new_n8951_ & ~new_n8954_;
  assign new_n9082_ = ~new_n9080_ & ~new_n9081_;
  assign new_n9083_ = new_n9004_ & ~new_n9082_;
  assign new_n9084_ = ~new_n9001_ & new_n9083_;
  assign new_n9085_ = ~new_n9078_ & ~new_n9084_;
  assign new_n9086_ = ~\b[26]  & ~new_n9085_;
  assign new_n9087_ = ~new_n8617_ & ~\quotient[29] ;
  assign new_n9088_ = ~new_n8627_ & new_n8949_;
  assign new_n9089_ = ~new_n8945_ & new_n9088_;
  assign new_n9090_ = ~new_n8946_ & ~new_n8949_;
  assign new_n9091_ = ~new_n9089_ & ~new_n9090_;
  assign new_n9092_ = new_n9004_ & ~new_n9091_;
  assign new_n9093_ = ~new_n9001_ & new_n9092_;
  assign new_n9094_ = ~new_n9087_ & ~new_n9093_;
  assign new_n9095_ = ~\b[25]  & ~new_n9094_;
  assign new_n9096_ = ~new_n8626_ & ~\quotient[29] ;
  assign new_n9097_ = ~new_n8636_ & new_n8944_;
  assign new_n9098_ = ~new_n8940_ & new_n9097_;
  assign new_n9099_ = ~new_n8941_ & ~new_n8944_;
  assign new_n9100_ = ~new_n9098_ & ~new_n9099_;
  assign new_n9101_ = new_n9004_ & ~new_n9100_;
  assign new_n9102_ = ~new_n9001_ & new_n9101_;
  assign new_n9103_ = ~new_n9096_ & ~new_n9102_;
  assign new_n9104_ = ~\b[24]  & ~new_n9103_;
  assign new_n9105_ = ~new_n8635_ & ~\quotient[29] ;
  assign new_n9106_ = ~new_n8645_ & new_n8939_;
  assign new_n9107_ = ~new_n8935_ & new_n9106_;
  assign new_n9108_ = ~new_n8936_ & ~new_n8939_;
  assign new_n9109_ = ~new_n9107_ & ~new_n9108_;
  assign new_n9110_ = new_n9004_ & ~new_n9109_;
  assign new_n9111_ = ~new_n9001_ & new_n9110_;
  assign new_n9112_ = ~new_n9105_ & ~new_n9111_;
  assign new_n9113_ = ~\b[23]  & ~new_n9112_;
  assign new_n9114_ = ~new_n8644_ & ~\quotient[29] ;
  assign new_n9115_ = ~new_n8654_ & new_n8934_;
  assign new_n9116_ = ~new_n8930_ & new_n9115_;
  assign new_n9117_ = ~new_n8931_ & ~new_n8934_;
  assign new_n9118_ = ~new_n9116_ & ~new_n9117_;
  assign new_n9119_ = new_n9004_ & ~new_n9118_;
  assign new_n9120_ = ~new_n9001_ & new_n9119_;
  assign new_n9121_ = ~new_n9114_ & ~new_n9120_;
  assign new_n9122_ = ~\b[22]  & ~new_n9121_;
  assign new_n9123_ = ~new_n8653_ & ~\quotient[29] ;
  assign new_n9124_ = ~new_n8663_ & new_n8929_;
  assign new_n9125_ = ~new_n8925_ & new_n9124_;
  assign new_n9126_ = ~new_n8926_ & ~new_n8929_;
  assign new_n9127_ = ~new_n9125_ & ~new_n9126_;
  assign new_n9128_ = new_n9004_ & ~new_n9127_;
  assign new_n9129_ = ~new_n9001_ & new_n9128_;
  assign new_n9130_ = ~new_n9123_ & ~new_n9129_;
  assign new_n9131_ = ~\b[21]  & ~new_n9130_;
  assign new_n9132_ = ~new_n8662_ & ~\quotient[29] ;
  assign new_n9133_ = ~new_n8672_ & new_n8924_;
  assign new_n9134_ = ~new_n8920_ & new_n9133_;
  assign new_n9135_ = ~new_n8921_ & ~new_n8924_;
  assign new_n9136_ = ~new_n9134_ & ~new_n9135_;
  assign new_n9137_ = new_n9004_ & ~new_n9136_;
  assign new_n9138_ = ~new_n9001_ & new_n9137_;
  assign new_n9139_ = ~new_n9132_ & ~new_n9138_;
  assign new_n9140_ = ~\b[20]  & ~new_n9139_;
  assign new_n9141_ = ~new_n8671_ & ~\quotient[29] ;
  assign new_n9142_ = ~new_n8681_ & new_n8919_;
  assign new_n9143_ = ~new_n8915_ & new_n9142_;
  assign new_n9144_ = ~new_n8916_ & ~new_n8919_;
  assign new_n9145_ = ~new_n9143_ & ~new_n9144_;
  assign new_n9146_ = new_n9004_ & ~new_n9145_;
  assign new_n9147_ = ~new_n9001_ & new_n9146_;
  assign new_n9148_ = ~new_n9141_ & ~new_n9147_;
  assign new_n9149_ = ~\b[19]  & ~new_n9148_;
  assign new_n9150_ = ~new_n8680_ & ~\quotient[29] ;
  assign new_n9151_ = ~new_n8690_ & new_n8914_;
  assign new_n9152_ = ~new_n8910_ & new_n9151_;
  assign new_n9153_ = ~new_n8911_ & ~new_n8914_;
  assign new_n9154_ = ~new_n9152_ & ~new_n9153_;
  assign new_n9155_ = new_n9004_ & ~new_n9154_;
  assign new_n9156_ = ~new_n9001_ & new_n9155_;
  assign new_n9157_ = ~new_n9150_ & ~new_n9156_;
  assign new_n9158_ = ~\b[18]  & ~new_n9157_;
  assign new_n9159_ = ~new_n8689_ & ~\quotient[29] ;
  assign new_n9160_ = ~new_n8699_ & new_n8909_;
  assign new_n9161_ = ~new_n8905_ & new_n9160_;
  assign new_n9162_ = ~new_n8906_ & ~new_n8909_;
  assign new_n9163_ = ~new_n9161_ & ~new_n9162_;
  assign new_n9164_ = new_n9004_ & ~new_n9163_;
  assign new_n9165_ = ~new_n9001_ & new_n9164_;
  assign new_n9166_ = ~new_n9159_ & ~new_n9165_;
  assign new_n9167_ = ~\b[17]  & ~new_n9166_;
  assign new_n9168_ = ~new_n8698_ & ~\quotient[29] ;
  assign new_n9169_ = ~new_n8708_ & new_n8904_;
  assign new_n9170_ = ~new_n8900_ & new_n9169_;
  assign new_n9171_ = ~new_n8901_ & ~new_n8904_;
  assign new_n9172_ = ~new_n9170_ & ~new_n9171_;
  assign new_n9173_ = new_n9004_ & ~new_n9172_;
  assign new_n9174_ = ~new_n9001_ & new_n9173_;
  assign new_n9175_ = ~new_n9168_ & ~new_n9174_;
  assign new_n9176_ = ~\b[16]  & ~new_n9175_;
  assign new_n9177_ = ~new_n8707_ & ~\quotient[29] ;
  assign new_n9178_ = ~new_n8717_ & new_n8899_;
  assign new_n9179_ = ~new_n8895_ & new_n9178_;
  assign new_n9180_ = ~new_n8896_ & ~new_n8899_;
  assign new_n9181_ = ~new_n9179_ & ~new_n9180_;
  assign new_n9182_ = new_n9004_ & ~new_n9181_;
  assign new_n9183_ = ~new_n9001_ & new_n9182_;
  assign new_n9184_ = ~new_n9177_ & ~new_n9183_;
  assign new_n9185_ = ~\b[15]  & ~new_n9184_;
  assign new_n9186_ = ~new_n8716_ & ~\quotient[29] ;
  assign new_n9187_ = ~new_n8726_ & new_n8894_;
  assign new_n9188_ = ~new_n8890_ & new_n9187_;
  assign new_n9189_ = ~new_n8891_ & ~new_n8894_;
  assign new_n9190_ = ~new_n9188_ & ~new_n9189_;
  assign new_n9191_ = new_n9004_ & ~new_n9190_;
  assign new_n9192_ = ~new_n9001_ & new_n9191_;
  assign new_n9193_ = ~new_n9186_ & ~new_n9192_;
  assign new_n9194_ = ~\b[14]  & ~new_n9193_;
  assign new_n9195_ = ~new_n8725_ & ~\quotient[29] ;
  assign new_n9196_ = ~new_n8735_ & new_n8889_;
  assign new_n9197_ = ~new_n8885_ & new_n9196_;
  assign new_n9198_ = ~new_n8886_ & ~new_n8889_;
  assign new_n9199_ = ~new_n9197_ & ~new_n9198_;
  assign new_n9200_ = new_n9004_ & ~new_n9199_;
  assign new_n9201_ = ~new_n9001_ & new_n9200_;
  assign new_n9202_ = ~new_n9195_ & ~new_n9201_;
  assign new_n9203_ = ~\b[13]  & ~new_n9202_;
  assign new_n9204_ = ~new_n8734_ & ~\quotient[29] ;
  assign new_n9205_ = ~new_n8744_ & new_n8884_;
  assign new_n9206_ = ~new_n8880_ & new_n9205_;
  assign new_n9207_ = ~new_n8881_ & ~new_n8884_;
  assign new_n9208_ = ~new_n9206_ & ~new_n9207_;
  assign new_n9209_ = new_n9004_ & ~new_n9208_;
  assign new_n9210_ = ~new_n9001_ & new_n9209_;
  assign new_n9211_ = ~new_n9204_ & ~new_n9210_;
  assign new_n9212_ = ~\b[12]  & ~new_n9211_;
  assign new_n9213_ = ~new_n8743_ & ~\quotient[29] ;
  assign new_n9214_ = ~new_n8753_ & new_n8879_;
  assign new_n9215_ = ~new_n8875_ & new_n9214_;
  assign new_n9216_ = ~new_n8876_ & ~new_n8879_;
  assign new_n9217_ = ~new_n9215_ & ~new_n9216_;
  assign new_n9218_ = new_n9004_ & ~new_n9217_;
  assign new_n9219_ = ~new_n9001_ & new_n9218_;
  assign new_n9220_ = ~new_n9213_ & ~new_n9219_;
  assign new_n9221_ = ~\b[11]  & ~new_n9220_;
  assign new_n9222_ = ~new_n8752_ & ~\quotient[29] ;
  assign new_n9223_ = ~new_n8762_ & new_n8874_;
  assign new_n9224_ = ~new_n8870_ & new_n9223_;
  assign new_n9225_ = ~new_n8871_ & ~new_n8874_;
  assign new_n9226_ = ~new_n9224_ & ~new_n9225_;
  assign new_n9227_ = new_n9004_ & ~new_n9226_;
  assign new_n9228_ = ~new_n9001_ & new_n9227_;
  assign new_n9229_ = ~new_n9222_ & ~new_n9228_;
  assign new_n9230_ = ~\b[10]  & ~new_n9229_;
  assign new_n9231_ = ~new_n8761_ & ~\quotient[29] ;
  assign new_n9232_ = ~new_n8771_ & new_n8869_;
  assign new_n9233_ = ~new_n8865_ & new_n9232_;
  assign new_n9234_ = ~new_n8866_ & ~new_n8869_;
  assign new_n9235_ = ~new_n9233_ & ~new_n9234_;
  assign new_n9236_ = new_n9004_ & ~new_n9235_;
  assign new_n9237_ = ~new_n9001_ & new_n9236_;
  assign new_n9238_ = ~new_n9231_ & ~new_n9237_;
  assign new_n9239_ = ~\b[9]  & ~new_n9238_;
  assign new_n9240_ = ~new_n8770_ & ~\quotient[29] ;
  assign new_n9241_ = ~new_n8780_ & new_n8864_;
  assign new_n9242_ = ~new_n8860_ & new_n9241_;
  assign new_n9243_ = ~new_n8861_ & ~new_n8864_;
  assign new_n9244_ = ~new_n9242_ & ~new_n9243_;
  assign new_n9245_ = new_n9004_ & ~new_n9244_;
  assign new_n9246_ = ~new_n9001_ & new_n9245_;
  assign new_n9247_ = ~new_n9240_ & ~new_n9246_;
  assign new_n9248_ = ~\b[8]  & ~new_n9247_;
  assign new_n9249_ = ~new_n8779_ & ~\quotient[29] ;
  assign new_n9250_ = ~new_n8789_ & new_n8859_;
  assign new_n9251_ = ~new_n8855_ & new_n9250_;
  assign new_n9252_ = ~new_n8856_ & ~new_n8859_;
  assign new_n9253_ = ~new_n9251_ & ~new_n9252_;
  assign new_n9254_ = new_n9004_ & ~new_n9253_;
  assign new_n9255_ = ~new_n9001_ & new_n9254_;
  assign new_n9256_ = ~new_n9249_ & ~new_n9255_;
  assign new_n9257_ = ~\b[7]  & ~new_n9256_;
  assign new_n9258_ = ~new_n8788_ & ~\quotient[29] ;
  assign new_n9259_ = ~new_n8798_ & new_n8854_;
  assign new_n9260_ = ~new_n8850_ & new_n9259_;
  assign new_n9261_ = ~new_n8851_ & ~new_n8854_;
  assign new_n9262_ = ~new_n9260_ & ~new_n9261_;
  assign new_n9263_ = new_n9004_ & ~new_n9262_;
  assign new_n9264_ = ~new_n9001_ & new_n9263_;
  assign new_n9265_ = ~new_n9258_ & ~new_n9264_;
  assign new_n9266_ = ~\b[6]  & ~new_n9265_;
  assign new_n9267_ = ~new_n8797_ & ~\quotient[29] ;
  assign new_n9268_ = ~new_n8807_ & new_n8849_;
  assign new_n9269_ = ~new_n8845_ & new_n9268_;
  assign new_n9270_ = ~new_n8846_ & ~new_n8849_;
  assign new_n9271_ = ~new_n9269_ & ~new_n9270_;
  assign new_n9272_ = new_n9004_ & ~new_n9271_;
  assign new_n9273_ = ~new_n9001_ & new_n9272_;
  assign new_n9274_ = ~new_n9267_ & ~new_n9273_;
  assign new_n9275_ = ~\b[5]  & ~new_n9274_;
  assign new_n9276_ = ~new_n8806_ & ~\quotient[29] ;
  assign new_n9277_ = ~new_n8815_ & new_n8844_;
  assign new_n9278_ = ~new_n8840_ & new_n9277_;
  assign new_n9279_ = ~new_n8841_ & ~new_n8844_;
  assign new_n9280_ = ~new_n9278_ & ~new_n9279_;
  assign new_n9281_ = new_n9004_ & ~new_n9280_;
  assign new_n9282_ = ~new_n9001_ & new_n9281_;
  assign new_n9283_ = ~new_n9276_ & ~new_n9282_;
  assign new_n9284_ = ~\b[4]  & ~new_n9283_;
  assign new_n9285_ = ~new_n8814_ & ~\quotient[29] ;
  assign new_n9286_ = ~new_n8835_ & new_n8839_;
  assign new_n9287_ = ~new_n8834_ & new_n9286_;
  assign new_n9288_ = ~new_n8836_ & ~new_n8839_;
  assign new_n9289_ = ~new_n9287_ & ~new_n9288_;
  assign new_n9290_ = new_n9004_ & ~new_n9289_;
  assign new_n9291_ = ~new_n9001_ & new_n9290_;
  assign new_n9292_ = ~new_n9285_ & ~new_n9291_;
  assign new_n9293_ = ~\b[3]  & ~new_n9292_;
  assign new_n9294_ = ~new_n8828_ & ~\quotient[29] ;
  assign new_n9295_ = ~new_n8831_ & new_n8833_;
  assign new_n9296_ = ~new_n8829_ & new_n9295_;
  assign new_n9297_ = new_n9004_ & ~new_n9296_;
  assign new_n9298_ = ~new_n8834_ & new_n9297_;
  assign new_n9299_ = ~new_n9001_ & new_n9298_;
  assign new_n9300_ = ~new_n9294_ & ~new_n9299_;
  assign new_n9301_ = ~\b[2]  & ~new_n9300_;
  assign new_n9302_ = \b[0]  & ~\b[35] ;
  assign new_n9303_ = new_n294_ & new_n9302_;
  assign new_n9304_ = new_n340_ & new_n9303_;
  assign new_n9305_ = new_n338_ & new_n9304_;
  assign new_n9306_ = ~new_n9001_ & new_n9305_;
  assign new_n9307_ = \a[29]  & ~new_n9306_;
  assign new_n9308_ = new_n413_ & new_n8833_;
  assign new_n9309_ = new_n411_ & new_n9308_;
  assign new_n9310_ = new_n422_ & new_n9309_;
  assign new_n9311_ = new_n408_ & new_n9310_;
  assign new_n9312_ = ~new_n9001_ & new_n9311_;
  assign new_n9313_ = ~new_n9307_ & ~new_n9312_;
  assign new_n9314_ = \b[1]  & ~new_n9313_;
  assign new_n9315_ = ~\b[1]  & ~new_n9312_;
  assign new_n9316_ = ~new_n9307_ & new_n9315_;
  assign new_n9317_ = ~new_n9314_ & ~new_n9316_;
  assign new_n9318_ = ~\a[28]  & \b[0] ;
  assign new_n9319_ = ~new_n9317_ & ~new_n9318_;
  assign new_n9320_ = ~\b[1]  & ~new_n9313_;
  assign new_n9321_ = ~new_n9319_ & ~new_n9320_;
  assign new_n9322_ = \b[2]  & ~new_n9299_;
  assign new_n9323_ = ~new_n9294_ & new_n9322_;
  assign new_n9324_ = ~new_n9301_ & ~new_n9323_;
  assign new_n9325_ = ~new_n9321_ & new_n9324_;
  assign new_n9326_ = ~new_n9301_ & ~new_n9325_;
  assign new_n9327_ = \b[3]  & ~new_n9291_;
  assign new_n9328_ = ~new_n9285_ & new_n9327_;
  assign new_n9329_ = ~new_n9293_ & ~new_n9328_;
  assign new_n9330_ = ~new_n9326_ & new_n9329_;
  assign new_n9331_ = ~new_n9293_ & ~new_n9330_;
  assign new_n9332_ = \b[4]  & ~new_n9282_;
  assign new_n9333_ = ~new_n9276_ & new_n9332_;
  assign new_n9334_ = ~new_n9284_ & ~new_n9333_;
  assign new_n9335_ = ~new_n9331_ & new_n9334_;
  assign new_n9336_ = ~new_n9284_ & ~new_n9335_;
  assign new_n9337_ = \b[5]  & ~new_n9273_;
  assign new_n9338_ = ~new_n9267_ & new_n9337_;
  assign new_n9339_ = ~new_n9275_ & ~new_n9338_;
  assign new_n9340_ = ~new_n9336_ & new_n9339_;
  assign new_n9341_ = ~new_n9275_ & ~new_n9340_;
  assign new_n9342_ = \b[6]  & ~new_n9264_;
  assign new_n9343_ = ~new_n9258_ & new_n9342_;
  assign new_n9344_ = ~new_n9266_ & ~new_n9343_;
  assign new_n9345_ = ~new_n9341_ & new_n9344_;
  assign new_n9346_ = ~new_n9266_ & ~new_n9345_;
  assign new_n9347_ = \b[7]  & ~new_n9255_;
  assign new_n9348_ = ~new_n9249_ & new_n9347_;
  assign new_n9349_ = ~new_n9257_ & ~new_n9348_;
  assign new_n9350_ = ~new_n9346_ & new_n9349_;
  assign new_n9351_ = ~new_n9257_ & ~new_n9350_;
  assign new_n9352_ = \b[8]  & ~new_n9246_;
  assign new_n9353_ = ~new_n9240_ & new_n9352_;
  assign new_n9354_ = ~new_n9248_ & ~new_n9353_;
  assign new_n9355_ = ~new_n9351_ & new_n9354_;
  assign new_n9356_ = ~new_n9248_ & ~new_n9355_;
  assign new_n9357_ = \b[9]  & ~new_n9237_;
  assign new_n9358_ = ~new_n9231_ & new_n9357_;
  assign new_n9359_ = ~new_n9239_ & ~new_n9358_;
  assign new_n9360_ = ~new_n9356_ & new_n9359_;
  assign new_n9361_ = ~new_n9239_ & ~new_n9360_;
  assign new_n9362_ = \b[10]  & ~new_n9228_;
  assign new_n9363_ = ~new_n9222_ & new_n9362_;
  assign new_n9364_ = ~new_n9230_ & ~new_n9363_;
  assign new_n9365_ = ~new_n9361_ & new_n9364_;
  assign new_n9366_ = ~new_n9230_ & ~new_n9365_;
  assign new_n9367_ = \b[11]  & ~new_n9219_;
  assign new_n9368_ = ~new_n9213_ & new_n9367_;
  assign new_n9369_ = ~new_n9221_ & ~new_n9368_;
  assign new_n9370_ = ~new_n9366_ & new_n9369_;
  assign new_n9371_ = ~new_n9221_ & ~new_n9370_;
  assign new_n9372_ = \b[12]  & ~new_n9210_;
  assign new_n9373_ = ~new_n9204_ & new_n9372_;
  assign new_n9374_ = ~new_n9212_ & ~new_n9373_;
  assign new_n9375_ = ~new_n9371_ & new_n9374_;
  assign new_n9376_ = ~new_n9212_ & ~new_n9375_;
  assign new_n9377_ = \b[13]  & ~new_n9201_;
  assign new_n9378_ = ~new_n9195_ & new_n9377_;
  assign new_n9379_ = ~new_n9203_ & ~new_n9378_;
  assign new_n9380_ = ~new_n9376_ & new_n9379_;
  assign new_n9381_ = ~new_n9203_ & ~new_n9380_;
  assign new_n9382_ = \b[14]  & ~new_n9192_;
  assign new_n9383_ = ~new_n9186_ & new_n9382_;
  assign new_n9384_ = ~new_n9194_ & ~new_n9383_;
  assign new_n9385_ = ~new_n9381_ & new_n9384_;
  assign new_n9386_ = ~new_n9194_ & ~new_n9385_;
  assign new_n9387_ = \b[15]  & ~new_n9183_;
  assign new_n9388_ = ~new_n9177_ & new_n9387_;
  assign new_n9389_ = ~new_n9185_ & ~new_n9388_;
  assign new_n9390_ = ~new_n9386_ & new_n9389_;
  assign new_n9391_ = ~new_n9185_ & ~new_n9390_;
  assign new_n9392_ = \b[16]  & ~new_n9174_;
  assign new_n9393_ = ~new_n9168_ & new_n9392_;
  assign new_n9394_ = ~new_n9176_ & ~new_n9393_;
  assign new_n9395_ = ~new_n9391_ & new_n9394_;
  assign new_n9396_ = ~new_n9176_ & ~new_n9395_;
  assign new_n9397_ = \b[17]  & ~new_n9165_;
  assign new_n9398_ = ~new_n9159_ & new_n9397_;
  assign new_n9399_ = ~new_n9167_ & ~new_n9398_;
  assign new_n9400_ = ~new_n9396_ & new_n9399_;
  assign new_n9401_ = ~new_n9167_ & ~new_n9400_;
  assign new_n9402_ = \b[18]  & ~new_n9156_;
  assign new_n9403_ = ~new_n9150_ & new_n9402_;
  assign new_n9404_ = ~new_n9158_ & ~new_n9403_;
  assign new_n9405_ = ~new_n9401_ & new_n9404_;
  assign new_n9406_ = ~new_n9158_ & ~new_n9405_;
  assign new_n9407_ = \b[19]  & ~new_n9147_;
  assign new_n9408_ = ~new_n9141_ & new_n9407_;
  assign new_n9409_ = ~new_n9149_ & ~new_n9408_;
  assign new_n9410_ = ~new_n9406_ & new_n9409_;
  assign new_n9411_ = ~new_n9149_ & ~new_n9410_;
  assign new_n9412_ = \b[20]  & ~new_n9138_;
  assign new_n9413_ = ~new_n9132_ & new_n9412_;
  assign new_n9414_ = ~new_n9140_ & ~new_n9413_;
  assign new_n9415_ = ~new_n9411_ & new_n9414_;
  assign new_n9416_ = ~new_n9140_ & ~new_n9415_;
  assign new_n9417_ = \b[21]  & ~new_n9129_;
  assign new_n9418_ = ~new_n9123_ & new_n9417_;
  assign new_n9419_ = ~new_n9131_ & ~new_n9418_;
  assign new_n9420_ = ~new_n9416_ & new_n9419_;
  assign new_n9421_ = ~new_n9131_ & ~new_n9420_;
  assign new_n9422_ = \b[22]  & ~new_n9120_;
  assign new_n9423_ = ~new_n9114_ & new_n9422_;
  assign new_n9424_ = ~new_n9122_ & ~new_n9423_;
  assign new_n9425_ = ~new_n9421_ & new_n9424_;
  assign new_n9426_ = ~new_n9122_ & ~new_n9425_;
  assign new_n9427_ = \b[23]  & ~new_n9111_;
  assign new_n9428_ = ~new_n9105_ & new_n9427_;
  assign new_n9429_ = ~new_n9113_ & ~new_n9428_;
  assign new_n9430_ = ~new_n9426_ & new_n9429_;
  assign new_n9431_ = ~new_n9113_ & ~new_n9430_;
  assign new_n9432_ = \b[24]  & ~new_n9102_;
  assign new_n9433_ = ~new_n9096_ & new_n9432_;
  assign new_n9434_ = ~new_n9104_ & ~new_n9433_;
  assign new_n9435_ = ~new_n9431_ & new_n9434_;
  assign new_n9436_ = ~new_n9104_ & ~new_n9435_;
  assign new_n9437_ = \b[25]  & ~new_n9093_;
  assign new_n9438_ = ~new_n9087_ & new_n9437_;
  assign new_n9439_ = ~new_n9095_ & ~new_n9438_;
  assign new_n9440_ = ~new_n9436_ & new_n9439_;
  assign new_n9441_ = ~new_n9095_ & ~new_n9440_;
  assign new_n9442_ = \b[26]  & ~new_n9084_;
  assign new_n9443_ = ~new_n9078_ & new_n9442_;
  assign new_n9444_ = ~new_n9086_ & ~new_n9443_;
  assign new_n9445_ = ~new_n9441_ & new_n9444_;
  assign new_n9446_ = ~new_n9086_ & ~new_n9445_;
  assign new_n9447_ = \b[27]  & ~new_n9075_;
  assign new_n9448_ = ~new_n9069_ & new_n9447_;
  assign new_n9449_ = ~new_n9077_ & ~new_n9448_;
  assign new_n9450_ = ~new_n9446_ & new_n9449_;
  assign new_n9451_ = ~new_n9077_ & ~new_n9450_;
  assign new_n9452_ = \b[28]  & ~new_n9066_;
  assign new_n9453_ = ~new_n9060_ & new_n9452_;
  assign new_n9454_ = ~new_n9068_ & ~new_n9453_;
  assign new_n9455_ = ~new_n9451_ & new_n9454_;
  assign new_n9456_ = ~new_n9068_ & ~new_n9455_;
  assign new_n9457_ = \b[29]  & ~new_n9057_;
  assign new_n9458_ = ~new_n9051_ & new_n9457_;
  assign new_n9459_ = ~new_n9059_ & ~new_n9458_;
  assign new_n9460_ = ~new_n9456_ & new_n9459_;
  assign new_n9461_ = ~new_n9059_ & ~new_n9460_;
  assign new_n9462_ = \b[30]  & ~new_n9048_;
  assign new_n9463_ = ~new_n9042_ & new_n9462_;
  assign new_n9464_ = ~new_n9050_ & ~new_n9463_;
  assign new_n9465_ = ~new_n9461_ & new_n9464_;
  assign new_n9466_ = ~new_n9050_ & ~new_n9465_;
  assign new_n9467_ = \b[31]  & ~new_n9039_;
  assign new_n9468_ = ~new_n9033_ & new_n9467_;
  assign new_n9469_ = ~new_n9041_ & ~new_n9468_;
  assign new_n9470_ = ~new_n9466_ & new_n9469_;
  assign new_n9471_ = ~new_n9041_ & ~new_n9470_;
  assign new_n9472_ = \b[32]  & ~new_n9030_;
  assign new_n9473_ = ~new_n9024_ & new_n9472_;
  assign new_n9474_ = ~new_n9032_ & ~new_n9473_;
  assign new_n9475_ = ~new_n9471_ & new_n9474_;
  assign new_n9476_ = ~new_n9032_ & ~new_n9475_;
  assign new_n9477_ = \b[33]  & ~new_n9021_;
  assign new_n9478_ = ~new_n9015_ & new_n9477_;
  assign new_n9479_ = ~new_n9023_ & ~new_n9478_;
  assign new_n9480_ = ~new_n9476_ & new_n9479_;
  assign new_n9481_ = ~new_n9023_ & ~new_n9480_;
  assign new_n9482_ = \b[34]  & ~new_n9012_;
  assign new_n9483_ = ~new_n9006_ & new_n9482_;
  assign new_n9484_ = ~new_n9014_ & ~new_n9483_;
  assign new_n9485_ = ~new_n9481_ & new_n9484_;
  assign new_n9486_ = ~new_n9014_ & ~new_n9485_;
  assign new_n9487_ = ~new_n8535_ & ~\quotient[29] ;
  assign new_n9488_ = ~new_n8537_ & new_n8999_;
  assign new_n9489_ = ~new_n8995_ & new_n9488_;
  assign new_n9490_ = ~new_n8996_ & ~new_n8999_;
  assign new_n9491_ = ~new_n9489_ & ~new_n9490_;
  assign new_n9492_ = \quotient[29]  & ~new_n9491_;
  assign new_n9493_ = ~new_n9487_ & ~new_n9492_;
  assign new_n9494_ = ~\b[35]  & ~new_n9493_;
  assign new_n9495_ = \b[35]  & ~new_n9487_;
  assign new_n9496_ = ~new_n9492_ & new_n9495_;
  assign new_n9497_ = new_n512_ & ~new_n9496_;
  assign new_n9498_ = ~new_n9494_ & new_n9497_;
  assign new_n9499_ = ~new_n9486_ & new_n9498_;
  assign new_n9500_ = new_n9004_ & ~new_n9493_;
  assign \quotient[28]  = new_n9499_ | new_n9500_;
  assign new_n9502_ = ~new_n9023_ & new_n9484_;
  assign new_n9503_ = ~new_n9480_ & new_n9502_;
  assign new_n9504_ = ~new_n9481_ & ~new_n9484_;
  assign new_n9505_ = ~new_n9503_ & ~new_n9504_;
  assign new_n9506_ = \quotient[28]  & ~new_n9505_;
  assign new_n9507_ = ~new_n9013_ & ~new_n9500_;
  assign new_n9508_ = ~new_n9499_ & new_n9507_;
  assign new_n9509_ = ~new_n9506_ & ~new_n9508_;
  assign new_n9510_ = ~new_n9014_ & ~new_n9496_;
  assign new_n9511_ = ~new_n9494_ & new_n9510_;
  assign new_n9512_ = ~new_n9485_ & new_n9511_;
  assign new_n9513_ = ~new_n9494_ & ~new_n9496_;
  assign new_n9514_ = ~new_n9486_ & ~new_n9513_;
  assign new_n9515_ = ~new_n9512_ & ~new_n9514_;
  assign new_n9516_ = \quotient[28]  & ~new_n9515_;
  assign new_n9517_ = ~new_n9493_ & ~new_n9500_;
  assign new_n9518_ = ~new_n9499_ & new_n9517_;
  assign new_n9519_ = ~new_n9516_ & ~new_n9518_;
  assign new_n9520_ = ~\b[36]  & ~new_n9519_;
  assign new_n9521_ = ~\b[35]  & ~new_n9509_;
  assign new_n9522_ = ~new_n9032_ & new_n9479_;
  assign new_n9523_ = ~new_n9475_ & new_n9522_;
  assign new_n9524_ = ~new_n9476_ & ~new_n9479_;
  assign new_n9525_ = ~new_n9523_ & ~new_n9524_;
  assign new_n9526_ = \quotient[28]  & ~new_n9525_;
  assign new_n9527_ = ~new_n9022_ & ~new_n9500_;
  assign new_n9528_ = ~new_n9499_ & new_n9527_;
  assign new_n9529_ = ~new_n9526_ & ~new_n9528_;
  assign new_n9530_ = ~\b[34]  & ~new_n9529_;
  assign new_n9531_ = ~new_n9041_ & new_n9474_;
  assign new_n9532_ = ~new_n9470_ & new_n9531_;
  assign new_n9533_ = ~new_n9471_ & ~new_n9474_;
  assign new_n9534_ = ~new_n9532_ & ~new_n9533_;
  assign new_n9535_ = \quotient[28]  & ~new_n9534_;
  assign new_n9536_ = ~new_n9031_ & ~new_n9500_;
  assign new_n9537_ = ~new_n9499_ & new_n9536_;
  assign new_n9538_ = ~new_n9535_ & ~new_n9537_;
  assign new_n9539_ = ~\b[33]  & ~new_n9538_;
  assign new_n9540_ = ~new_n9050_ & new_n9469_;
  assign new_n9541_ = ~new_n9465_ & new_n9540_;
  assign new_n9542_ = ~new_n9466_ & ~new_n9469_;
  assign new_n9543_ = ~new_n9541_ & ~new_n9542_;
  assign new_n9544_ = \quotient[28]  & ~new_n9543_;
  assign new_n9545_ = ~new_n9040_ & ~new_n9500_;
  assign new_n9546_ = ~new_n9499_ & new_n9545_;
  assign new_n9547_ = ~new_n9544_ & ~new_n9546_;
  assign new_n9548_ = ~\b[32]  & ~new_n9547_;
  assign new_n9549_ = ~new_n9059_ & new_n9464_;
  assign new_n9550_ = ~new_n9460_ & new_n9549_;
  assign new_n9551_ = ~new_n9461_ & ~new_n9464_;
  assign new_n9552_ = ~new_n9550_ & ~new_n9551_;
  assign new_n9553_ = \quotient[28]  & ~new_n9552_;
  assign new_n9554_ = ~new_n9049_ & ~new_n9500_;
  assign new_n9555_ = ~new_n9499_ & new_n9554_;
  assign new_n9556_ = ~new_n9553_ & ~new_n9555_;
  assign new_n9557_ = ~\b[31]  & ~new_n9556_;
  assign new_n9558_ = ~new_n9068_ & new_n9459_;
  assign new_n9559_ = ~new_n9455_ & new_n9558_;
  assign new_n9560_ = ~new_n9456_ & ~new_n9459_;
  assign new_n9561_ = ~new_n9559_ & ~new_n9560_;
  assign new_n9562_ = \quotient[28]  & ~new_n9561_;
  assign new_n9563_ = ~new_n9058_ & ~new_n9500_;
  assign new_n9564_ = ~new_n9499_ & new_n9563_;
  assign new_n9565_ = ~new_n9562_ & ~new_n9564_;
  assign new_n9566_ = ~\b[30]  & ~new_n9565_;
  assign new_n9567_ = ~new_n9077_ & new_n9454_;
  assign new_n9568_ = ~new_n9450_ & new_n9567_;
  assign new_n9569_ = ~new_n9451_ & ~new_n9454_;
  assign new_n9570_ = ~new_n9568_ & ~new_n9569_;
  assign new_n9571_ = \quotient[28]  & ~new_n9570_;
  assign new_n9572_ = ~new_n9067_ & ~new_n9500_;
  assign new_n9573_ = ~new_n9499_ & new_n9572_;
  assign new_n9574_ = ~new_n9571_ & ~new_n9573_;
  assign new_n9575_ = ~\b[29]  & ~new_n9574_;
  assign new_n9576_ = ~new_n9086_ & new_n9449_;
  assign new_n9577_ = ~new_n9445_ & new_n9576_;
  assign new_n9578_ = ~new_n9446_ & ~new_n9449_;
  assign new_n9579_ = ~new_n9577_ & ~new_n9578_;
  assign new_n9580_ = \quotient[28]  & ~new_n9579_;
  assign new_n9581_ = ~new_n9076_ & ~new_n9500_;
  assign new_n9582_ = ~new_n9499_ & new_n9581_;
  assign new_n9583_ = ~new_n9580_ & ~new_n9582_;
  assign new_n9584_ = ~\b[28]  & ~new_n9583_;
  assign new_n9585_ = ~new_n9095_ & new_n9444_;
  assign new_n9586_ = ~new_n9440_ & new_n9585_;
  assign new_n9587_ = ~new_n9441_ & ~new_n9444_;
  assign new_n9588_ = ~new_n9586_ & ~new_n9587_;
  assign new_n9589_ = \quotient[28]  & ~new_n9588_;
  assign new_n9590_ = ~new_n9085_ & ~new_n9500_;
  assign new_n9591_ = ~new_n9499_ & new_n9590_;
  assign new_n9592_ = ~new_n9589_ & ~new_n9591_;
  assign new_n9593_ = ~\b[27]  & ~new_n9592_;
  assign new_n9594_ = ~new_n9104_ & new_n9439_;
  assign new_n9595_ = ~new_n9435_ & new_n9594_;
  assign new_n9596_ = ~new_n9436_ & ~new_n9439_;
  assign new_n9597_ = ~new_n9595_ & ~new_n9596_;
  assign new_n9598_ = \quotient[28]  & ~new_n9597_;
  assign new_n9599_ = ~new_n9094_ & ~new_n9500_;
  assign new_n9600_ = ~new_n9499_ & new_n9599_;
  assign new_n9601_ = ~new_n9598_ & ~new_n9600_;
  assign new_n9602_ = ~\b[26]  & ~new_n9601_;
  assign new_n9603_ = ~new_n9113_ & new_n9434_;
  assign new_n9604_ = ~new_n9430_ & new_n9603_;
  assign new_n9605_ = ~new_n9431_ & ~new_n9434_;
  assign new_n9606_ = ~new_n9604_ & ~new_n9605_;
  assign new_n9607_ = \quotient[28]  & ~new_n9606_;
  assign new_n9608_ = ~new_n9103_ & ~new_n9500_;
  assign new_n9609_ = ~new_n9499_ & new_n9608_;
  assign new_n9610_ = ~new_n9607_ & ~new_n9609_;
  assign new_n9611_ = ~\b[25]  & ~new_n9610_;
  assign new_n9612_ = ~new_n9122_ & new_n9429_;
  assign new_n9613_ = ~new_n9425_ & new_n9612_;
  assign new_n9614_ = ~new_n9426_ & ~new_n9429_;
  assign new_n9615_ = ~new_n9613_ & ~new_n9614_;
  assign new_n9616_ = \quotient[28]  & ~new_n9615_;
  assign new_n9617_ = ~new_n9112_ & ~new_n9500_;
  assign new_n9618_ = ~new_n9499_ & new_n9617_;
  assign new_n9619_ = ~new_n9616_ & ~new_n9618_;
  assign new_n9620_ = ~\b[24]  & ~new_n9619_;
  assign new_n9621_ = ~new_n9131_ & new_n9424_;
  assign new_n9622_ = ~new_n9420_ & new_n9621_;
  assign new_n9623_ = ~new_n9421_ & ~new_n9424_;
  assign new_n9624_ = ~new_n9622_ & ~new_n9623_;
  assign new_n9625_ = \quotient[28]  & ~new_n9624_;
  assign new_n9626_ = ~new_n9121_ & ~new_n9500_;
  assign new_n9627_ = ~new_n9499_ & new_n9626_;
  assign new_n9628_ = ~new_n9625_ & ~new_n9627_;
  assign new_n9629_ = ~\b[23]  & ~new_n9628_;
  assign new_n9630_ = ~new_n9140_ & new_n9419_;
  assign new_n9631_ = ~new_n9415_ & new_n9630_;
  assign new_n9632_ = ~new_n9416_ & ~new_n9419_;
  assign new_n9633_ = ~new_n9631_ & ~new_n9632_;
  assign new_n9634_ = \quotient[28]  & ~new_n9633_;
  assign new_n9635_ = ~new_n9130_ & ~new_n9500_;
  assign new_n9636_ = ~new_n9499_ & new_n9635_;
  assign new_n9637_ = ~new_n9634_ & ~new_n9636_;
  assign new_n9638_ = ~\b[22]  & ~new_n9637_;
  assign new_n9639_ = ~new_n9149_ & new_n9414_;
  assign new_n9640_ = ~new_n9410_ & new_n9639_;
  assign new_n9641_ = ~new_n9411_ & ~new_n9414_;
  assign new_n9642_ = ~new_n9640_ & ~new_n9641_;
  assign new_n9643_ = \quotient[28]  & ~new_n9642_;
  assign new_n9644_ = ~new_n9139_ & ~new_n9500_;
  assign new_n9645_ = ~new_n9499_ & new_n9644_;
  assign new_n9646_ = ~new_n9643_ & ~new_n9645_;
  assign new_n9647_ = ~\b[21]  & ~new_n9646_;
  assign new_n9648_ = ~new_n9158_ & new_n9409_;
  assign new_n9649_ = ~new_n9405_ & new_n9648_;
  assign new_n9650_ = ~new_n9406_ & ~new_n9409_;
  assign new_n9651_ = ~new_n9649_ & ~new_n9650_;
  assign new_n9652_ = \quotient[28]  & ~new_n9651_;
  assign new_n9653_ = ~new_n9148_ & ~new_n9500_;
  assign new_n9654_ = ~new_n9499_ & new_n9653_;
  assign new_n9655_ = ~new_n9652_ & ~new_n9654_;
  assign new_n9656_ = ~\b[20]  & ~new_n9655_;
  assign new_n9657_ = ~new_n9167_ & new_n9404_;
  assign new_n9658_ = ~new_n9400_ & new_n9657_;
  assign new_n9659_ = ~new_n9401_ & ~new_n9404_;
  assign new_n9660_ = ~new_n9658_ & ~new_n9659_;
  assign new_n9661_ = \quotient[28]  & ~new_n9660_;
  assign new_n9662_ = ~new_n9157_ & ~new_n9500_;
  assign new_n9663_ = ~new_n9499_ & new_n9662_;
  assign new_n9664_ = ~new_n9661_ & ~new_n9663_;
  assign new_n9665_ = ~\b[19]  & ~new_n9664_;
  assign new_n9666_ = ~new_n9176_ & new_n9399_;
  assign new_n9667_ = ~new_n9395_ & new_n9666_;
  assign new_n9668_ = ~new_n9396_ & ~new_n9399_;
  assign new_n9669_ = ~new_n9667_ & ~new_n9668_;
  assign new_n9670_ = \quotient[28]  & ~new_n9669_;
  assign new_n9671_ = ~new_n9166_ & ~new_n9500_;
  assign new_n9672_ = ~new_n9499_ & new_n9671_;
  assign new_n9673_ = ~new_n9670_ & ~new_n9672_;
  assign new_n9674_ = ~\b[18]  & ~new_n9673_;
  assign new_n9675_ = ~new_n9185_ & new_n9394_;
  assign new_n9676_ = ~new_n9390_ & new_n9675_;
  assign new_n9677_ = ~new_n9391_ & ~new_n9394_;
  assign new_n9678_ = ~new_n9676_ & ~new_n9677_;
  assign new_n9679_ = \quotient[28]  & ~new_n9678_;
  assign new_n9680_ = ~new_n9175_ & ~new_n9500_;
  assign new_n9681_ = ~new_n9499_ & new_n9680_;
  assign new_n9682_ = ~new_n9679_ & ~new_n9681_;
  assign new_n9683_ = ~\b[17]  & ~new_n9682_;
  assign new_n9684_ = ~new_n9194_ & new_n9389_;
  assign new_n9685_ = ~new_n9385_ & new_n9684_;
  assign new_n9686_ = ~new_n9386_ & ~new_n9389_;
  assign new_n9687_ = ~new_n9685_ & ~new_n9686_;
  assign new_n9688_ = \quotient[28]  & ~new_n9687_;
  assign new_n9689_ = ~new_n9184_ & ~new_n9500_;
  assign new_n9690_ = ~new_n9499_ & new_n9689_;
  assign new_n9691_ = ~new_n9688_ & ~new_n9690_;
  assign new_n9692_ = ~\b[16]  & ~new_n9691_;
  assign new_n9693_ = ~new_n9203_ & new_n9384_;
  assign new_n9694_ = ~new_n9380_ & new_n9693_;
  assign new_n9695_ = ~new_n9381_ & ~new_n9384_;
  assign new_n9696_ = ~new_n9694_ & ~new_n9695_;
  assign new_n9697_ = \quotient[28]  & ~new_n9696_;
  assign new_n9698_ = ~new_n9193_ & ~new_n9500_;
  assign new_n9699_ = ~new_n9499_ & new_n9698_;
  assign new_n9700_ = ~new_n9697_ & ~new_n9699_;
  assign new_n9701_ = ~\b[15]  & ~new_n9700_;
  assign new_n9702_ = ~new_n9212_ & new_n9379_;
  assign new_n9703_ = ~new_n9375_ & new_n9702_;
  assign new_n9704_ = ~new_n9376_ & ~new_n9379_;
  assign new_n9705_ = ~new_n9703_ & ~new_n9704_;
  assign new_n9706_ = \quotient[28]  & ~new_n9705_;
  assign new_n9707_ = ~new_n9202_ & ~new_n9500_;
  assign new_n9708_ = ~new_n9499_ & new_n9707_;
  assign new_n9709_ = ~new_n9706_ & ~new_n9708_;
  assign new_n9710_ = ~\b[14]  & ~new_n9709_;
  assign new_n9711_ = ~new_n9221_ & new_n9374_;
  assign new_n9712_ = ~new_n9370_ & new_n9711_;
  assign new_n9713_ = ~new_n9371_ & ~new_n9374_;
  assign new_n9714_ = ~new_n9712_ & ~new_n9713_;
  assign new_n9715_ = \quotient[28]  & ~new_n9714_;
  assign new_n9716_ = ~new_n9211_ & ~new_n9500_;
  assign new_n9717_ = ~new_n9499_ & new_n9716_;
  assign new_n9718_ = ~new_n9715_ & ~new_n9717_;
  assign new_n9719_ = ~\b[13]  & ~new_n9718_;
  assign new_n9720_ = ~new_n9230_ & new_n9369_;
  assign new_n9721_ = ~new_n9365_ & new_n9720_;
  assign new_n9722_ = ~new_n9366_ & ~new_n9369_;
  assign new_n9723_ = ~new_n9721_ & ~new_n9722_;
  assign new_n9724_ = \quotient[28]  & ~new_n9723_;
  assign new_n9725_ = ~new_n9220_ & ~new_n9500_;
  assign new_n9726_ = ~new_n9499_ & new_n9725_;
  assign new_n9727_ = ~new_n9724_ & ~new_n9726_;
  assign new_n9728_ = ~\b[12]  & ~new_n9727_;
  assign new_n9729_ = ~new_n9239_ & new_n9364_;
  assign new_n9730_ = ~new_n9360_ & new_n9729_;
  assign new_n9731_ = ~new_n9361_ & ~new_n9364_;
  assign new_n9732_ = ~new_n9730_ & ~new_n9731_;
  assign new_n9733_ = \quotient[28]  & ~new_n9732_;
  assign new_n9734_ = ~new_n9229_ & ~new_n9500_;
  assign new_n9735_ = ~new_n9499_ & new_n9734_;
  assign new_n9736_ = ~new_n9733_ & ~new_n9735_;
  assign new_n9737_ = ~\b[11]  & ~new_n9736_;
  assign new_n9738_ = ~new_n9248_ & new_n9359_;
  assign new_n9739_ = ~new_n9355_ & new_n9738_;
  assign new_n9740_ = ~new_n9356_ & ~new_n9359_;
  assign new_n9741_ = ~new_n9739_ & ~new_n9740_;
  assign new_n9742_ = \quotient[28]  & ~new_n9741_;
  assign new_n9743_ = ~new_n9238_ & ~new_n9500_;
  assign new_n9744_ = ~new_n9499_ & new_n9743_;
  assign new_n9745_ = ~new_n9742_ & ~new_n9744_;
  assign new_n9746_ = ~\b[10]  & ~new_n9745_;
  assign new_n9747_ = ~new_n9257_ & new_n9354_;
  assign new_n9748_ = ~new_n9350_ & new_n9747_;
  assign new_n9749_ = ~new_n9351_ & ~new_n9354_;
  assign new_n9750_ = ~new_n9748_ & ~new_n9749_;
  assign new_n9751_ = \quotient[28]  & ~new_n9750_;
  assign new_n9752_ = ~new_n9247_ & ~new_n9500_;
  assign new_n9753_ = ~new_n9499_ & new_n9752_;
  assign new_n9754_ = ~new_n9751_ & ~new_n9753_;
  assign new_n9755_ = ~\b[9]  & ~new_n9754_;
  assign new_n9756_ = ~new_n9266_ & new_n9349_;
  assign new_n9757_ = ~new_n9345_ & new_n9756_;
  assign new_n9758_ = ~new_n9346_ & ~new_n9349_;
  assign new_n9759_ = ~new_n9757_ & ~new_n9758_;
  assign new_n9760_ = \quotient[28]  & ~new_n9759_;
  assign new_n9761_ = ~new_n9256_ & ~new_n9500_;
  assign new_n9762_ = ~new_n9499_ & new_n9761_;
  assign new_n9763_ = ~new_n9760_ & ~new_n9762_;
  assign new_n9764_ = ~\b[8]  & ~new_n9763_;
  assign new_n9765_ = ~new_n9275_ & new_n9344_;
  assign new_n9766_ = ~new_n9340_ & new_n9765_;
  assign new_n9767_ = ~new_n9341_ & ~new_n9344_;
  assign new_n9768_ = ~new_n9766_ & ~new_n9767_;
  assign new_n9769_ = \quotient[28]  & ~new_n9768_;
  assign new_n9770_ = ~new_n9265_ & ~new_n9500_;
  assign new_n9771_ = ~new_n9499_ & new_n9770_;
  assign new_n9772_ = ~new_n9769_ & ~new_n9771_;
  assign new_n9773_ = ~\b[7]  & ~new_n9772_;
  assign new_n9774_ = ~new_n9284_ & new_n9339_;
  assign new_n9775_ = ~new_n9335_ & new_n9774_;
  assign new_n9776_ = ~new_n9336_ & ~new_n9339_;
  assign new_n9777_ = ~new_n9775_ & ~new_n9776_;
  assign new_n9778_ = \quotient[28]  & ~new_n9777_;
  assign new_n9779_ = ~new_n9274_ & ~new_n9500_;
  assign new_n9780_ = ~new_n9499_ & new_n9779_;
  assign new_n9781_ = ~new_n9778_ & ~new_n9780_;
  assign new_n9782_ = ~\b[6]  & ~new_n9781_;
  assign new_n9783_ = ~new_n9293_ & new_n9334_;
  assign new_n9784_ = ~new_n9330_ & new_n9783_;
  assign new_n9785_ = ~new_n9331_ & ~new_n9334_;
  assign new_n9786_ = ~new_n9784_ & ~new_n9785_;
  assign new_n9787_ = \quotient[28]  & ~new_n9786_;
  assign new_n9788_ = ~new_n9283_ & ~new_n9500_;
  assign new_n9789_ = ~new_n9499_ & new_n9788_;
  assign new_n9790_ = ~new_n9787_ & ~new_n9789_;
  assign new_n9791_ = ~\b[5]  & ~new_n9790_;
  assign new_n9792_ = ~new_n9301_ & new_n9329_;
  assign new_n9793_ = ~new_n9325_ & new_n9792_;
  assign new_n9794_ = ~new_n9326_ & ~new_n9329_;
  assign new_n9795_ = ~new_n9793_ & ~new_n9794_;
  assign new_n9796_ = \quotient[28]  & ~new_n9795_;
  assign new_n9797_ = ~new_n9292_ & ~new_n9500_;
  assign new_n9798_ = ~new_n9499_ & new_n9797_;
  assign new_n9799_ = ~new_n9796_ & ~new_n9798_;
  assign new_n9800_ = ~\b[4]  & ~new_n9799_;
  assign new_n9801_ = ~new_n9320_ & new_n9324_;
  assign new_n9802_ = ~new_n9319_ & new_n9801_;
  assign new_n9803_ = ~new_n9321_ & ~new_n9324_;
  assign new_n9804_ = ~new_n9802_ & ~new_n9803_;
  assign new_n9805_ = \quotient[28]  & ~new_n9804_;
  assign new_n9806_ = ~new_n9300_ & ~new_n9500_;
  assign new_n9807_ = ~new_n9499_ & new_n9806_;
  assign new_n9808_ = ~new_n9805_ & ~new_n9807_;
  assign new_n9809_ = ~\b[3]  & ~new_n9808_;
  assign new_n9810_ = ~new_n9316_ & new_n9318_;
  assign new_n9811_ = ~new_n9314_ & new_n9810_;
  assign new_n9812_ = ~new_n9319_ & ~new_n9811_;
  assign new_n9813_ = \quotient[28]  & new_n9812_;
  assign new_n9814_ = ~new_n9313_ & ~new_n9500_;
  assign new_n9815_ = ~new_n9499_ & new_n9814_;
  assign new_n9816_ = ~new_n9813_ & ~new_n9815_;
  assign new_n9817_ = ~\b[2]  & ~new_n9816_;
  assign new_n9818_ = \b[0]  & \quotient[28] ;
  assign new_n9819_ = \a[28]  & ~new_n9818_;
  assign new_n9820_ = new_n9318_ & \quotient[28] ;
  assign new_n9821_ = ~new_n9819_ & ~new_n9820_;
  assign new_n9822_ = \b[1]  & ~new_n9821_;
  assign new_n9823_ = ~\b[1]  & ~new_n9820_;
  assign new_n9824_ = ~new_n9819_ & new_n9823_;
  assign new_n9825_ = ~new_n9822_ & ~new_n9824_;
  assign new_n9826_ = ~\a[27]  & \b[0] ;
  assign new_n9827_ = ~new_n9825_ & ~new_n9826_;
  assign new_n9828_ = ~\b[1]  & ~new_n9821_;
  assign new_n9829_ = ~new_n9827_ & ~new_n9828_;
  assign new_n9830_ = \b[2]  & ~new_n9815_;
  assign new_n9831_ = ~new_n9813_ & new_n9830_;
  assign new_n9832_ = ~new_n9817_ & ~new_n9831_;
  assign new_n9833_ = ~new_n9829_ & new_n9832_;
  assign new_n9834_ = ~new_n9817_ & ~new_n9833_;
  assign new_n9835_ = \b[3]  & ~new_n9807_;
  assign new_n9836_ = ~new_n9805_ & new_n9835_;
  assign new_n9837_ = ~new_n9809_ & ~new_n9836_;
  assign new_n9838_ = ~new_n9834_ & new_n9837_;
  assign new_n9839_ = ~new_n9809_ & ~new_n9838_;
  assign new_n9840_ = \b[4]  & ~new_n9798_;
  assign new_n9841_ = ~new_n9796_ & new_n9840_;
  assign new_n9842_ = ~new_n9800_ & ~new_n9841_;
  assign new_n9843_ = ~new_n9839_ & new_n9842_;
  assign new_n9844_ = ~new_n9800_ & ~new_n9843_;
  assign new_n9845_ = \b[5]  & ~new_n9789_;
  assign new_n9846_ = ~new_n9787_ & new_n9845_;
  assign new_n9847_ = ~new_n9791_ & ~new_n9846_;
  assign new_n9848_ = ~new_n9844_ & new_n9847_;
  assign new_n9849_ = ~new_n9791_ & ~new_n9848_;
  assign new_n9850_ = \b[6]  & ~new_n9780_;
  assign new_n9851_ = ~new_n9778_ & new_n9850_;
  assign new_n9852_ = ~new_n9782_ & ~new_n9851_;
  assign new_n9853_ = ~new_n9849_ & new_n9852_;
  assign new_n9854_ = ~new_n9782_ & ~new_n9853_;
  assign new_n9855_ = \b[7]  & ~new_n9771_;
  assign new_n9856_ = ~new_n9769_ & new_n9855_;
  assign new_n9857_ = ~new_n9773_ & ~new_n9856_;
  assign new_n9858_ = ~new_n9854_ & new_n9857_;
  assign new_n9859_ = ~new_n9773_ & ~new_n9858_;
  assign new_n9860_ = \b[8]  & ~new_n9762_;
  assign new_n9861_ = ~new_n9760_ & new_n9860_;
  assign new_n9862_ = ~new_n9764_ & ~new_n9861_;
  assign new_n9863_ = ~new_n9859_ & new_n9862_;
  assign new_n9864_ = ~new_n9764_ & ~new_n9863_;
  assign new_n9865_ = \b[9]  & ~new_n9753_;
  assign new_n9866_ = ~new_n9751_ & new_n9865_;
  assign new_n9867_ = ~new_n9755_ & ~new_n9866_;
  assign new_n9868_ = ~new_n9864_ & new_n9867_;
  assign new_n9869_ = ~new_n9755_ & ~new_n9868_;
  assign new_n9870_ = \b[10]  & ~new_n9744_;
  assign new_n9871_ = ~new_n9742_ & new_n9870_;
  assign new_n9872_ = ~new_n9746_ & ~new_n9871_;
  assign new_n9873_ = ~new_n9869_ & new_n9872_;
  assign new_n9874_ = ~new_n9746_ & ~new_n9873_;
  assign new_n9875_ = \b[11]  & ~new_n9735_;
  assign new_n9876_ = ~new_n9733_ & new_n9875_;
  assign new_n9877_ = ~new_n9737_ & ~new_n9876_;
  assign new_n9878_ = ~new_n9874_ & new_n9877_;
  assign new_n9879_ = ~new_n9737_ & ~new_n9878_;
  assign new_n9880_ = \b[12]  & ~new_n9726_;
  assign new_n9881_ = ~new_n9724_ & new_n9880_;
  assign new_n9882_ = ~new_n9728_ & ~new_n9881_;
  assign new_n9883_ = ~new_n9879_ & new_n9882_;
  assign new_n9884_ = ~new_n9728_ & ~new_n9883_;
  assign new_n9885_ = \b[13]  & ~new_n9717_;
  assign new_n9886_ = ~new_n9715_ & new_n9885_;
  assign new_n9887_ = ~new_n9719_ & ~new_n9886_;
  assign new_n9888_ = ~new_n9884_ & new_n9887_;
  assign new_n9889_ = ~new_n9719_ & ~new_n9888_;
  assign new_n9890_ = \b[14]  & ~new_n9708_;
  assign new_n9891_ = ~new_n9706_ & new_n9890_;
  assign new_n9892_ = ~new_n9710_ & ~new_n9891_;
  assign new_n9893_ = ~new_n9889_ & new_n9892_;
  assign new_n9894_ = ~new_n9710_ & ~new_n9893_;
  assign new_n9895_ = \b[15]  & ~new_n9699_;
  assign new_n9896_ = ~new_n9697_ & new_n9895_;
  assign new_n9897_ = ~new_n9701_ & ~new_n9896_;
  assign new_n9898_ = ~new_n9894_ & new_n9897_;
  assign new_n9899_ = ~new_n9701_ & ~new_n9898_;
  assign new_n9900_ = \b[16]  & ~new_n9690_;
  assign new_n9901_ = ~new_n9688_ & new_n9900_;
  assign new_n9902_ = ~new_n9692_ & ~new_n9901_;
  assign new_n9903_ = ~new_n9899_ & new_n9902_;
  assign new_n9904_ = ~new_n9692_ & ~new_n9903_;
  assign new_n9905_ = \b[17]  & ~new_n9681_;
  assign new_n9906_ = ~new_n9679_ & new_n9905_;
  assign new_n9907_ = ~new_n9683_ & ~new_n9906_;
  assign new_n9908_ = ~new_n9904_ & new_n9907_;
  assign new_n9909_ = ~new_n9683_ & ~new_n9908_;
  assign new_n9910_ = \b[18]  & ~new_n9672_;
  assign new_n9911_ = ~new_n9670_ & new_n9910_;
  assign new_n9912_ = ~new_n9674_ & ~new_n9911_;
  assign new_n9913_ = ~new_n9909_ & new_n9912_;
  assign new_n9914_ = ~new_n9674_ & ~new_n9913_;
  assign new_n9915_ = \b[19]  & ~new_n9663_;
  assign new_n9916_ = ~new_n9661_ & new_n9915_;
  assign new_n9917_ = ~new_n9665_ & ~new_n9916_;
  assign new_n9918_ = ~new_n9914_ & new_n9917_;
  assign new_n9919_ = ~new_n9665_ & ~new_n9918_;
  assign new_n9920_ = \b[20]  & ~new_n9654_;
  assign new_n9921_ = ~new_n9652_ & new_n9920_;
  assign new_n9922_ = ~new_n9656_ & ~new_n9921_;
  assign new_n9923_ = ~new_n9919_ & new_n9922_;
  assign new_n9924_ = ~new_n9656_ & ~new_n9923_;
  assign new_n9925_ = \b[21]  & ~new_n9645_;
  assign new_n9926_ = ~new_n9643_ & new_n9925_;
  assign new_n9927_ = ~new_n9647_ & ~new_n9926_;
  assign new_n9928_ = ~new_n9924_ & new_n9927_;
  assign new_n9929_ = ~new_n9647_ & ~new_n9928_;
  assign new_n9930_ = \b[22]  & ~new_n9636_;
  assign new_n9931_ = ~new_n9634_ & new_n9930_;
  assign new_n9932_ = ~new_n9638_ & ~new_n9931_;
  assign new_n9933_ = ~new_n9929_ & new_n9932_;
  assign new_n9934_ = ~new_n9638_ & ~new_n9933_;
  assign new_n9935_ = \b[23]  & ~new_n9627_;
  assign new_n9936_ = ~new_n9625_ & new_n9935_;
  assign new_n9937_ = ~new_n9629_ & ~new_n9936_;
  assign new_n9938_ = ~new_n9934_ & new_n9937_;
  assign new_n9939_ = ~new_n9629_ & ~new_n9938_;
  assign new_n9940_ = \b[24]  & ~new_n9618_;
  assign new_n9941_ = ~new_n9616_ & new_n9940_;
  assign new_n9942_ = ~new_n9620_ & ~new_n9941_;
  assign new_n9943_ = ~new_n9939_ & new_n9942_;
  assign new_n9944_ = ~new_n9620_ & ~new_n9943_;
  assign new_n9945_ = \b[25]  & ~new_n9609_;
  assign new_n9946_ = ~new_n9607_ & new_n9945_;
  assign new_n9947_ = ~new_n9611_ & ~new_n9946_;
  assign new_n9948_ = ~new_n9944_ & new_n9947_;
  assign new_n9949_ = ~new_n9611_ & ~new_n9948_;
  assign new_n9950_ = \b[26]  & ~new_n9600_;
  assign new_n9951_ = ~new_n9598_ & new_n9950_;
  assign new_n9952_ = ~new_n9602_ & ~new_n9951_;
  assign new_n9953_ = ~new_n9949_ & new_n9952_;
  assign new_n9954_ = ~new_n9602_ & ~new_n9953_;
  assign new_n9955_ = \b[27]  & ~new_n9591_;
  assign new_n9956_ = ~new_n9589_ & new_n9955_;
  assign new_n9957_ = ~new_n9593_ & ~new_n9956_;
  assign new_n9958_ = ~new_n9954_ & new_n9957_;
  assign new_n9959_ = ~new_n9593_ & ~new_n9958_;
  assign new_n9960_ = \b[28]  & ~new_n9582_;
  assign new_n9961_ = ~new_n9580_ & new_n9960_;
  assign new_n9962_ = ~new_n9584_ & ~new_n9961_;
  assign new_n9963_ = ~new_n9959_ & new_n9962_;
  assign new_n9964_ = ~new_n9584_ & ~new_n9963_;
  assign new_n9965_ = \b[29]  & ~new_n9573_;
  assign new_n9966_ = ~new_n9571_ & new_n9965_;
  assign new_n9967_ = ~new_n9575_ & ~new_n9966_;
  assign new_n9968_ = ~new_n9964_ & new_n9967_;
  assign new_n9969_ = ~new_n9575_ & ~new_n9968_;
  assign new_n9970_ = \b[30]  & ~new_n9564_;
  assign new_n9971_ = ~new_n9562_ & new_n9970_;
  assign new_n9972_ = ~new_n9566_ & ~new_n9971_;
  assign new_n9973_ = ~new_n9969_ & new_n9972_;
  assign new_n9974_ = ~new_n9566_ & ~new_n9973_;
  assign new_n9975_ = \b[31]  & ~new_n9555_;
  assign new_n9976_ = ~new_n9553_ & new_n9975_;
  assign new_n9977_ = ~new_n9557_ & ~new_n9976_;
  assign new_n9978_ = ~new_n9974_ & new_n9977_;
  assign new_n9979_ = ~new_n9557_ & ~new_n9978_;
  assign new_n9980_ = \b[32]  & ~new_n9546_;
  assign new_n9981_ = ~new_n9544_ & new_n9980_;
  assign new_n9982_ = ~new_n9548_ & ~new_n9981_;
  assign new_n9983_ = ~new_n9979_ & new_n9982_;
  assign new_n9984_ = ~new_n9548_ & ~new_n9983_;
  assign new_n9985_ = \b[33]  & ~new_n9537_;
  assign new_n9986_ = ~new_n9535_ & new_n9985_;
  assign new_n9987_ = ~new_n9539_ & ~new_n9986_;
  assign new_n9988_ = ~new_n9984_ & new_n9987_;
  assign new_n9989_ = ~new_n9539_ & ~new_n9988_;
  assign new_n9990_ = \b[34]  & ~new_n9528_;
  assign new_n9991_ = ~new_n9526_ & new_n9990_;
  assign new_n9992_ = ~new_n9530_ & ~new_n9991_;
  assign new_n9993_ = ~new_n9989_ & new_n9992_;
  assign new_n9994_ = ~new_n9530_ & ~new_n9993_;
  assign new_n9995_ = \b[35]  & ~new_n9508_;
  assign new_n9996_ = ~new_n9506_ & new_n9995_;
  assign new_n9997_ = ~new_n9521_ & ~new_n9996_;
  assign new_n9998_ = ~new_n9994_ & new_n9997_;
  assign new_n9999_ = ~new_n9521_ & ~new_n9998_;
  assign new_n10000_ = \b[36]  & ~new_n9518_;
  assign new_n10001_ = ~new_n9516_ & new_n10000_;
  assign new_n10002_ = ~new_n9520_ & ~new_n10001_;
  assign new_n10003_ = ~new_n9999_ & new_n10002_;
  assign new_n10004_ = ~new_n9520_ & ~new_n10003_;
  assign \quotient[27]  = new_n599_ & ~new_n10004_;
  assign new_n10006_ = ~new_n9509_ & ~\quotient[27] ;
  assign new_n10007_ = ~new_n9530_ & new_n9997_;
  assign new_n10008_ = ~new_n9993_ & new_n10007_;
  assign new_n10009_ = ~new_n9994_ & ~new_n9997_;
  assign new_n10010_ = ~new_n10008_ & ~new_n10009_;
  assign new_n10011_ = new_n599_ & ~new_n10010_;
  assign new_n10012_ = ~new_n10004_ & new_n10011_;
  assign new_n10013_ = ~new_n10006_ & ~new_n10012_;
  assign new_n10014_ = ~new_n9519_ & ~\quotient[27] ;
  assign new_n10015_ = ~new_n9521_ & new_n10002_;
  assign new_n10016_ = ~new_n9998_ & new_n10015_;
  assign new_n10017_ = ~new_n9999_ & ~new_n10002_;
  assign new_n10018_ = ~new_n10016_ & ~new_n10017_;
  assign new_n10019_ = \quotient[27]  & ~new_n10018_;
  assign new_n10020_ = ~new_n10014_ & ~new_n10019_;
  assign new_n10021_ = ~\b[37]  & ~new_n10020_;
  assign new_n10022_ = ~\b[36]  & ~new_n10013_;
  assign new_n10023_ = ~new_n9529_ & ~\quotient[27] ;
  assign new_n10024_ = ~new_n9539_ & new_n9992_;
  assign new_n10025_ = ~new_n9988_ & new_n10024_;
  assign new_n10026_ = ~new_n9989_ & ~new_n9992_;
  assign new_n10027_ = ~new_n10025_ & ~new_n10026_;
  assign new_n10028_ = new_n599_ & ~new_n10027_;
  assign new_n10029_ = ~new_n10004_ & new_n10028_;
  assign new_n10030_ = ~new_n10023_ & ~new_n10029_;
  assign new_n10031_ = ~\b[35]  & ~new_n10030_;
  assign new_n10032_ = ~new_n9538_ & ~\quotient[27] ;
  assign new_n10033_ = ~new_n9548_ & new_n9987_;
  assign new_n10034_ = ~new_n9983_ & new_n10033_;
  assign new_n10035_ = ~new_n9984_ & ~new_n9987_;
  assign new_n10036_ = ~new_n10034_ & ~new_n10035_;
  assign new_n10037_ = new_n599_ & ~new_n10036_;
  assign new_n10038_ = ~new_n10004_ & new_n10037_;
  assign new_n10039_ = ~new_n10032_ & ~new_n10038_;
  assign new_n10040_ = ~\b[34]  & ~new_n10039_;
  assign new_n10041_ = ~new_n9547_ & ~\quotient[27] ;
  assign new_n10042_ = ~new_n9557_ & new_n9982_;
  assign new_n10043_ = ~new_n9978_ & new_n10042_;
  assign new_n10044_ = ~new_n9979_ & ~new_n9982_;
  assign new_n10045_ = ~new_n10043_ & ~new_n10044_;
  assign new_n10046_ = new_n599_ & ~new_n10045_;
  assign new_n10047_ = ~new_n10004_ & new_n10046_;
  assign new_n10048_ = ~new_n10041_ & ~new_n10047_;
  assign new_n10049_ = ~\b[33]  & ~new_n10048_;
  assign new_n10050_ = ~new_n9556_ & ~\quotient[27] ;
  assign new_n10051_ = ~new_n9566_ & new_n9977_;
  assign new_n10052_ = ~new_n9973_ & new_n10051_;
  assign new_n10053_ = ~new_n9974_ & ~new_n9977_;
  assign new_n10054_ = ~new_n10052_ & ~new_n10053_;
  assign new_n10055_ = new_n599_ & ~new_n10054_;
  assign new_n10056_ = ~new_n10004_ & new_n10055_;
  assign new_n10057_ = ~new_n10050_ & ~new_n10056_;
  assign new_n10058_ = ~\b[32]  & ~new_n10057_;
  assign new_n10059_ = ~new_n9565_ & ~\quotient[27] ;
  assign new_n10060_ = ~new_n9575_ & new_n9972_;
  assign new_n10061_ = ~new_n9968_ & new_n10060_;
  assign new_n10062_ = ~new_n9969_ & ~new_n9972_;
  assign new_n10063_ = ~new_n10061_ & ~new_n10062_;
  assign new_n10064_ = new_n599_ & ~new_n10063_;
  assign new_n10065_ = ~new_n10004_ & new_n10064_;
  assign new_n10066_ = ~new_n10059_ & ~new_n10065_;
  assign new_n10067_ = ~\b[31]  & ~new_n10066_;
  assign new_n10068_ = ~new_n9574_ & ~\quotient[27] ;
  assign new_n10069_ = ~new_n9584_ & new_n9967_;
  assign new_n10070_ = ~new_n9963_ & new_n10069_;
  assign new_n10071_ = ~new_n9964_ & ~new_n9967_;
  assign new_n10072_ = ~new_n10070_ & ~new_n10071_;
  assign new_n10073_ = new_n599_ & ~new_n10072_;
  assign new_n10074_ = ~new_n10004_ & new_n10073_;
  assign new_n10075_ = ~new_n10068_ & ~new_n10074_;
  assign new_n10076_ = ~\b[30]  & ~new_n10075_;
  assign new_n10077_ = ~new_n9583_ & ~\quotient[27] ;
  assign new_n10078_ = ~new_n9593_ & new_n9962_;
  assign new_n10079_ = ~new_n9958_ & new_n10078_;
  assign new_n10080_ = ~new_n9959_ & ~new_n9962_;
  assign new_n10081_ = ~new_n10079_ & ~new_n10080_;
  assign new_n10082_ = new_n599_ & ~new_n10081_;
  assign new_n10083_ = ~new_n10004_ & new_n10082_;
  assign new_n10084_ = ~new_n10077_ & ~new_n10083_;
  assign new_n10085_ = ~\b[29]  & ~new_n10084_;
  assign new_n10086_ = ~new_n9592_ & ~\quotient[27] ;
  assign new_n10087_ = ~new_n9602_ & new_n9957_;
  assign new_n10088_ = ~new_n9953_ & new_n10087_;
  assign new_n10089_ = ~new_n9954_ & ~new_n9957_;
  assign new_n10090_ = ~new_n10088_ & ~new_n10089_;
  assign new_n10091_ = new_n599_ & ~new_n10090_;
  assign new_n10092_ = ~new_n10004_ & new_n10091_;
  assign new_n10093_ = ~new_n10086_ & ~new_n10092_;
  assign new_n10094_ = ~\b[28]  & ~new_n10093_;
  assign new_n10095_ = ~new_n9601_ & ~\quotient[27] ;
  assign new_n10096_ = ~new_n9611_ & new_n9952_;
  assign new_n10097_ = ~new_n9948_ & new_n10096_;
  assign new_n10098_ = ~new_n9949_ & ~new_n9952_;
  assign new_n10099_ = ~new_n10097_ & ~new_n10098_;
  assign new_n10100_ = new_n599_ & ~new_n10099_;
  assign new_n10101_ = ~new_n10004_ & new_n10100_;
  assign new_n10102_ = ~new_n10095_ & ~new_n10101_;
  assign new_n10103_ = ~\b[27]  & ~new_n10102_;
  assign new_n10104_ = ~new_n9610_ & ~\quotient[27] ;
  assign new_n10105_ = ~new_n9620_ & new_n9947_;
  assign new_n10106_ = ~new_n9943_ & new_n10105_;
  assign new_n10107_ = ~new_n9944_ & ~new_n9947_;
  assign new_n10108_ = ~new_n10106_ & ~new_n10107_;
  assign new_n10109_ = new_n599_ & ~new_n10108_;
  assign new_n10110_ = ~new_n10004_ & new_n10109_;
  assign new_n10111_ = ~new_n10104_ & ~new_n10110_;
  assign new_n10112_ = ~\b[26]  & ~new_n10111_;
  assign new_n10113_ = ~new_n9619_ & ~\quotient[27] ;
  assign new_n10114_ = ~new_n9629_ & new_n9942_;
  assign new_n10115_ = ~new_n9938_ & new_n10114_;
  assign new_n10116_ = ~new_n9939_ & ~new_n9942_;
  assign new_n10117_ = ~new_n10115_ & ~new_n10116_;
  assign new_n10118_ = new_n599_ & ~new_n10117_;
  assign new_n10119_ = ~new_n10004_ & new_n10118_;
  assign new_n10120_ = ~new_n10113_ & ~new_n10119_;
  assign new_n10121_ = ~\b[25]  & ~new_n10120_;
  assign new_n10122_ = ~new_n9628_ & ~\quotient[27] ;
  assign new_n10123_ = ~new_n9638_ & new_n9937_;
  assign new_n10124_ = ~new_n9933_ & new_n10123_;
  assign new_n10125_ = ~new_n9934_ & ~new_n9937_;
  assign new_n10126_ = ~new_n10124_ & ~new_n10125_;
  assign new_n10127_ = new_n599_ & ~new_n10126_;
  assign new_n10128_ = ~new_n10004_ & new_n10127_;
  assign new_n10129_ = ~new_n10122_ & ~new_n10128_;
  assign new_n10130_ = ~\b[24]  & ~new_n10129_;
  assign new_n10131_ = ~new_n9637_ & ~\quotient[27] ;
  assign new_n10132_ = ~new_n9647_ & new_n9932_;
  assign new_n10133_ = ~new_n9928_ & new_n10132_;
  assign new_n10134_ = ~new_n9929_ & ~new_n9932_;
  assign new_n10135_ = ~new_n10133_ & ~new_n10134_;
  assign new_n10136_ = new_n599_ & ~new_n10135_;
  assign new_n10137_ = ~new_n10004_ & new_n10136_;
  assign new_n10138_ = ~new_n10131_ & ~new_n10137_;
  assign new_n10139_ = ~\b[23]  & ~new_n10138_;
  assign new_n10140_ = ~new_n9646_ & ~\quotient[27] ;
  assign new_n10141_ = ~new_n9656_ & new_n9927_;
  assign new_n10142_ = ~new_n9923_ & new_n10141_;
  assign new_n10143_ = ~new_n9924_ & ~new_n9927_;
  assign new_n10144_ = ~new_n10142_ & ~new_n10143_;
  assign new_n10145_ = new_n599_ & ~new_n10144_;
  assign new_n10146_ = ~new_n10004_ & new_n10145_;
  assign new_n10147_ = ~new_n10140_ & ~new_n10146_;
  assign new_n10148_ = ~\b[22]  & ~new_n10147_;
  assign new_n10149_ = ~new_n9655_ & ~\quotient[27] ;
  assign new_n10150_ = ~new_n9665_ & new_n9922_;
  assign new_n10151_ = ~new_n9918_ & new_n10150_;
  assign new_n10152_ = ~new_n9919_ & ~new_n9922_;
  assign new_n10153_ = ~new_n10151_ & ~new_n10152_;
  assign new_n10154_ = new_n599_ & ~new_n10153_;
  assign new_n10155_ = ~new_n10004_ & new_n10154_;
  assign new_n10156_ = ~new_n10149_ & ~new_n10155_;
  assign new_n10157_ = ~\b[21]  & ~new_n10156_;
  assign new_n10158_ = ~new_n9664_ & ~\quotient[27] ;
  assign new_n10159_ = ~new_n9674_ & new_n9917_;
  assign new_n10160_ = ~new_n9913_ & new_n10159_;
  assign new_n10161_ = ~new_n9914_ & ~new_n9917_;
  assign new_n10162_ = ~new_n10160_ & ~new_n10161_;
  assign new_n10163_ = new_n599_ & ~new_n10162_;
  assign new_n10164_ = ~new_n10004_ & new_n10163_;
  assign new_n10165_ = ~new_n10158_ & ~new_n10164_;
  assign new_n10166_ = ~\b[20]  & ~new_n10165_;
  assign new_n10167_ = ~new_n9673_ & ~\quotient[27] ;
  assign new_n10168_ = ~new_n9683_ & new_n9912_;
  assign new_n10169_ = ~new_n9908_ & new_n10168_;
  assign new_n10170_ = ~new_n9909_ & ~new_n9912_;
  assign new_n10171_ = ~new_n10169_ & ~new_n10170_;
  assign new_n10172_ = new_n599_ & ~new_n10171_;
  assign new_n10173_ = ~new_n10004_ & new_n10172_;
  assign new_n10174_ = ~new_n10167_ & ~new_n10173_;
  assign new_n10175_ = ~\b[19]  & ~new_n10174_;
  assign new_n10176_ = ~new_n9682_ & ~\quotient[27] ;
  assign new_n10177_ = ~new_n9692_ & new_n9907_;
  assign new_n10178_ = ~new_n9903_ & new_n10177_;
  assign new_n10179_ = ~new_n9904_ & ~new_n9907_;
  assign new_n10180_ = ~new_n10178_ & ~new_n10179_;
  assign new_n10181_ = new_n599_ & ~new_n10180_;
  assign new_n10182_ = ~new_n10004_ & new_n10181_;
  assign new_n10183_ = ~new_n10176_ & ~new_n10182_;
  assign new_n10184_ = ~\b[18]  & ~new_n10183_;
  assign new_n10185_ = ~new_n9691_ & ~\quotient[27] ;
  assign new_n10186_ = ~new_n9701_ & new_n9902_;
  assign new_n10187_ = ~new_n9898_ & new_n10186_;
  assign new_n10188_ = ~new_n9899_ & ~new_n9902_;
  assign new_n10189_ = ~new_n10187_ & ~new_n10188_;
  assign new_n10190_ = new_n599_ & ~new_n10189_;
  assign new_n10191_ = ~new_n10004_ & new_n10190_;
  assign new_n10192_ = ~new_n10185_ & ~new_n10191_;
  assign new_n10193_ = ~\b[17]  & ~new_n10192_;
  assign new_n10194_ = ~new_n9700_ & ~\quotient[27] ;
  assign new_n10195_ = ~new_n9710_ & new_n9897_;
  assign new_n10196_ = ~new_n9893_ & new_n10195_;
  assign new_n10197_ = ~new_n9894_ & ~new_n9897_;
  assign new_n10198_ = ~new_n10196_ & ~new_n10197_;
  assign new_n10199_ = new_n599_ & ~new_n10198_;
  assign new_n10200_ = ~new_n10004_ & new_n10199_;
  assign new_n10201_ = ~new_n10194_ & ~new_n10200_;
  assign new_n10202_ = ~\b[16]  & ~new_n10201_;
  assign new_n10203_ = ~new_n9709_ & ~\quotient[27] ;
  assign new_n10204_ = ~new_n9719_ & new_n9892_;
  assign new_n10205_ = ~new_n9888_ & new_n10204_;
  assign new_n10206_ = ~new_n9889_ & ~new_n9892_;
  assign new_n10207_ = ~new_n10205_ & ~new_n10206_;
  assign new_n10208_ = new_n599_ & ~new_n10207_;
  assign new_n10209_ = ~new_n10004_ & new_n10208_;
  assign new_n10210_ = ~new_n10203_ & ~new_n10209_;
  assign new_n10211_ = ~\b[15]  & ~new_n10210_;
  assign new_n10212_ = ~new_n9718_ & ~\quotient[27] ;
  assign new_n10213_ = ~new_n9728_ & new_n9887_;
  assign new_n10214_ = ~new_n9883_ & new_n10213_;
  assign new_n10215_ = ~new_n9884_ & ~new_n9887_;
  assign new_n10216_ = ~new_n10214_ & ~new_n10215_;
  assign new_n10217_ = new_n599_ & ~new_n10216_;
  assign new_n10218_ = ~new_n10004_ & new_n10217_;
  assign new_n10219_ = ~new_n10212_ & ~new_n10218_;
  assign new_n10220_ = ~\b[14]  & ~new_n10219_;
  assign new_n10221_ = ~new_n9727_ & ~\quotient[27] ;
  assign new_n10222_ = ~new_n9737_ & new_n9882_;
  assign new_n10223_ = ~new_n9878_ & new_n10222_;
  assign new_n10224_ = ~new_n9879_ & ~new_n9882_;
  assign new_n10225_ = ~new_n10223_ & ~new_n10224_;
  assign new_n10226_ = new_n599_ & ~new_n10225_;
  assign new_n10227_ = ~new_n10004_ & new_n10226_;
  assign new_n10228_ = ~new_n10221_ & ~new_n10227_;
  assign new_n10229_ = ~\b[13]  & ~new_n10228_;
  assign new_n10230_ = ~new_n9736_ & ~\quotient[27] ;
  assign new_n10231_ = ~new_n9746_ & new_n9877_;
  assign new_n10232_ = ~new_n9873_ & new_n10231_;
  assign new_n10233_ = ~new_n9874_ & ~new_n9877_;
  assign new_n10234_ = ~new_n10232_ & ~new_n10233_;
  assign new_n10235_ = new_n599_ & ~new_n10234_;
  assign new_n10236_ = ~new_n10004_ & new_n10235_;
  assign new_n10237_ = ~new_n10230_ & ~new_n10236_;
  assign new_n10238_ = ~\b[12]  & ~new_n10237_;
  assign new_n10239_ = ~new_n9745_ & ~\quotient[27] ;
  assign new_n10240_ = ~new_n9755_ & new_n9872_;
  assign new_n10241_ = ~new_n9868_ & new_n10240_;
  assign new_n10242_ = ~new_n9869_ & ~new_n9872_;
  assign new_n10243_ = ~new_n10241_ & ~new_n10242_;
  assign new_n10244_ = new_n599_ & ~new_n10243_;
  assign new_n10245_ = ~new_n10004_ & new_n10244_;
  assign new_n10246_ = ~new_n10239_ & ~new_n10245_;
  assign new_n10247_ = ~\b[11]  & ~new_n10246_;
  assign new_n10248_ = ~new_n9754_ & ~\quotient[27] ;
  assign new_n10249_ = ~new_n9764_ & new_n9867_;
  assign new_n10250_ = ~new_n9863_ & new_n10249_;
  assign new_n10251_ = ~new_n9864_ & ~new_n9867_;
  assign new_n10252_ = ~new_n10250_ & ~new_n10251_;
  assign new_n10253_ = new_n599_ & ~new_n10252_;
  assign new_n10254_ = ~new_n10004_ & new_n10253_;
  assign new_n10255_ = ~new_n10248_ & ~new_n10254_;
  assign new_n10256_ = ~\b[10]  & ~new_n10255_;
  assign new_n10257_ = ~new_n9763_ & ~\quotient[27] ;
  assign new_n10258_ = ~new_n9773_ & new_n9862_;
  assign new_n10259_ = ~new_n9858_ & new_n10258_;
  assign new_n10260_ = ~new_n9859_ & ~new_n9862_;
  assign new_n10261_ = ~new_n10259_ & ~new_n10260_;
  assign new_n10262_ = new_n599_ & ~new_n10261_;
  assign new_n10263_ = ~new_n10004_ & new_n10262_;
  assign new_n10264_ = ~new_n10257_ & ~new_n10263_;
  assign new_n10265_ = ~\b[9]  & ~new_n10264_;
  assign new_n10266_ = ~new_n9772_ & ~\quotient[27] ;
  assign new_n10267_ = ~new_n9782_ & new_n9857_;
  assign new_n10268_ = ~new_n9853_ & new_n10267_;
  assign new_n10269_ = ~new_n9854_ & ~new_n9857_;
  assign new_n10270_ = ~new_n10268_ & ~new_n10269_;
  assign new_n10271_ = new_n599_ & ~new_n10270_;
  assign new_n10272_ = ~new_n10004_ & new_n10271_;
  assign new_n10273_ = ~new_n10266_ & ~new_n10272_;
  assign new_n10274_ = ~\b[8]  & ~new_n10273_;
  assign new_n10275_ = ~new_n9781_ & ~\quotient[27] ;
  assign new_n10276_ = ~new_n9791_ & new_n9852_;
  assign new_n10277_ = ~new_n9848_ & new_n10276_;
  assign new_n10278_ = ~new_n9849_ & ~new_n9852_;
  assign new_n10279_ = ~new_n10277_ & ~new_n10278_;
  assign new_n10280_ = new_n599_ & ~new_n10279_;
  assign new_n10281_ = ~new_n10004_ & new_n10280_;
  assign new_n10282_ = ~new_n10275_ & ~new_n10281_;
  assign new_n10283_ = ~\b[7]  & ~new_n10282_;
  assign new_n10284_ = ~new_n9790_ & ~\quotient[27] ;
  assign new_n10285_ = ~new_n9800_ & new_n9847_;
  assign new_n10286_ = ~new_n9843_ & new_n10285_;
  assign new_n10287_ = ~new_n9844_ & ~new_n9847_;
  assign new_n10288_ = ~new_n10286_ & ~new_n10287_;
  assign new_n10289_ = new_n599_ & ~new_n10288_;
  assign new_n10290_ = ~new_n10004_ & new_n10289_;
  assign new_n10291_ = ~new_n10284_ & ~new_n10290_;
  assign new_n10292_ = ~\b[6]  & ~new_n10291_;
  assign new_n10293_ = ~new_n9799_ & ~\quotient[27] ;
  assign new_n10294_ = ~new_n9809_ & new_n9842_;
  assign new_n10295_ = ~new_n9838_ & new_n10294_;
  assign new_n10296_ = ~new_n9839_ & ~new_n9842_;
  assign new_n10297_ = ~new_n10295_ & ~new_n10296_;
  assign new_n10298_ = new_n599_ & ~new_n10297_;
  assign new_n10299_ = ~new_n10004_ & new_n10298_;
  assign new_n10300_ = ~new_n10293_ & ~new_n10299_;
  assign new_n10301_ = ~\b[5]  & ~new_n10300_;
  assign new_n10302_ = ~new_n9808_ & ~\quotient[27] ;
  assign new_n10303_ = ~new_n9817_ & new_n9837_;
  assign new_n10304_ = ~new_n9833_ & new_n10303_;
  assign new_n10305_ = ~new_n9834_ & ~new_n9837_;
  assign new_n10306_ = ~new_n10304_ & ~new_n10305_;
  assign new_n10307_ = new_n599_ & ~new_n10306_;
  assign new_n10308_ = ~new_n10004_ & new_n10307_;
  assign new_n10309_ = ~new_n10302_ & ~new_n10308_;
  assign new_n10310_ = ~\b[4]  & ~new_n10309_;
  assign new_n10311_ = ~new_n9816_ & ~\quotient[27] ;
  assign new_n10312_ = ~new_n9828_ & new_n9832_;
  assign new_n10313_ = ~new_n9827_ & new_n10312_;
  assign new_n10314_ = ~new_n9829_ & ~new_n9832_;
  assign new_n10315_ = ~new_n10313_ & ~new_n10314_;
  assign new_n10316_ = new_n599_ & ~new_n10315_;
  assign new_n10317_ = ~new_n10004_ & new_n10316_;
  assign new_n10318_ = ~new_n10311_ & ~new_n10317_;
  assign new_n10319_ = ~\b[3]  & ~new_n10318_;
  assign new_n10320_ = ~new_n9821_ & ~\quotient[27] ;
  assign new_n10321_ = ~new_n9824_ & new_n9826_;
  assign new_n10322_ = ~new_n9822_ & new_n10321_;
  assign new_n10323_ = new_n599_ & ~new_n10322_;
  assign new_n10324_ = ~new_n9827_ & new_n10323_;
  assign new_n10325_ = ~new_n10004_ & new_n10324_;
  assign new_n10326_ = ~new_n10320_ & ~new_n10325_;
  assign new_n10327_ = ~\b[2]  & ~new_n10326_;
  assign new_n10328_ = \b[0]  & ~\b[37] ;
  assign new_n10329_ = new_n293_ & new_n10328_;
  assign new_n10330_ = new_n291_ & new_n10329_;
  assign new_n10331_ = new_n302_ & new_n10330_;
  assign new_n10332_ = new_n288_ & new_n10331_;
  assign new_n10333_ = ~new_n10004_ & new_n10332_;
  assign new_n10334_ = \a[27]  & ~new_n10333_;
  assign new_n10335_ = new_n411_ & new_n9826_;
  assign new_n10336_ = new_n422_ & new_n10335_;
  assign new_n10337_ = new_n408_ & new_n10336_;
  assign new_n10338_ = ~new_n10004_ & new_n10337_;
  assign new_n10339_ = ~new_n10334_ & ~new_n10338_;
  assign new_n10340_ = \b[1]  & ~new_n10339_;
  assign new_n10341_ = ~\b[1]  & ~new_n10338_;
  assign new_n10342_ = ~new_n10334_ & new_n10341_;
  assign new_n10343_ = ~new_n10340_ & ~new_n10342_;
  assign new_n10344_ = ~\a[26]  & \b[0] ;
  assign new_n10345_ = ~new_n10343_ & ~new_n10344_;
  assign new_n10346_ = ~\b[1]  & ~new_n10339_;
  assign new_n10347_ = ~new_n10345_ & ~new_n10346_;
  assign new_n10348_ = \b[2]  & ~new_n10325_;
  assign new_n10349_ = ~new_n10320_ & new_n10348_;
  assign new_n10350_ = ~new_n10327_ & ~new_n10349_;
  assign new_n10351_ = ~new_n10347_ & new_n10350_;
  assign new_n10352_ = ~new_n10327_ & ~new_n10351_;
  assign new_n10353_ = \b[3]  & ~new_n10317_;
  assign new_n10354_ = ~new_n10311_ & new_n10353_;
  assign new_n10355_ = ~new_n10319_ & ~new_n10354_;
  assign new_n10356_ = ~new_n10352_ & new_n10355_;
  assign new_n10357_ = ~new_n10319_ & ~new_n10356_;
  assign new_n10358_ = \b[4]  & ~new_n10308_;
  assign new_n10359_ = ~new_n10302_ & new_n10358_;
  assign new_n10360_ = ~new_n10310_ & ~new_n10359_;
  assign new_n10361_ = ~new_n10357_ & new_n10360_;
  assign new_n10362_ = ~new_n10310_ & ~new_n10361_;
  assign new_n10363_ = \b[5]  & ~new_n10299_;
  assign new_n10364_ = ~new_n10293_ & new_n10363_;
  assign new_n10365_ = ~new_n10301_ & ~new_n10364_;
  assign new_n10366_ = ~new_n10362_ & new_n10365_;
  assign new_n10367_ = ~new_n10301_ & ~new_n10366_;
  assign new_n10368_ = \b[6]  & ~new_n10290_;
  assign new_n10369_ = ~new_n10284_ & new_n10368_;
  assign new_n10370_ = ~new_n10292_ & ~new_n10369_;
  assign new_n10371_ = ~new_n10367_ & new_n10370_;
  assign new_n10372_ = ~new_n10292_ & ~new_n10371_;
  assign new_n10373_ = \b[7]  & ~new_n10281_;
  assign new_n10374_ = ~new_n10275_ & new_n10373_;
  assign new_n10375_ = ~new_n10283_ & ~new_n10374_;
  assign new_n10376_ = ~new_n10372_ & new_n10375_;
  assign new_n10377_ = ~new_n10283_ & ~new_n10376_;
  assign new_n10378_ = \b[8]  & ~new_n10272_;
  assign new_n10379_ = ~new_n10266_ & new_n10378_;
  assign new_n10380_ = ~new_n10274_ & ~new_n10379_;
  assign new_n10381_ = ~new_n10377_ & new_n10380_;
  assign new_n10382_ = ~new_n10274_ & ~new_n10381_;
  assign new_n10383_ = \b[9]  & ~new_n10263_;
  assign new_n10384_ = ~new_n10257_ & new_n10383_;
  assign new_n10385_ = ~new_n10265_ & ~new_n10384_;
  assign new_n10386_ = ~new_n10382_ & new_n10385_;
  assign new_n10387_ = ~new_n10265_ & ~new_n10386_;
  assign new_n10388_ = \b[10]  & ~new_n10254_;
  assign new_n10389_ = ~new_n10248_ & new_n10388_;
  assign new_n10390_ = ~new_n10256_ & ~new_n10389_;
  assign new_n10391_ = ~new_n10387_ & new_n10390_;
  assign new_n10392_ = ~new_n10256_ & ~new_n10391_;
  assign new_n10393_ = \b[11]  & ~new_n10245_;
  assign new_n10394_ = ~new_n10239_ & new_n10393_;
  assign new_n10395_ = ~new_n10247_ & ~new_n10394_;
  assign new_n10396_ = ~new_n10392_ & new_n10395_;
  assign new_n10397_ = ~new_n10247_ & ~new_n10396_;
  assign new_n10398_ = \b[12]  & ~new_n10236_;
  assign new_n10399_ = ~new_n10230_ & new_n10398_;
  assign new_n10400_ = ~new_n10238_ & ~new_n10399_;
  assign new_n10401_ = ~new_n10397_ & new_n10400_;
  assign new_n10402_ = ~new_n10238_ & ~new_n10401_;
  assign new_n10403_ = \b[13]  & ~new_n10227_;
  assign new_n10404_ = ~new_n10221_ & new_n10403_;
  assign new_n10405_ = ~new_n10229_ & ~new_n10404_;
  assign new_n10406_ = ~new_n10402_ & new_n10405_;
  assign new_n10407_ = ~new_n10229_ & ~new_n10406_;
  assign new_n10408_ = \b[14]  & ~new_n10218_;
  assign new_n10409_ = ~new_n10212_ & new_n10408_;
  assign new_n10410_ = ~new_n10220_ & ~new_n10409_;
  assign new_n10411_ = ~new_n10407_ & new_n10410_;
  assign new_n10412_ = ~new_n10220_ & ~new_n10411_;
  assign new_n10413_ = \b[15]  & ~new_n10209_;
  assign new_n10414_ = ~new_n10203_ & new_n10413_;
  assign new_n10415_ = ~new_n10211_ & ~new_n10414_;
  assign new_n10416_ = ~new_n10412_ & new_n10415_;
  assign new_n10417_ = ~new_n10211_ & ~new_n10416_;
  assign new_n10418_ = \b[16]  & ~new_n10200_;
  assign new_n10419_ = ~new_n10194_ & new_n10418_;
  assign new_n10420_ = ~new_n10202_ & ~new_n10419_;
  assign new_n10421_ = ~new_n10417_ & new_n10420_;
  assign new_n10422_ = ~new_n10202_ & ~new_n10421_;
  assign new_n10423_ = \b[17]  & ~new_n10191_;
  assign new_n10424_ = ~new_n10185_ & new_n10423_;
  assign new_n10425_ = ~new_n10193_ & ~new_n10424_;
  assign new_n10426_ = ~new_n10422_ & new_n10425_;
  assign new_n10427_ = ~new_n10193_ & ~new_n10426_;
  assign new_n10428_ = \b[18]  & ~new_n10182_;
  assign new_n10429_ = ~new_n10176_ & new_n10428_;
  assign new_n10430_ = ~new_n10184_ & ~new_n10429_;
  assign new_n10431_ = ~new_n10427_ & new_n10430_;
  assign new_n10432_ = ~new_n10184_ & ~new_n10431_;
  assign new_n10433_ = \b[19]  & ~new_n10173_;
  assign new_n10434_ = ~new_n10167_ & new_n10433_;
  assign new_n10435_ = ~new_n10175_ & ~new_n10434_;
  assign new_n10436_ = ~new_n10432_ & new_n10435_;
  assign new_n10437_ = ~new_n10175_ & ~new_n10436_;
  assign new_n10438_ = \b[20]  & ~new_n10164_;
  assign new_n10439_ = ~new_n10158_ & new_n10438_;
  assign new_n10440_ = ~new_n10166_ & ~new_n10439_;
  assign new_n10441_ = ~new_n10437_ & new_n10440_;
  assign new_n10442_ = ~new_n10166_ & ~new_n10441_;
  assign new_n10443_ = \b[21]  & ~new_n10155_;
  assign new_n10444_ = ~new_n10149_ & new_n10443_;
  assign new_n10445_ = ~new_n10157_ & ~new_n10444_;
  assign new_n10446_ = ~new_n10442_ & new_n10445_;
  assign new_n10447_ = ~new_n10157_ & ~new_n10446_;
  assign new_n10448_ = \b[22]  & ~new_n10146_;
  assign new_n10449_ = ~new_n10140_ & new_n10448_;
  assign new_n10450_ = ~new_n10148_ & ~new_n10449_;
  assign new_n10451_ = ~new_n10447_ & new_n10450_;
  assign new_n10452_ = ~new_n10148_ & ~new_n10451_;
  assign new_n10453_ = \b[23]  & ~new_n10137_;
  assign new_n10454_ = ~new_n10131_ & new_n10453_;
  assign new_n10455_ = ~new_n10139_ & ~new_n10454_;
  assign new_n10456_ = ~new_n10452_ & new_n10455_;
  assign new_n10457_ = ~new_n10139_ & ~new_n10456_;
  assign new_n10458_ = \b[24]  & ~new_n10128_;
  assign new_n10459_ = ~new_n10122_ & new_n10458_;
  assign new_n10460_ = ~new_n10130_ & ~new_n10459_;
  assign new_n10461_ = ~new_n10457_ & new_n10460_;
  assign new_n10462_ = ~new_n10130_ & ~new_n10461_;
  assign new_n10463_ = \b[25]  & ~new_n10119_;
  assign new_n10464_ = ~new_n10113_ & new_n10463_;
  assign new_n10465_ = ~new_n10121_ & ~new_n10464_;
  assign new_n10466_ = ~new_n10462_ & new_n10465_;
  assign new_n10467_ = ~new_n10121_ & ~new_n10466_;
  assign new_n10468_ = \b[26]  & ~new_n10110_;
  assign new_n10469_ = ~new_n10104_ & new_n10468_;
  assign new_n10470_ = ~new_n10112_ & ~new_n10469_;
  assign new_n10471_ = ~new_n10467_ & new_n10470_;
  assign new_n10472_ = ~new_n10112_ & ~new_n10471_;
  assign new_n10473_ = \b[27]  & ~new_n10101_;
  assign new_n10474_ = ~new_n10095_ & new_n10473_;
  assign new_n10475_ = ~new_n10103_ & ~new_n10474_;
  assign new_n10476_ = ~new_n10472_ & new_n10475_;
  assign new_n10477_ = ~new_n10103_ & ~new_n10476_;
  assign new_n10478_ = \b[28]  & ~new_n10092_;
  assign new_n10479_ = ~new_n10086_ & new_n10478_;
  assign new_n10480_ = ~new_n10094_ & ~new_n10479_;
  assign new_n10481_ = ~new_n10477_ & new_n10480_;
  assign new_n10482_ = ~new_n10094_ & ~new_n10481_;
  assign new_n10483_ = \b[29]  & ~new_n10083_;
  assign new_n10484_ = ~new_n10077_ & new_n10483_;
  assign new_n10485_ = ~new_n10085_ & ~new_n10484_;
  assign new_n10486_ = ~new_n10482_ & new_n10485_;
  assign new_n10487_ = ~new_n10085_ & ~new_n10486_;
  assign new_n10488_ = \b[30]  & ~new_n10074_;
  assign new_n10489_ = ~new_n10068_ & new_n10488_;
  assign new_n10490_ = ~new_n10076_ & ~new_n10489_;
  assign new_n10491_ = ~new_n10487_ & new_n10490_;
  assign new_n10492_ = ~new_n10076_ & ~new_n10491_;
  assign new_n10493_ = \b[31]  & ~new_n10065_;
  assign new_n10494_ = ~new_n10059_ & new_n10493_;
  assign new_n10495_ = ~new_n10067_ & ~new_n10494_;
  assign new_n10496_ = ~new_n10492_ & new_n10495_;
  assign new_n10497_ = ~new_n10067_ & ~new_n10496_;
  assign new_n10498_ = \b[32]  & ~new_n10056_;
  assign new_n10499_ = ~new_n10050_ & new_n10498_;
  assign new_n10500_ = ~new_n10058_ & ~new_n10499_;
  assign new_n10501_ = ~new_n10497_ & new_n10500_;
  assign new_n10502_ = ~new_n10058_ & ~new_n10501_;
  assign new_n10503_ = \b[33]  & ~new_n10047_;
  assign new_n10504_ = ~new_n10041_ & new_n10503_;
  assign new_n10505_ = ~new_n10049_ & ~new_n10504_;
  assign new_n10506_ = ~new_n10502_ & new_n10505_;
  assign new_n10507_ = ~new_n10049_ & ~new_n10506_;
  assign new_n10508_ = \b[34]  & ~new_n10038_;
  assign new_n10509_ = ~new_n10032_ & new_n10508_;
  assign new_n10510_ = ~new_n10040_ & ~new_n10509_;
  assign new_n10511_ = ~new_n10507_ & new_n10510_;
  assign new_n10512_ = ~new_n10040_ & ~new_n10511_;
  assign new_n10513_ = \b[35]  & ~new_n10029_;
  assign new_n10514_ = ~new_n10023_ & new_n10513_;
  assign new_n10515_ = ~new_n10031_ & ~new_n10514_;
  assign new_n10516_ = ~new_n10512_ & new_n10515_;
  assign new_n10517_ = ~new_n10031_ & ~new_n10516_;
  assign new_n10518_ = \b[36]  & ~new_n10012_;
  assign new_n10519_ = ~new_n10006_ & new_n10518_;
  assign new_n10520_ = ~new_n10022_ & ~new_n10519_;
  assign new_n10521_ = ~new_n10517_ & new_n10520_;
  assign new_n10522_ = ~new_n10022_ & ~new_n10521_;
  assign new_n10523_ = \b[37]  & ~new_n10014_;
  assign new_n10524_ = ~new_n10019_ & new_n10523_;
  assign new_n10525_ = ~new_n10021_ & ~new_n10524_;
  assign new_n10526_ = ~new_n10522_ & new_n10525_;
  assign new_n10527_ = ~new_n10021_ & ~new_n10526_;
  assign new_n10528_ = new_n291_ & new_n293_;
  assign new_n10529_ = new_n302_ & new_n10528_;
  assign new_n10530_ = new_n288_ & new_n10529_;
  assign \quotient[26]  = ~new_n10527_ & new_n10530_;
  assign new_n10532_ = ~new_n10013_ & ~\quotient[26] ;
  assign new_n10533_ = ~new_n10031_ & new_n10520_;
  assign new_n10534_ = ~new_n10516_ & new_n10533_;
  assign new_n10535_ = ~new_n10517_ & ~new_n10520_;
  assign new_n10536_ = ~new_n10534_ & ~new_n10535_;
  assign new_n10537_ = new_n10530_ & ~new_n10536_;
  assign new_n10538_ = ~new_n10527_ & new_n10537_;
  assign new_n10539_ = ~new_n10532_ & ~new_n10538_;
  assign new_n10540_ = ~\b[37]  & ~new_n10539_;
  assign new_n10541_ = ~new_n10030_ & ~\quotient[26] ;
  assign new_n10542_ = ~new_n10040_ & new_n10515_;
  assign new_n10543_ = ~new_n10511_ & new_n10542_;
  assign new_n10544_ = ~new_n10512_ & ~new_n10515_;
  assign new_n10545_ = ~new_n10543_ & ~new_n10544_;
  assign new_n10546_ = new_n10530_ & ~new_n10545_;
  assign new_n10547_ = ~new_n10527_ & new_n10546_;
  assign new_n10548_ = ~new_n10541_ & ~new_n10547_;
  assign new_n10549_ = ~\b[36]  & ~new_n10548_;
  assign new_n10550_ = ~new_n10039_ & ~\quotient[26] ;
  assign new_n10551_ = ~new_n10049_ & new_n10510_;
  assign new_n10552_ = ~new_n10506_ & new_n10551_;
  assign new_n10553_ = ~new_n10507_ & ~new_n10510_;
  assign new_n10554_ = ~new_n10552_ & ~new_n10553_;
  assign new_n10555_ = new_n10530_ & ~new_n10554_;
  assign new_n10556_ = ~new_n10527_ & new_n10555_;
  assign new_n10557_ = ~new_n10550_ & ~new_n10556_;
  assign new_n10558_ = ~\b[35]  & ~new_n10557_;
  assign new_n10559_ = ~new_n10048_ & ~\quotient[26] ;
  assign new_n10560_ = ~new_n10058_ & new_n10505_;
  assign new_n10561_ = ~new_n10501_ & new_n10560_;
  assign new_n10562_ = ~new_n10502_ & ~new_n10505_;
  assign new_n10563_ = ~new_n10561_ & ~new_n10562_;
  assign new_n10564_ = new_n10530_ & ~new_n10563_;
  assign new_n10565_ = ~new_n10527_ & new_n10564_;
  assign new_n10566_ = ~new_n10559_ & ~new_n10565_;
  assign new_n10567_ = ~\b[34]  & ~new_n10566_;
  assign new_n10568_ = ~new_n10057_ & ~\quotient[26] ;
  assign new_n10569_ = ~new_n10067_ & new_n10500_;
  assign new_n10570_ = ~new_n10496_ & new_n10569_;
  assign new_n10571_ = ~new_n10497_ & ~new_n10500_;
  assign new_n10572_ = ~new_n10570_ & ~new_n10571_;
  assign new_n10573_ = new_n10530_ & ~new_n10572_;
  assign new_n10574_ = ~new_n10527_ & new_n10573_;
  assign new_n10575_ = ~new_n10568_ & ~new_n10574_;
  assign new_n10576_ = ~\b[33]  & ~new_n10575_;
  assign new_n10577_ = ~new_n10066_ & ~\quotient[26] ;
  assign new_n10578_ = ~new_n10076_ & new_n10495_;
  assign new_n10579_ = ~new_n10491_ & new_n10578_;
  assign new_n10580_ = ~new_n10492_ & ~new_n10495_;
  assign new_n10581_ = ~new_n10579_ & ~new_n10580_;
  assign new_n10582_ = new_n10530_ & ~new_n10581_;
  assign new_n10583_ = ~new_n10527_ & new_n10582_;
  assign new_n10584_ = ~new_n10577_ & ~new_n10583_;
  assign new_n10585_ = ~\b[32]  & ~new_n10584_;
  assign new_n10586_ = ~new_n10075_ & ~\quotient[26] ;
  assign new_n10587_ = ~new_n10085_ & new_n10490_;
  assign new_n10588_ = ~new_n10486_ & new_n10587_;
  assign new_n10589_ = ~new_n10487_ & ~new_n10490_;
  assign new_n10590_ = ~new_n10588_ & ~new_n10589_;
  assign new_n10591_ = new_n10530_ & ~new_n10590_;
  assign new_n10592_ = ~new_n10527_ & new_n10591_;
  assign new_n10593_ = ~new_n10586_ & ~new_n10592_;
  assign new_n10594_ = ~\b[31]  & ~new_n10593_;
  assign new_n10595_ = ~new_n10084_ & ~\quotient[26] ;
  assign new_n10596_ = ~new_n10094_ & new_n10485_;
  assign new_n10597_ = ~new_n10481_ & new_n10596_;
  assign new_n10598_ = ~new_n10482_ & ~new_n10485_;
  assign new_n10599_ = ~new_n10597_ & ~new_n10598_;
  assign new_n10600_ = new_n10530_ & ~new_n10599_;
  assign new_n10601_ = ~new_n10527_ & new_n10600_;
  assign new_n10602_ = ~new_n10595_ & ~new_n10601_;
  assign new_n10603_ = ~\b[30]  & ~new_n10602_;
  assign new_n10604_ = ~new_n10093_ & ~\quotient[26] ;
  assign new_n10605_ = ~new_n10103_ & new_n10480_;
  assign new_n10606_ = ~new_n10476_ & new_n10605_;
  assign new_n10607_ = ~new_n10477_ & ~new_n10480_;
  assign new_n10608_ = ~new_n10606_ & ~new_n10607_;
  assign new_n10609_ = new_n10530_ & ~new_n10608_;
  assign new_n10610_ = ~new_n10527_ & new_n10609_;
  assign new_n10611_ = ~new_n10604_ & ~new_n10610_;
  assign new_n10612_ = ~\b[29]  & ~new_n10611_;
  assign new_n10613_ = ~new_n10102_ & ~\quotient[26] ;
  assign new_n10614_ = ~new_n10112_ & new_n10475_;
  assign new_n10615_ = ~new_n10471_ & new_n10614_;
  assign new_n10616_ = ~new_n10472_ & ~new_n10475_;
  assign new_n10617_ = ~new_n10615_ & ~new_n10616_;
  assign new_n10618_ = new_n10530_ & ~new_n10617_;
  assign new_n10619_ = ~new_n10527_ & new_n10618_;
  assign new_n10620_ = ~new_n10613_ & ~new_n10619_;
  assign new_n10621_ = ~\b[28]  & ~new_n10620_;
  assign new_n10622_ = ~new_n10111_ & ~\quotient[26] ;
  assign new_n10623_ = ~new_n10121_ & new_n10470_;
  assign new_n10624_ = ~new_n10466_ & new_n10623_;
  assign new_n10625_ = ~new_n10467_ & ~new_n10470_;
  assign new_n10626_ = ~new_n10624_ & ~new_n10625_;
  assign new_n10627_ = new_n10530_ & ~new_n10626_;
  assign new_n10628_ = ~new_n10527_ & new_n10627_;
  assign new_n10629_ = ~new_n10622_ & ~new_n10628_;
  assign new_n10630_ = ~\b[27]  & ~new_n10629_;
  assign new_n10631_ = ~new_n10120_ & ~\quotient[26] ;
  assign new_n10632_ = ~new_n10130_ & new_n10465_;
  assign new_n10633_ = ~new_n10461_ & new_n10632_;
  assign new_n10634_ = ~new_n10462_ & ~new_n10465_;
  assign new_n10635_ = ~new_n10633_ & ~new_n10634_;
  assign new_n10636_ = new_n10530_ & ~new_n10635_;
  assign new_n10637_ = ~new_n10527_ & new_n10636_;
  assign new_n10638_ = ~new_n10631_ & ~new_n10637_;
  assign new_n10639_ = ~\b[26]  & ~new_n10638_;
  assign new_n10640_ = ~new_n10129_ & ~\quotient[26] ;
  assign new_n10641_ = ~new_n10139_ & new_n10460_;
  assign new_n10642_ = ~new_n10456_ & new_n10641_;
  assign new_n10643_ = ~new_n10457_ & ~new_n10460_;
  assign new_n10644_ = ~new_n10642_ & ~new_n10643_;
  assign new_n10645_ = new_n10530_ & ~new_n10644_;
  assign new_n10646_ = ~new_n10527_ & new_n10645_;
  assign new_n10647_ = ~new_n10640_ & ~new_n10646_;
  assign new_n10648_ = ~\b[25]  & ~new_n10647_;
  assign new_n10649_ = ~new_n10138_ & ~\quotient[26] ;
  assign new_n10650_ = ~new_n10148_ & new_n10455_;
  assign new_n10651_ = ~new_n10451_ & new_n10650_;
  assign new_n10652_ = ~new_n10452_ & ~new_n10455_;
  assign new_n10653_ = ~new_n10651_ & ~new_n10652_;
  assign new_n10654_ = new_n10530_ & ~new_n10653_;
  assign new_n10655_ = ~new_n10527_ & new_n10654_;
  assign new_n10656_ = ~new_n10649_ & ~new_n10655_;
  assign new_n10657_ = ~\b[24]  & ~new_n10656_;
  assign new_n10658_ = ~new_n10147_ & ~\quotient[26] ;
  assign new_n10659_ = ~new_n10157_ & new_n10450_;
  assign new_n10660_ = ~new_n10446_ & new_n10659_;
  assign new_n10661_ = ~new_n10447_ & ~new_n10450_;
  assign new_n10662_ = ~new_n10660_ & ~new_n10661_;
  assign new_n10663_ = new_n10530_ & ~new_n10662_;
  assign new_n10664_ = ~new_n10527_ & new_n10663_;
  assign new_n10665_ = ~new_n10658_ & ~new_n10664_;
  assign new_n10666_ = ~\b[23]  & ~new_n10665_;
  assign new_n10667_ = ~new_n10156_ & ~\quotient[26] ;
  assign new_n10668_ = ~new_n10166_ & new_n10445_;
  assign new_n10669_ = ~new_n10441_ & new_n10668_;
  assign new_n10670_ = ~new_n10442_ & ~new_n10445_;
  assign new_n10671_ = ~new_n10669_ & ~new_n10670_;
  assign new_n10672_ = new_n10530_ & ~new_n10671_;
  assign new_n10673_ = ~new_n10527_ & new_n10672_;
  assign new_n10674_ = ~new_n10667_ & ~new_n10673_;
  assign new_n10675_ = ~\b[22]  & ~new_n10674_;
  assign new_n10676_ = ~new_n10165_ & ~\quotient[26] ;
  assign new_n10677_ = ~new_n10175_ & new_n10440_;
  assign new_n10678_ = ~new_n10436_ & new_n10677_;
  assign new_n10679_ = ~new_n10437_ & ~new_n10440_;
  assign new_n10680_ = ~new_n10678_ & ~new_n10679_;
  assign new_n10681_ = new_n10530_ & ~new_n10680_;
  assign new_n10682_ = ~new_n10527_ & new_n10681_;
  assign new_n10683_ = ~new_n10676_ & ~new_n10682_;
  assign new_n10684_ = ~\b[21]  & ~new_n10683_;
  assign new_n10685_ = ~new_n10174_ & ~\quotient[26] ;
  assign new_n10686_ = ~new_n10184_ & new_n10435_;
  assign new_n10687_ = ~new_n10431_ & new_n10686_;
  assign new_n10688_ = ~new_n10432_ & ~new_n10435_;
  assign new_n10689_ = ~new_n10687_ & ~new_n10688_;
  assign new_n10690_ = new_n10530_ & ~new_n10689_;
  assign new_n10691_ = ~new_n10527_ & new_n10690_;
  assign new_n10692_ = ~new_n10685_ & ~new_n10691_;
  assign new_n10693_ = ~\b[20]  & ~new_n10692_;
  assign new_n10694_ = ~new_n10183_ & ~\quotient[26] ;
  assign new_n10695_ = ~new_n10193_ & new_n10430_;
  assign new_n10696_ = ~new_n10426_ & new_n10695_;
  assign new_n10697_ = ~new_n10427_ & ~new_n10430_;
  assign new_n10698_ = ~new_n10696_ & ~new_n10697_;
  assign new_n10699_ = new_n10530_ & ~new_n10698_;
  assign new_n10700_ = ~new_n10527_ & new_n10699_;
  assign new_n10701_ = ~new_n10694_ & ~new_n10700_;
  assign new_n10702_ = ~\b[19]  & ~new_n10701_;
  assign new_n10703_ = ~new_n10192_ & ~\quotient[26] ;
  assign new_n10704_ = ~new_n10202_ & new_n10425_;
  assign new_n10705_ = ~new_n10421_ & new_n10704_;
  assign new_n10706_ = ~new_n10422_ & ~new_n10425_;
  assign new_n10707_ = ~new_n10705_ & ~new_n10706_;
  assign new_n10708_ = new_n10530_ & ~new_n10707_;
  assign new_n10709_ = ~new_n10527_ & new_n10708_;
  assign new_n10710_ = ~new_n10703_ & ~new_n10709_;
  assign new_n10711_ = ~\b[18]  & ~new_n10710_;
  assign new_n10712_ = ~new_n10201_ & ~\quotient[26] ;
  assign new_n10713_ = ~new_n10211_ & new_n10420_;
  assign new_n10714_ = ~new_n10416_ & new_n10713_;
  assign new_n10715_ = ~new_n10417_ & ~new_n10420_;
  assign new_n10716_ = ~new_n10714_ & ~new_n10715_;
  assign new_n10717_ = new_n10530_ & ~new_n10716_;
  assign new_n10718_ = ~new_n10527_ & new_n10717_;
  assign new_n10719_ = ~new_n10712_ & ~new_n10718_;
  assign new_n10720_ = ~\b[17]  & ~new_n10719_;
  assign new_n10721_ = ~new_n10210_ & ~\quotient[26] ;
  assign new_n10722_ = ~new_n10220_ & new_n10415_;
  assign new_n10723_ = ~new_n10411_ & new_n10722_;
  assign new_n10724_ = ~new_n10412_ & ~new_n10415_;
  assign new_n10725_ = ~new_n10723_ & ~new_n10724_;
  assign new_n10726_ = new_n10530_ & ~new_n10725_;
  assign new_n10727_ = ~new_n10527_ & new_n10726_;
  assign new_n10728_ = ~new_n10721_ & ~new_n10727_;
  assign new_n10729_ = ~\b[16]  & ~new_n10728_;
  assign new_n10730_ = ~new_n10219_ & ~\quotient[26] ;
  assign new_n10731_ = ~new_n10229_ & new_n10410_;
  assign new_n10732_ = ~new_n10406_ & new_n10731_;
  assign new_n10733_ = ~new_n10407_ & ~new_n10410_;
  assign new_n10734_ = ~new_n10732_ & ~new_n10733_;
  assign new_n10735_ = new_n10530_ & ~new_n10734_;
  assign new_n10736_ = ~new_n10527_ & new_n10735_;
  assign new_n10737_ = ~new_n10730_ & ~new_n10736_;
  assign new_n10738_ = ~\b[15]  & ~new_n10737_;
  assign new_n10739_ = ~new_n10228_ & ~\quotient[26] ;
  assign new_n10740_ = ~new_n10238_ & new_n10405_;
  assign new_n10741_ = ~new_n10401_ & new_n10740_;
  assign new_n10742_ = ~new_n10402_ & ~new_n10405_;
  assign new_n10743_ = ~new_n10741_ & ~new_n10742_;
  assign new_n10744_ = new_n10530_ & ~new_n10743_;
  assign new_n10745_ = ~new_n10527_ & new_n10744_;
  assign new_n10746_ = ~new_n10739_ & ~new_n10745_;
  assign new_n10747_ = ~\b[14]  & ~new_n10746_;
  assign new_n10748_ = ~new_n10237_ & ~\quotient[26] ;
  assign new_n10749_ = ~new_n10247_ & new_n10400_;
  assign new_n10750_ = ~new_n10396_ & new_n10749_;
  assign new_n10751_ = ~new_n10397_ & ~new_n10400_;
  assign new_n10752_ = ~new_n10750_ & ~new_n10751_;
  assign new_n10753_ = new_n10530_ & ~new_n10752_;
  assign new_n10754_ = ~new_n10527_ & new_n10753_;
  assign new_n10755_ = ~new_n10748_ & ~new_n10754_;
  assign new_n10756_ = ~\b[13]  & ~new_n10755_;
  assign new_n10757_ = ~new_n10246_ & ~\quotient[26] ;
  assign new_n10758_ = ~new_n10256_ & new_n10395_;
  assign new_n10759_ = ~new_n10391_ & new_n10758_;
  assign new_n10760_ = ~new_n10392_ & ~new_n10395_;
  assign new_n10761_ = ~new_n10759_ & ~new_n10760_;
  assign new_n10762_ = new_n10530_ & ~new_n10761_;
  assign new_n10763_ = ~new_n10527_ & new_n10762_;
  assign new_n10764_ = ~new_n10757_ & ~new_n10763_;
  assign new_n10765_ = ~\b[12]  & ~new_n10764_;
  assign new_n10766_ = ~new_n10255_ & ~\quotient[26] ;
  assign new_n10767_ = ~new_n10265_ & new_n10390_;
  assign new_n10768_ = ~new_n10386_ & new_n10767_;
  assign new_n10769_ = ~new_n10387_ & ~new_n10390_;
  assign new_n10770_ = ~new_n10768_ & ~new_n10769_;
  assign new_n10771_ = new_n10530_ & ~new_n10770_;
  assign new_n10772_ = ~new_n10527_ & new_n10771_;
  assign new_n10773_ = ~new_n10766_ & ~new_n10772_;
  assign new_n10774_ = ~\b[11]  & ~new_n10773_;
  assign new_n10775_ = ~new_n10264_ & ~\quotient[26] ;
  assign new_n10776_ = ~new_n10274_ & new_n10385_;
  assign new_n10777_ = ~new_n10381_ & new_n10776_;
  assign new_n10778_ = ~new_n10382_ & ~new_n10385_;
  assign new_n10779_ = ~new_n10777_ & ~new_n10778_;
  assign new_n10780_ = new_n10530_ & ~new_n10779_;
  assign new_n10781_ = ~new_n10527_ & new_n10780_;
  assign new_n10782_ = ~new_n10775_ & ~new_n10781_;
  assign new_n10783_ = ~\b[10]  & ~new_n10782_;
  assign new_n10784_ = ~new_n10273_ & ~\quotient[26] ;
  assign new_n10785_ = ~new_n10283_ & new_n10380_;
  assign new_n10786_ = ~new_n10376_ & new_n10785_;
  assign new_n10787_ = ~new_n10377_ & ~new_n10380_;
  assign new_n10788_ = ~new_n10786_ & ~new_n10787_;
  assign new_n10789_ = new_n10530_ & ~new_n10788_;
  assign new_n10790_ = ~new_n10527_ & new_n10789_;
  assign new_n10791_ = ~new_n10784_ & ~new_n10790_;
  assign new_n10792_ = ~\b[9]  & ~new_n10791_;
  assign new_n10793_ = ~new_n10282_ & ~\quotient[26] ;
  assign new_n10794_ = ~new_n10292_ & new_n10375_;
  assign new_n10795_ = ~new_n10371_ & new_n10794_;
  assign new_n10796_ = ~new_n10372_ & ~new_n10375_;
  assign new_n10797_ = ~new_n10795_ & ~new_n10796_;
  assign new_n10798_ = new_n10530_ & ~new_n10797_;
  assign new_n10799_ = ~new_n10527_ & new_n10798_;
  assign new_n10800_ = ~new_n10793_ & ~new_n10799_;
  assign new_n10801_ = ~\b[8]  & ~new_n10800_;
  assign new_n10802_ = ~new_n10291_ & ~\quotient[26] ;
  assign new_n10803_ = ~new_n10301_ & new_n10370_;
  assign new_n10804_ = ~new_n10366_ & new_n10803_;
  assign new_n10805_ = ~new_n10367_ & ~new_n10370_;
  assign new_n10806_ = ~new_n10804_ & ~new_n10805_;
  assign new_n10807_ = new_n10530_ & ~new_n10806_;
  assign new_n10808_ = ~new_n10527_ & new_n10807_;
  assign new_n10809_ = ~new_n10802_ & ~new_n10808_;
  assign new_n10810_ = ~\b[7]  & ~new_n10809_;
  assign new_n10811_ = ~new_n10300_ & ~\quotient[26] ;
  assign new_n10812_ = ~new_n10310_ & new_n10365_;
  assign new_n10813_ = ~new_n10361_ & new_n10812_;
  assign new_n10814_ = ~new_n10362_ & ~new_n10365_;
  assign new_n10815_ = ~new_n10813_ & ~new_n10814_;
  assign new_n10816_ = new_n10530_ & ~new_n10815_;
  assign new_n10817_ = ~new_n10527_ & new_n10816_;
  assign new_n10818_ = ~new_n10811_ & ~new_n10817_;
  assign new_n10819_ = ~\b[6]  & ~new_n10818_;
  assign new_n10820_ = ~new_n10309_ & ~\quotient[26] ;
  assign new_n10821_ = ~new_n10319_ & new_n10360_;
  assign new_n10822_ = ~new_n10356_ & new_n10821_;
  assign new_n10823_ = ~new_n10357_ & ~new_n10360_;
  assign new_n10824_ = ~new_n10822_ & ~new_n10823_;
  assign new_n10825_ = new_n10530_ & ~new_n10824_;
  assign new_n10826_ = ~new_n10527_ & new_n10825_;
  assign new_n10827_ = ~new_n10820_ & ~new_n10826_;
  assign new_n10828_ = ~\b[5]  & ~new_n10827_;
  assign new_n10829_ = ~new_n10318_ & ~\quotient[26] ;
  assign new_n10830_ = ~new_n10327_ & new_n10355_;
  assign new_n10831_ = ~new_n10351_ & new_n10830_;
  assign new_n10832_ = ~new_n10352_ & ~new_n10355_;
  assign new_n10833_ = ~new_n10831_ & ~new_n10832_;
  assign new_n10834_ = new_n10530_ & ~new_n10833_;
  assign new_n10835_ = ~new_n10527_ & new_n10834_;
  assign new_n10836_ = ~new_n10829_ & ~new_n10835_;
  assign new_n10837_ = ~\b[4]  & ~new_n10836_;
  assign new_n10838_ = ~new_n10326_ & ~\quotient[26] ;
  assign new_n10839_ = ~new_n10346_ & new_n10350_;
  assign new_n10840_ = ~new_n10345_ & new_n10839_;
  assign new_n10841_ = ~new_n10347_ & ~new_n10350_;
  assign new_n10842_ = ~new_n10840_ & ~new_n10841_;
  assign new_n10843_ = new_n10530_ & ~new_n10842_;
  assign new_n10844_ = ~new_n10527_ & new_n10843_;
  assign new_n10845_ = ~new_n10838_ & ~new_n10844_;
  assign new_n10846_ = ~\b[3]  & ~new_n10845_;
  assign new_n10847_ = ~new_n10339_ & ~\quotient[26] ;
  assign new_n10848_ = ~new_n10342_ & new_n10344_;
  assign new_n10849_ = ~new_n10340_ & new_n10848_;
  assign new_n10850_ = new_n10530_ & ~new_n10849_;
  assign new_n10851_ = ~new_n10345_ & new_n10850_;
  assign new_n10852_ = ~new_n10527_ & new_n10851_;
  assign new_n10853_ = ~new_n10847_ & ~new_n10852_;
  assign new_n10854_ = ~\b[2]  & ~new_n10853_;
  assign new_n10855_ = \b[0]  & ~\b[38] ;
  assign new_n10856_ = new_n410_ & new_n10855_;
  assign new_n10857_ = new_n421_ & new_n10856_;
  assign new_n10858_ = new_n597_ & new_n10857_;
  assign new_n10859_ = new_n595_ & new_n10858_;
  assign new_n10860_ = ~new_n10527_ & new_n10859_;
  assign new_n10861_ = \a[26]  & ~new_n10860_;
  assign new_n10862_ = new_n293_ & new_n10344_;
  assign new_n10863_ = new_n291_ & new_n10862_;
  assign new_n10864_ = new_n302_ & new_n10863_;
  assign new_n10865_ = new_n288_ & new_n10864_;
  assign new_n10866_ = ~new_n10527_ & new_n10865_;
  assign new_n10867_ = ~new_n10861_ & ~new_n10866_;
  assign new_n10868_ = \b[1]  & ~new_n10867_;
  assign new_n10869_ = ~\b[1]  & ~new_n10866_;
  assign new_n10870_ = ~new_n10861_ & new_n10869_;
  assign new_n10871_ = ~new_n10868_ & ~new_n10870_;
  assign new_n10872_ = ~\a[25]  & \b[0] ;
  assign new_n10873_ = ~new_n10871_ & ~new_n10872_;
  assign new_n10874_ = ~\b[1]  & ~new_n10867_;
  assign new_n10875_ = ~new_n10873_ & ~new_n10874_;
  assign new_n10876_ = \b[2]  & ~new_n10852_;
  assign new_n10877_ = ~new_n10847_ & new_n10876_;
  assign new_n10878_ = ~new_n10854_ & ~new_n10877_;
  assign new_n10879_ = ~new_n10875_ & new_n10878_;
  assign new_n10880_ = ~new_n10854_ & ~new_n10879_;
  assign new_n10881_ = \b[3]  & ~new_n10844_;
  assign new_n10882_ = ~new_n10838_ & new_n10881_;
  assign new_n10883_ = ~new_n10846_ & ~new_n10882_;
  assign new_n10884_ = ~new_n10880_ & new_n10883_;
  assign new_n10885_ = ~new_n10846_ & ~new_n10884_;
  assign new_n10886_ = \b[4]  & ~new_n10835_;
  assign new_n10887_ = ~new_n10829_ & new_n10886_;
  assign new_n10888_ = ~new_n10837_ & ~new_n10887_;
  assign new_n10889_ = ~new_n10885_ & new_n10888_;
  assign new_n10890_ = ~new_n10837_ & ~new_n10889_;
  assign new_n10891_ = \b[5]  & ~new_n10826_;
  assign new_n10892_ = ~new_n10820_ & new_n10891_;
  assign new_n10893_ = ~new_n10828_ & ~new_n10892_;
  assign new_n10894_ = ~new_n10890_ & new_n10893_;
  assign new_n10895_ = ~new_n10828_ & ~new_n10894_;
  assign new_n10896_ = \b[6]  & ~new_n10817_;
  assign new_n10897_ = ~new_n10811_ & new_n10896_;
  assign new_n10898_ = ~new_n10819_ & ~new_n10897_;
  assign new_n10899_ = ~new_n10895_ & new_n10898_;
  assign new_n10900_ = ~new_n10819_ & ~new_n10899_;
  assign new_n10901_ = \b[7]  & ~new_n10808_;
  assign new_n10902_ = ~new_n10802_ & new_n10901_;
  assign new_n10903_ = ~new_n10810_ & ~new_n10902_;
  assign new_n10904_ = ~new_n10900_ & new_n10903_;
  assign new_n10905_ = ~new_n10810_ & ~new_n10904_;
  assign new_n10906_ = \b[8]  & ~new_n10799_;
  assign new_n10907_ = ~new_n10793_ & new_n10906_;
  assign new_n10908_ = ~new_n10801_ & ~new_n10907_;
  assign new_n10909_ = ~new_n10905_ & new_n10908_;
  assign new_n10910_ = ~new_n10801_ & ~new_n10909_;
  assign new_n10911_ = \b[9]  & ~new_n10790_;
  assign new_n10912_ = ~new_n10784_ & new_n10911_;
  assign new_n10913_ = ~new_n10792_ & ~new_n10912_;
  assign new_n10914_ = ~new_n10910_ & new_n10913_;
  assign new_n10915_ = ~new_n10792_ & ~new_n10914_;
  assign new_n10916_ = \b[10]  & ~new_n10781_;
  assign new_n10917_ = ~new_n10775_ & new_n10916_;
  assign new_n10918_ = ~new_n10783_ & ~new_n10917_;
  assign new_n10919_ = ~new_n10915_ & new_n10918_;
  assign new_n10920_ = ~new_n10783_ & ~new_n10919_;
  assign new_n10921_ = \b[11]  & ~new_n10772_;
  assign new_n10922_ = ~new_n10766_ & new_n10921_;
  assign new_n10923_ = ~new_n10774_ & ~new_n10922_;
  assign new_n10924_ = ~new_n10920_ & new_n10923_;
  assign new_n10925_ = ~new_n10774_ & ~new_n10924_;
  assign new_n10926_ = \b[12]  & ~new_n10763_;
  assign new_n10927_ = ~new_n10757_ & new_n10926_;
  assign new_n10928_ = ~new_n10765_ & ~new_n10927_;
  assign new_n10929_ = ~new_n10925_ & new_n10928_;
  assign new_n10930_ = ~new_n10765_ & ~new_n10929_;
  assign new_n10931_ = \b[13]  & ~new_n10754_;
  assign new_n10932_ = ~new_n10748_ & new_n10931_;
  assign new_n10933_ = ~new_n10756_ & ~new_n10932_;
  assign new_n10934_ = ~new_n10930_ & new_n10933_;
  assign new_n10935_ = ~new_n10756_ & ~new_n10934_;
  assign new_n10936_ = \b[14]  & ~new_n10745_;
  assign new_n10937_ = ~new_n10739_ & new_n10936_;
  assign new_n10938_ = ~new_n10747_ & ~new_n10937_;
  assign new_n10939_ = ~new_n10935_ & new_n10938_;
  assign new_n10940_ = ~new_n10747_ & ~new_n10939_;
  assign new_n10941_ = \b[15]  & ~new_n10736_;
  assign new_n10942_ = ~new_n10730_ & new_n10941_;
  assign new_n10943_ = ~new_n10738_ & ~new_n10942_;
  assign new_n10944_ = ~new_n10940_ & new_n10943_;
  assign new_n10945_ = ~new_n10738_ & ~new_n10944_;
  assign new_n10946_ = \b[16]  & ~new_n10727_;
  assign new_n10947_ = ~new_n10721_ & new_n10946_;
  assign new_n10948_ = ~new_n10729_ & ~new_n10947_;
  assign new_n10949_ = ~new_n10945_ & new_n10948_;
  assign new_n10950_ = ~new_n10729_ & ~new_n10949_;
  assign new_n10951_ = \b[17]  & ~new_n10718_;
  assign new_n10952_ = ~new_n10712_ & new_n10951_;
  assign new_n10953_ = ~new_n10720_ & ~new_n10952_;
  assign new_n10954_ = ~new_n10950_ & new_n10953_;
  assign new_n10955_ = ~new_n10720_ & ~new_n10954_;
  assign new_n10956_ = \b[18]  & ~new_n10709_;
  assign new_n10957_ = ~new_n10703_ & new_n10956_;
  assign new_n10958_ = ~new_n10711_ & ~new_n10957_;
  assign new_n10959_ = ~new_n10955_ & new_n10958_;
  assign new_n10960_ = ~new_n10711_ & ~new_n10959_;
  assign new_n10961_ = \b[19]  & ~new_n10700_;
  assign new_n10962_ = ~new_n10694_ & new_n10961_;
  assign new_n10963_ = ~new_n10702_ & ~new_n10962_;
  assign new_n10964_ = ~new_n10960_ & new_n10963_;
  assign new_n10965_ = ~new_n10702_ & ~new_n10964_;
  assign new_n10966_ = \b[20]  & ~new_n10691_;
  assign new_n10967_ = ~new_n10685_ & new_n10966_;
  assign new_n10968_ = ~new_n10693_ & ~new_n10967_;
  assign new_n10969_ = ~new_n10965_ & new_n10968_;
  assign new_n10970_ = ~new_n10693_ & ~new_n10969_;
  assign new_n10971_ = \b[21]  & ~new_n10682_;
  assign new_n10972_ = ~new_n10676_ & new_n10971_;
  assign new_n10973_ = ~new_n10684_ & ~new_n10972_;
  assign new_n10974_ = ~new_n10970_ & new_n10973_;
  assign new_n10975_ = ~new_n10684_ & ~new_n10974_;
  assign new_n10976_ = \b[22]  & ~new_n10673_;
  assign new_n10977_ = ~new_n10667_ & new_n10976_;
  assign new_n10978_ = ~new_n10675_ & ~new_n10977_;
  assign new_n10979_ = ~new_n10975_ & new_n10978_;
  assign new_n10980_ = ~new_n10675_ & ~new_n10979_;
  assign new_n10981_ = \b[23]  & ~new_n10664_;
  assign new_n10982_ = ~new_n10658_ & new_n10981_;
  assign new_n10983_ = ~new_n10666_ & ~new_n10982_;
  assign new_n10984_ = ~new_n10980_ & new_n10983_;
  assign new_n10985_ = ~new_n10666_ & ~new_n10984_;
  assign new_n10986_ = \b[24]  & ~new_n10655_;
  assign new_n10987_ = ~new_n10649_ & new_n10986_;
  assign new_n10988_ = ~new_n10657_ & ~new_n10987_;
  assign new_n10989_ = ~new_n10985_ & new_n10988_;
  assign new_n10990_ = ~new_n10657_ & ~new_n10989_;
  assign new_n10991_ = \b[25]  & ~new_n10646_;
  assign new_n10992_ = ~new_n10640_ & new_n10991_;
  assign new_n10993_ = ~new_n10648_ & ~new_n10992_;
  assign new_n10994_ = ~new_n10990_ & new_n10993_;
  assign new_n10995_ = ~new_n10648_ & ~new_n10994_;
  assign new_n10996_ = \b[26]  & ~new_n10637_;
  assign new_n10997_ = ~new_n10631_ & new_n10996_;
  assign new_n10998_ = ~new_n10639_ & ~new_n10997_;
  assign new_n10999_ = ~new_n10995_ & new_n10998_;
  assign new_n11000_ = ~new_n10639_ & ~new_n10999_;
  assign new_n11001_ = \b[27]  & ~new_n10628_;
  assign new_n11002_ = ~new_n10622_ & new_n11001_;
  assign new_n11003_ = ~new_n10630_ & ~new_n11002_;
  assign new_n11004_ = ~new_n11000_ & new_n11003_;
  assign new_n11005_ = ~new_n10630_ & ~new_n11004_;
  assign new_n11006_ = \b[28]  & ~new_n10619_;
  assign new_n11007_ = ~new_n10613_ & new_n11006_;
  assign new_n11008_ = ~new_n10621_ & ~new_n11007_;
  assign new_n11009_ = ~new_n11005_ & new_n11008_;
  assign new_n11010_ = ~new_n10621_ & ~new_n11009_;
  assign new_n11011_ = \b[29]  & ~new_n10610_;
  assign new_n11012_ = ~new_n10604_ & new_n11011_;
  assign new_n11013_ = ~new_n10612_ & ~new_n11012_;
  assign new_n11014_ = ~new_n11010_ & new_n11013_;
  assign new_n11015_ = ~new_n10612_ & ~new_n11014_;
  assign new_n11016_ = \b[30]  & ~new_n10601_;
  assign new_n11017_ = ~new_n10595_ & new_n11016_;
  assign new_n11018_ = ~new_n10603_ & ~new_n11017_;
  assign new_n11019_ = ~new_n11015_ & new_n11018_;
  assign new_n11020_ = ~new_n10603_ & ~new_n11019_;
  assign new_n11021_ = \b[31]  & ~new_n10592_;
  assign new_n11022_ = ~new_n10586_ & new_n11021_;
  assign new_n11023_ = ~new_n10594_ & ~new_n11022_;
  assign new_n11024_ = ~new_n11020_ & new_n11023_;
  assign new_n11025_ = ~new_n10594_ & ~new_n11024_;
  assign new_n11026_ = \b[32]  & ~new_n10583_;
  assign new_n11027_ = ~new_n10577_ & new_n11026_;
  assign new_n11028_ = ~new_n10585_ & ~new_n11027_;
  assign new_n11029_ = ~new_n11025_ & new_n11028_;
  assign new_n11030_ = ~new_n10585_ & ~new_n11029_;
  assign new_n11031_ = \b[33]  & ~new_n10574_;
  assign new_n11032_ = ~new_n10568_ & new_n11031_;
  assign new_n11033_ = ~new_n10576_ & ~new_n11032_;
  assign new_n11034_ = ~new_n11030_ & new_n11033_;
  assign new_n11035_ = ~new_n10576_ & ~new_n11034_;
  assign new_n11036_ = \b[34]  & ~new_n10565_;
  assign new_n11037_ = ~new_n10559_ & new_n11036_;
  assign new_n11038_ = ~new_n10567_ & ~new_n11037_;
  assign new_n11039_ = ~new_n11035_ & new_n11038_;
  assign new_n11040_ = ~new_n10567_ & ~new_n11039_;
  assign new_n11041_ = \b[35]  & ~new_n10556_;
  assign new_n11042_ = ~new_n10550_ & new_n11041_;
  assign new_n11043_ = ~new_n10558_ & ~new_n11042_;
  assign new_n11044_ = ~new_n11040_ & new_n11043_;
  assign new_n11045_ = ~new_n10558_ & ~new_n11044_;
  assign new_n11046_ = \b[36]  & ~new_n10547_;
  assign new_n11047_ = ~new_n10541_ & new_n11046_;
  assign new_n11048_ = ~new_n10549_ & ~new_n11047_;
  assign new_n11049_ = ~new_n11045_ & new_n11048_;
  assign new_n11050_ = ~new_n10549_ & ~new_n11049_;
  assign new_n11051_ = \b[37]  & ~new_n10538_;
  assign new_n11052_ = ~new_n10532_ & new_n11051_;
  assign new_n11053_ = ~new_n10540_ & ~new_n11052_;
  assign new_n11054_ = ~new_n11050_ & new_n11053_;
  assign new_n11055_ = ~new_n10540_ & ~new_n11054_;
  assign new_n11056_ = ~new_n10020_ & ~\quotient[26] ;
  assign new_n11057_ = ~new_n10022_ & new_n10525_;
  assign new_n11058_ = ~new_n10521_ & new_n11057_;
  assign new_n11059_ = ~new_n10522_ & ~new_n10525_;
  assign new_n11060_ = ~new_n11058_ & ~new_n11059_;
  assign new_n11061_ = \quotient[26]  & ~new_n11060_;
  assign new_n11062_ = ~new_n11056_ & ~new_n11061_;
  assign new_n11063_ = ~\b[38]  & ~new_n11062_;
  assign new_n11064_ = \b[38]  & ~new_n11056_;
  assign new_n11065_ = ~new_n11061_ & new_n11064_;
  assign new_n11066_ = new_n410_ & new_n421_;
  assign new_n11067_ = new_n597_ & new_n11066_;
  assign new_n11068_ = new_n595_ & new_n11067_;
  assign new_n11069_ = ~new_n11065_ & new_n11068_;
  assign new_n11070_ = ~new_n11063_ & new_n11069_;
  assign new_n11071_ = ~new_n11055_ & new_n11070_;
  assign new_n11072_ = new_n10530_ & ~new_n11062_;
  assign \quotient[25]  = new_n11071_ | new_n11072_;
  assign new_n11074_ = ~new_n10549_ & new_n11053_;
  assign new_n11075_ = ~new_n11049_ & new_n11074_;
  assign new_n11076_ = ~new_n11050_ & ~new_n11053_;
  assign new_n11077_ = ~new_n11075_ & ~new_n11076_;
  assign new_n11078_ = \quotient[25]  & ~new_n11077_;
  assign new_n11079_ = ~new_n10539_ & ~new_n11072_;
  assign new_n11080_ = ~new_n11071_ & new_n11079_;
  assign new_n11081_ = ~new_n11078_ & ~new_n11080_;
  assign new_n11082_ = ~new_n10540_ & ~new_n11065_;
  assign new_n11083_ = ~new_n11063_ & new_n11082_;
  assign new_n11084_ = ~new_n11054_ & new_n11083_;
  assign new_n11085_ = ~new_n11063_ & ~new_n11065_;
  assign new_n11086_ = ~new_n11055_ & ~new_n11085_;
  assign new_n11087_ = ~new_n11084_ & ~new_n11086_;
  assign new_n11088_ = \quotient[25]  & ~new_n11087_;
  assign new_n11089_ = ~new_n11062_ & ~new_n11072_;
  assign new_n11090_ = ~new_n11071_ & new_n11089_;
  assign new_n11091_ = ~new_n11088_ & ~new_n11090_;
  assign new_n11092_ = ~\b[39]  & ~new_n11091_;
  assign new_n11093_ = ~\b[38]  & ~new_n11081_;
  assign new_n11094_ = ~new_n10558_ & new_n11048_;
  assign new_n11095_ = ~new_n11044_ & new_n11094_;
  assign new_n11096_ = ~new_n11045_ & ~new_n11048_;
  assign new_n11097_ = ~new_n11095_ & ~new_n11096_;
  assign new_n11098_ = \quotient[25]  & ~new_n11097_;
  assign new_n11099_ = ~new_n10548_ & ~new_n11072_;
  assign new_n11100_ = ~new_n11071_ & new_n11099_;
  assign new_n11101_ = ~new_n11098_ & ~new_n11100_;
  assign new_n11102_ = ~\b[37]  & ~new_n11101_;
  assign new_n11103_ = ~new_n10567_ & new_n11043_;
  assign new_n11104_ = ~new_n11039_ & new_n11103_;
  assign new_n11105_ = ~new_n11040_ & ~new_n11043_;
  assign new_n11106_ = ~new_n11104_ & ~new_n11105_;
  assign new_n11107_ = \quotient[25]  & ~new_n11106_;
  assign new_n11108_ = ~new_n10557_ & ~new_n11072_;
  assign new_n11109_ = ~new_n11071_ & new_n11108_;
  assign new_n11110_ = ~new_n11107_ & ~new_n11109_;
  assign new_n11111_ = ~\b[36]  & ~new_n11110_;
  assign new_n11112_ = ~new_n10576_ & new_n11038_;
  assign new_n11113_ = ~new_n11034_ & new_n11112_;
  assign new_n11114_ = ~new_n11035_ & ~new_n11038_;
  assign new_n11115_ = ~new_n11113_ & ~new_n11114_;
  assign new_n11116_ = \quotient[25]  & ~new_n11115_;
  assign new_n11117_ = ~new_n10566_ & ~new_n11072_;
  assign new_n11118_ = ~new_n11071_ & new_n11117_;
  assign new_n11119_ = ~new_n11116_ & ~new_n11118_;
  assign new_n11120_ = ~\b[35]  & ~new_n11119_;
  assign new_n11121_ = ~new_n10585_ & new_n11033_;
  assign new_n11122_ = ~new_n11029_ & new_n11121_;
  assign new_n11123_ = ~new_n11030_ & ~new_n11033_;
  assign new_n11124_ = ~new_n11122_ & ~new_n11123_;
  assign new_n11125_ = \quotient[25]  & ~new_n11124_;
  assign new_n11126_ = ~new_n10575_ & ~new_n11072_;
  assign new_n11127_ = ~new_n11071_ & new_n11126_;
  assign new_n11128_ = ~new_n11125_ & ~new_n11127_;
  assign new_n11129_ = ~\b[34]  & ~new_n11128_;
  assign new_n11130_ = ~new_n10594_ & new_n11028_;
  assign new_n11131_ = ~new_n11024_ & new_n11130_;
  assign new_n11132_ = ~new_n11025_ & ~new_n11028_;
  assign new_n11133_ = ~new_n11131_ & ~new_n11132_;
  assign new_n11134_ = \quotient[25]  & ~new_n11133_;
  assign new_n11135_ = ~new_n10584_ & ~new_n11072_;
  assign new_n11136_ = ~new_n11071_ & new_n11135_;
  assign new_n11137_ = ~new_n11134_ & ~new_n11136_;
  assign new_n11138_ = ~\b[33]  & ~new_n11137_;
  assign new_n11139_ = ~new_n10603_ & new_n11023_;
  assign new_n11140_ = ~new_n11019_ & new_n11139_;
  assign new_n11141_ = ~new_n11020_ & ~new_n11023_;
  assign new_n11142_ = ~new_n11140_ & ~new_n11141_;
  assign new_n11143_ = \quotient[25]  & ~new_n11142_;
  assign new_n11144_ = ~new_n10593_ & ~new_n11072_;
  assign new_n11145_ = ~new_n11071_ & new_n11144_;
  assign new_n11146_ = ~new_n11143_ & ~new_n11145_;
  assign new_n11147_ = ~\b[32]  & ~new_n11146_;
  assign new_n11148_ = ~new_n10612_ & new_n11018_;
  assign new_n11149_ = ~new_n11014_ & new_n11148_;
  assign new_n11150_ = ~new_n11015_ & ~new_n11018_;
  assign new_n11151_ = ~new_n11149_ & ~new_n11150_;
  assign new_n11152_ = \quotient[25]  & ~new_n11151_;
  assign new_n11153_ = ~new_n10602_ & ~new_n11072_;
  assign new_n11154_ = ~new_n11071_ & new_n11153_;
  assign new_n11155_ = ~new_n11152_ & ~new_n11154_;
  assign new_n11156_ = ~\b[31]  & ~new_n11155_;
  assign new_n11157_ = ~new_n10621_ & new_n11013_;
  assign new_n11158_ = ~new_n11009_ & new_n11157_;
  assign new_n11159_ = ~new_n11010_ & ~new_n11013_;
  assign new_n11160_ = ~new_n11158_ & ~new_n11159_;
  assign new_n11161_ = \quotient[25]  & ~new_n11160_;
  assign new_n11162_ = ~new_n10611_ & ~new_n11072_;
  assign new_n11163_ = ~new_n11071_ & new_n11162_;
  assign new_n11164_ = ~new_n11161_ & ~new_n11163_;
  assign new_n11165_ = ~\b[30]  & ~new_n11164_;
  assign new_n11166_ = ~new_n10630_ & new_n11008_;
  assign new_n11167_ = ~new_n11004_ & new_n11166_;
  assign new_n11168_ = ~new_n11005_ & ~new_n11008_;
  assign new_n11169_ = ~new_n11167_ & ~new_n11168_;
  assign new_n11170_ = \quotient[25]  & ~new_n11169_;
  assign new_n11171_ = ~new_n10620_ & ~new_n11072_;
  assign new_n11172_ = ~new_n11071_ & new_n11171_;
  assign new_n11173_ = ~new_n11170_ & ~new_n11172_;
  assign new_n11174_ = ~\b[29]  & ~new_n11173_;
  assign new_n11175_ = ~new_n10639_ & new_n11003_;
  assign new_n11176_ = ~new_n10999_ & new_n11175_;
  assign new_n11177_ = ~new_n11000_ & ~new_n11003_;
  assign new_n11178_ = ~new_n11176_ & ~new_n11177_;
  assign new_n11179_ = \quotient[25]  & ~new_n11178_;
  assign new_n11180_ = ~new_n10629_ & ~new_n11072_;
  assign new_n11181_ = ~new_n11071_ & new_n11180_;
  assign new_n11182_ = ~new_n11179_ & ~new_n11181_;
  assign new_n11183_ = ~\b[28]  & ~new_n11182_;
  assign new_n11184_ = ~new_n10648_ & new_n10998_;
  assign new_n11185_ = ~new_n10994_ & new_n11184_;
  assign new_n11186_ = ~new_n10995_ & ~new_n10998_;
  assign new_n11187_ = ~new_n11185_ & ~new_n11186_;
  assign new_n11188_ = \quotient[25]  & ~new_n11187_;
  assign new_n11189_ = ~new_n10638_ & ~new_n11072_;
  assign new_n11190_ = ~new_n11071_ & new_n11189_;
  assign new_n11191_ = ~new_n11188_ & ~new_n11190_;
  assign new_n11192_ = ~\b[27]  & ~new_n11191_;
  assign new_n11193_ = ~new_n10657_ & new_n10993_;
  assign new_n11194_ = ~new_n10989_ & new_n11193_;
  assign new_n11195_ = ~new_n10990_ & ~new_n10993_;
  assign new_n11196_ = ~new_n11194_ & ~new_n11195_;
  assign new_n11197_ = \quotient[25]  & ~new_n11196_;
  assign new_n11198_ = ~new_n10647_ & ~new_n11072_;
  assign new_n11199_ = ~new_n11071_ & new_n11198_;
  assign new_n11200_ = ~new_n11197_ & ~new_n11199_;
  assign new_n11201_ = ~\b[26]  & ~new_n11200_;
  assign new_n11202_ = ~new_n10666_ & new_n10988_;
  assign new_n11203_ = ~new_n10984_ & new_n11202_;
  assign new_n11204_ = ~new_n10985_ & ~new_n10988_;
  assign new_n11205_ = ~new_n11203_ & ~new_n11204_;
  assign new_n11206_ = \quotient[25]  & ~new_n11205_;
  assign new_n11207_ = ~new_n10656_ & ~new_n11072_;
  assign new_n11208_ = ~new_n11071_ & new_n11207_;
  assign new_n11209_ = ~new_n11206_ & ~new_n11208_;
  assign new_n11210_ = ~\b[25]  & ~new_n11209_;
  assign new_n11211_ = ~new_n10675_ & new_n10983_;
  assign new_n11212_ = ~new_n10979_ & new_n11211_;
  assign new_n11213_ = ~new_n10980_ & ~new_n10983_;
  assign new_n11214_ = ~new_n11212_ & ~new_n11213_;
  assign new_n11215_ = \quotient[25]  & ~new_n11214_;
  assign new_n11216_ = ~new_n10665_ & ~new_n11072_;
  assign new_n11217_ = ~new_n11071_ & new_n11216_;
  assign new_n11218_ = ~new_n11215_ & ~new_n11217_;
  assign new_n11219_ = ~\b[24]  & ~new_n11218_;
  assign new_n11220_ = ~new_n10684_ & new_n10978_;
  assign new_n11221_ = ~new_n10974_ & new_n11220_;
  assign new_n11222_ = ~new_n10975_ & ~new_n10978_;
  assign new_n11223_ = ~new_n11221_ & ~new_n11222_;
  assign new_n11224_ = \quotient[25]  & ~new_n11223_;
  assign new_n11225_ = ~new_n10674_ & ~new_n11072_;
  assign new_n11226_ = ~new_n11071_ & new_n11225_;
  assign new_n11227_ = ~new_n11224_ & ~new_n11226_;
  assign new_n11228_ = ~\b[23]  & ~new_n11227_;
  assign new_n11229_ = ~new_n10693_ & new_n10973_;
  assign new_n11230_ = ~new_n10969_ & new_n11229_;
  assign new_n11231_ = ~new_n10970_ & ~new_n10973_;
  assign new_n11232_ = ~new_n11230_ & ~new_n11231_;
  assign new_n11233_ = \quotient[25]  & ~new_n11232_;
  assign new_n11234_ = ~new_n10683_ & ~new_n11072_;
  assign new_n11235_ = ~new_n11071_ & new_n11234_;
  assign new_n11236_ = ~new_n11233_ & ~new_n11235_;
  assign new_n11237_ = ~\b[22]  & ~new_n11236_;
  assign new_n11238_ = ~new_n10702_ & new_n10968_;
  assign new_n11239_ = ~new_n10964_ & new_n11238_;
  assign new_n11240_ = ~new_n10965_ & ~new_n10968_;
  assign new_n11241_ = ~new_n11239_ & ~new_n11240_;
  assign new_n11242_ = \quotient[25]  & ~new_n11241_;
  assign new_n11243_ = ~new_n10692_ & ~new_n11072_;
  assign new_n11244_ = ~new_n11071_ & new_n11243_;
  assign new_n11245_ = ~new_n11242_ & ~new_n11244_;
  assign new_n11246_ = ~\b[21]  & ~new_n11245_;
  assign new_n11247_ = ~new_n10711_ & new_n10963_;
  assign new_n11248_ = ~new_n10959_ & new_n11247_;
  assign new_n11249_ = ~new_n10960_ & ~new_n10963_;
  assign new_n11250_ = ~new_n11248_ & ~new_n11249_;
  assign new_n11251_ = \quotient[25]  & ~new_n11250_;
  assign new_n11252_ = ~new_n10701_ & ~new_n11072_;
  assign new_n11253_ = ~new_n11071_ & new_n11252_;
  assign new_n11254_ = ~new_n11251_ & ~new_n11253_;
  assign new_n11255_ = ~\b[20]  & ~new_n11254_;
  assign new_n11256_ = ~new_n10720_ & new_n10958_;
  assign new_n11257_ = ~new_n10954_ & new_n11256_;
  assign new_n11258_ = ~new_n10955_ & ~new_n10958_;
  assign new_n11259_ = ~new_n11257_ & ~new_n11258_;
  assign new_n11260_ = \quotient[25]  & ~new_n11259_;
  assign new_n11261_ = ~new_n10710_ & ~new_n11072_;
  assign new_n11262_ = ~new_n11071_ & new_n11261_;
  assign new_n11263_ = ~new_n11260_ & ~new_n11262_;
  assign new_n11264_ = ~\b[19]  & ~new_n11263_;
  assign new_n11265_ = ~new_n10729_ & new_n10953_;
  assign new_n11266_ = ~new_n10949_ & new_n11265_;
  assign new_n11267_ = ~new_n10950_ & ~new_n10953_;
  assign new_n11268_ = ~new_n11266_ & ~new_n11267_;
  assign new_n11269_ = \quotient[25]  & ~new_n11268_;
  assign new_n11270_ = ~new_n10719_ & ~new_n11072_;
  assign new_n11271_ = ~new_n11071_ & new_n11270_;
  assign new_n11272_ = ~new_n11269_ & ~new_n11271_;
  assign new_n11273_ = ~\b[18]  & ~new_n11272_;
  assign new_n11274_ = ~new_n10738_ & new_n10948_;
  assign new_n11275_ = ~new_n10944_ & new_n11274_;
  assign new_n11276_ = ~new_n10945_ & ~new_n10948_;
  assign new_n11277_ = ~new_n11275_ & ~new_n11276_;
  assign new_n11278_ = \quotient[25]  & ~new_n11277_;
  assign new_n11279_ = ~new_n10728_ & ~new_n11072_;
  assign new_n11280_ = ~new_n11071_ & new_n11279_;
  assign new_n11281_ = ~new_n11278_ & ~new_n11280_;
  assign new_n11282_ = ~\b[17]  & ~new_n11281_;
  assign new_n11283_ = ~new_n10747_ & new_n10943_;
  assign new_n11284_ = ~new_n10939_ & new_n11283_;
  assign new_n11285_ = ~new_n10940_ & ~new_n10943_;
  assign new_n11286_ = ~new_n11284_ & ~new_n11285_;
  assign new_n11287_ = \quotient[25]  & ~new_n11286_;
  assign new_n11288_ = ~new_n10737_ & ~new_n11072_;
  assign new_n11289_ = ~new_n11071_ & new_n11288_;
  assign new_n11290_ = ~new_n11287_ & ~new_n11289_;
  assign new_n11291_ = ~\b[16]  & ~new_n11290_;
  assign new_n11292_ = ~new_n10756_ & new_n10938_;
  assign new_n11293_ = ~new_n10934_ & new_n11292_;
  assign new_n11294_ = ~new_n10935_ & ~new_n10938_;
  assign new_n11295_ = ~new_n11293_ & ~new_n11294_;
  assign new_n11296_ = \quotient[25]  & ~new_n11295_;
  assign new_n11297_ = ~new_n10746_ & ~new_n11072_;
  assign new_n11298_ = ~new_n11071_ & new_n11297_;
  assign new_n11299_ = ~new_n11296_ & ~new_n11298_;
  assign new_n11300_ = ~\b[15]  & ~new_n11299_;
  assign new_n11301_ = ~new_n10765_ & new_n10933_;
  assign new_n11302_ = ~new_n10929_ & new_n11301_;
  assign new_n11303_ = ~new_n10930_ & ~new_n10933_;
  assign new_n11304_ = ~new_n11302_ & ~new_n11303_;
  assign new_n11305_ = \quotient[25]  & ~new_n11304_;
  assign new_n11306_ = ~new_n10755_ & ~new_n11072_;
  assign new_n11307_ = ~new_n11071_ & new_n11306_;
  assign new_n11308_ = ~new_n11305_ & ~new_n11307_;
  assign new_n11309_ = ~\b[14]  & ~new_n11308_;
  assign new_n11310_ = ~new_n10774_ & new_n10928_;
  assign new_n11311_ = ~new_n10924_ & new_n11310_;
  assign new_n11312_ = ~new_n10925_ & ~new_n10928_;
  assign new_n11313_ = ~new_n11311_ & ~new_n11312_;
  assign new_n11314_ = \quotient[25]  & ~new_n11313_;
  assign new_n11315_ = ~new_n10764_ & ~new_n11072_;
  assign new_n11316_ = ~new_n11071_ & new_n11315_;
  assign new_n11317_ = ~new_n11314_ & ~new_n11316_;
  assign new_n11318_ = ~\b[13]  & ~new_n11317_;
  assign new_n11319_ = ~new_n10783_ & new_n10923_;
  assign new_n11320_ = ~new_n10919_ & new_n11319_;
  assign new_n11321_ = ~new_n10920_ & ~new_n10923_;
  assign new_n11322_ = ~new_n11320_ & ~new_n11321_;
  assign new_n11323_ = \quotient[25]  & ~new_n11322_;
  assign new_n11324_ = ~new_n10773_ & ~new_n11072_;
  assign new_n11325_ = ~new_n11071_ & new_n11324_;
  assign new_n11326_ = ~new_n11323_ & ~new_n11325_;
  assign new_n11327_ = ~\b[12]  & ~new_n11326_;
  assign new_n11328_ = ~new_n10792_ & new_n10918_;
  assign new_n11329_ = ~new_n10914_ & new_n11328_;
  assign new_n11330_ = ~new_n10915_ & ~new_n10918_;
  assign new_n11331_ = ~new_n11329_ & ~new_n11330_;
  assign new_n11332_ = \quotient[25]  & ~new_n11331_;
  assign new_n11333_ = ~new_n10782_ & ~new_n11072_;
  assign new_n11334_ = ~new_n11071_ & new_n11333_;
  assign new_n11335_ = ~new_n11332_ & ~new_n11334_;
  assign new_n11336_ = ~\b[11]  & ~new_n11335_;
  assign new_n11337_ = ~new_n10801_ & new_n10913_;
  assign new_n11338_ = ~new_n10909_ & new_n11337_;
  assign new_n11339_ = ~new_n10910_ & ~new_n10913_;
  assign new_n11340_ = ~new_n11338_ & ~new_n11339_;
  assign new_n11341_ = \quotient[25]  & ~new_n11340_;
  assign new_n11342_ = ~new_n10791_ & ~new_n11072_;
  assign new_n11343_ = ~new_n11071_ & new_n11342_;
  assign new_n11344_ = ~new_n11341_ & ~new_n11343_;
  assign new_n11345_ = ~\b[10]  & ~new_n11344_;
  assign new_n11346_ = ~new_n10810_ & new_n10908_;
  assign new_n11347_ = ~new_n10904_ & new_n11346_;
  assign new_n11348_ = ~new_n10905_ & ~new_n10908_;
  assign new_n11349_ = ~new_n11347_ & ~new_n11348_;
  assign new_n11350_ = \quotient[25]  & ~new_n11349_;
  assign new_n11351_ = ~new_n10800_ & ~new_n11072_;
  assign new_n11352_ = ~new_n11071_ & new_n11351_;
  assign new_n11353_ = ~new_n11350_ & ~new_n11352_;
  assign new_n11354_ = ~\b[9]  & ~new_n11353_;
  assign new_n11355_ = ~new_n10819_ & new_n10903_;
  assign new_n11356_ = ~new_n10899_ & new_n11355_;
  assign new_n11357_ = ~new_n10900_ & ~new_n10903_;
  assign new_n11358_ = ~new_n11356_ & ~new_n11357_;
  assign new_n11359_ = \quotient[25]  & ~new_n11358_;
  assign new_n11360_ = ~new_n10809_ & ~new_n11072_;
  assign new_n11361_ = ~new_n11071_ & new_n11360_;
  assign new_n11362_ = ~new_n11359_ & ~new_n11361_;
  assign new_n11363_ = ~\b[8]  & ~new_n11362_;
  assign new_n11364_ = ~new_n10828_ & new_n10898_;
  assign new_n11365_ = ~new_n10894_ & new_n11364_;
  assign new_n11366_ = ~new_n10895_ & ~new_n10898_;
  assign new_n11367_ = ~new_n11365_ & ~new_n11366_;
  assign new_n11368_ = \quotient[25]  & ~new_n11367_;
  assign new_n11369_ = ~new_n10818_ & ~new_n11072_;
  assign new_n11370_ = ~new_n11071_ & new_n11369_;
  assign new_n11371_ = ~new_n11368_ & ~new_n11370_;
  assign new_n11372_ = ~\b[7]  & ~new_n11371_;
  assign new_n11373_ = ~new_n10837_ & new_n10893_;
  assign new_n11374_ = ~new_n10889_ & new_n11373_;
  assign new_n11375_ = ~new_n10890_ & ~new_n10893_;
  assign new_n11376_ = ~new_n11374_ & ~new_n11375_;
  assign new_n11377_ = \quotient[25]  & ~new_n11376_;
  assign new_n11378_ = ~new_n10827_ & ~new_n11072_;
  assign new_n11379_ = ~new_n11071_ & new_n11378_;
  assign new_n11380_ = ~new_n11377_ & ~new_n11379_;
  assign new_n11381_ = ~\b[6]  & ~new_n11380_;
  assign new_n11382_ = ~new_n10846_ & new_n10888_;
  assign new_n11383_ = ~new_n10884_ & new_n11382_;
  assign new_n11384_ = ~new_n10885_ & ~new_n10888_;
  assign new_n11385_ = ~new_n11383_ & ~new_n11384_;
  assign new_n11386_ = \quotient[25]  & ~new_n11385_;
  assign new_n11387_ = ~new_n10836_ & ~new_n11072_;
  assign new_n11388_ = ~new_n11071_ & new_n11387_;
  assign new_n11389_ = ~new_n11386_ & ~new_n11388_;
  assign new_n11390_ = ~\b[5]  & ~new_n11389_;
  assign new_n11391_ = ~new_n10854_ & new_n10883_;
  assign new_n11392_ = ~new_n10879_ & new_n11391_;
  assign new_n11393_ = ~new_n10880_ & ~new_n10883_;
  assign new_n11394_ = ~new_n11392_ & ~new_n11393_;
  assign new_n11395_ = \quotient[25]  & ~new_n11394_;
  assign new_n11396_ = ~new_n10845_ & ~new_n11072_;
  assign new_n11397_ = ~new_n11071_ & new_n11396_;
  assign new_n11398_ = ~new_n11395_ & ~new_n11397_;
  assign new_n11399_ = ~\b[4]  & ~new_n11398_;
  assign new_n11400_ = ~new_n10874_ & new_n10878_;
  assign new_n11401_ = ~new_n10873_ & new_n11400_;
  assign new_n11402_ = ~new_n10875_ & ~new_n10878_;
  assign new_n11403_ = ~new_n11401_ & ~new_n11402_;
  assign new_n11404_ = \quotient[25]  & ~new_n11403_;
  assign new_n11405_ = ~new_n10853_ & ~new_n11072_;
  assign new_n11406_ = ~new_n11071_ & new_n11405_;
  assign new_n11407_ = ~new_n11404_ & ~new_n11406_;
  assign new_n11408_ = ~\b[3]  & ~new_n11407_;
  assign new_n11409_ = ~new_n10870_ & new_n10872_;
  assign new_n11410_ = ~new_n10868_ & new_n11409_;
  assign new_n11411_ = ~new_n10873_ & ~new_n11410_;
  assign new_n11412_ = \quotient[25]  & new_n11411_;
  assign new_n11413_ = ~new_n10867_ & ~new_n11072_;
  assign new_n11414_ = ~new_n11071_ & new_n11413_;
  assign new_n11415_ = ~new_n11412_ & ~new_n11414_;
  assign new_n11416_ = ~\b[2]  & ~new_n11415_;
  assign new_n11417_ = \b[0]  & \quotient[25] ;
  assign new_n11418_ = \a[25]  & ~new_n11417_;
  assign new_n11419_ = new_n10872_ & \quotient[25] ;
  assign new_n11420_ = ~new_n11418_ & ~new_n11419_;
  assign new_n11421_ = \b[1]  & ~new_n11420_;
  assign new_n11422_ = ~\b[1]  & ~new_n11419_;
  assign new_n11423_ = ~new_n11418_ & new_n11422_;
  assign new_n11424_ = ~new_n11421_ & ~new_n11423_;
  assign new_n11425_ = ~\a[24]  & \b[0] ;
  assign new_n11426_ = ~new_n11424_ & ~new_n11425_;
  assign new_n11427_ = ~\b[1]  & ~new_n11420_;
  assign new_n11428_ = ~new_n11426_ & ~new_n11427_;
  assign new_n11429_ = \b[2]  & ~new_n11414_;
  assign new_n11430_ = ~new_n11412_ & new_n11429_;
  assign new_n11431_ = ~new_n11416_ & ~new_n11430_;
  assign new_n11432_ = ~new_n11428_ & new_n11431_;
  assign new_n11433_ = ~new_n11416_ & ~new_n11432_;
  assign new_n11434_ = \b[3]  & ~new_n11406_;
  assign new_n11435_ = ~new_n11404_ & new_n11434_;
  assign new_n11436_ = ~new_n11408_ & ~new_n11435_;
  assign new_n11437_ = ~new_n11433_ & new_n11436_;
  assign new_n11438_ = ~new_n11408_ & ~new_n11437_;
  assign new_n11439_ = \b[4]  & ~new_n11397_;
  assign new_n11440_ = ~new_n11395_ & new_n11439_;
  assign new_n11441_ = ~new_n11399_ & ~new_n11440_;
  assign new_n11442_ = ~new_n11438_ & new_n11441_;
  assign new_n11443_ = ~new_n11399_ & ~new_n11442_;
  assign new_n11444_ = \b[5]  & ~new_n11388_;
  assign new_n11445_ = ~new_n11386_ & new_n11444_;
  assign new_n11446_ = ~new_n11390_ & ~new_n11445_;
  assign new_n11447_ = ~new_n11443_ & new_n11446_;
  assign new_n11448_ = ~new_n11390_ & ~new_n11447_;
  assign new_n11449_ = \b[6]  & ~new_n11379_;
  assign new_n11450_ = ~new_n11377_ & new_n11449_;
  assign new_n11451_ = ~new_n11381_ & ~new_n11450_;
  assign new_n11452_ = ~new_n11448_ & new_n11451_;
  assign new_n11453_ = ~new_n11381_ & ~new_n11452_;
  assign new_n11454_ = \b[7]  & ~new_n11370_;
  assign new_n11455_ = ~new_n11368_ & new_n11454_;
  assign new_n11456_ = ~new_n11372_ & ~new_n11455_;
  assign new_n11457_ = ~new_n11453_ & new_n11456_;
  assign new_n11458_ = ~new_n11372_ & ~new_n11457_;
  assign new_n11459_ = \b[8]  & ~new_n11361_;
  assign new_n11460_ = ~new_n11359_ & new_n11459_;
  assign new_n11461_ = ~new_n11363_ & ~new_n11460_;
  assign new_n11462_ = ~new_n11458_ & new_n11461_;
  assign new_n11463_ = ~new_n11363_ & ~new_n11462_;
  assign new_n11464_ = \b[9]  & ~new_n11352_;
  assign new_n11465_ = ~new_n11350_ & new_n11464_;
  assign new_n11466_ = ~new_n11354_ & ~new_n11465_;
  assign new_n11467_ = ~new_n11463_ & new_n11466_;
  assign new_n11468_ = ~new_n11354_ & ~new_n11467_;
  assign new_n11469_ = \b[10]  & ~new_n11343_;
  assign new_n11470_ = ~new_n11341_ & new_n11469_;
  assign new_n11471_ = ~new_n11345_ & ~new_n11470_;
  assign new_n11472_ = ~new_n11468_ & new_n11471_;
  assign new_n11473_ = ~new_n11345_ & ~new_n11472_;
  assign new_n11474_ = \b[11]  & ~new_n11334_;
  assign new_n11475_ = ~new_n11332_ & new_n11474_;
  assign new_n11476_ = ~new_n11336_ & ~new_n11475_;
  assign new_n11477_ = ~new_n11473_ & new_n11476_;
  assign new_n11478_ = ~new_n11336_ & ~new_n11477_;
  assign new_n11479_ = \b[12]  & ~new_n11325_;
  assign new_n11480_ = ~new_n11323_ & new_n11479_;
  assign new_n11481_ = ~new_n11327_ & ~new_n11480_;
  assign new_n11482_ = ~new_n11478_ & new_n11481_;
  assign new_n11483_ = ~new_n11327_ & ~new_n11482_;
  assign new_n11484_ = \b[13]  & ~new_n11316_;
  assign new_n11485_ = ~new_n11314_ & new_n11484_;
  assign new_n11486_ = ~new_n11318_ & ~new_n11485_;
  assign new_n11487_ = ~new_n11483_ & new_n11486_;
  assign new_n11488_ = ~new_n11318_ & ~new_n11487_;
  assign new_n11489_ = \b[14]  & ~new_n11307_;
  assign new_n11490_ = ~new_n11305_ & new_n11489_;
  assign new_n11491_ = ~new_n11309_ & ~new_n11490_;
  assign new_n11492_ = ~new_n11488_ & new_n11491_;
  assign new_n11493_ = ~new_n11309_ & ~new_n11492_;
  assign new_n11494_ = \b[15]  & ~new_n11298_;
  assign new_n11495_ = ~new_n11296_ & new_n11494_;
  assign new_n11496_ = ~new_n11300_ & ~new_n11495_;
  assign new_n11497_ = ~new_n11493_ & new_n11496_;
  assign new_n11498_ = ~new_n11300_ & ~new_n11497_;
  assign new_n11499_ = \b[16]  & ~new_n11289_;
  assign new_n11500_ = ~new_n11287_ & new_n11499_;
  assign new_n11501_ = ~new_n11291_ & ~new_n11500_;
  assign new_n11502_ = ~new_n11498_ & new_n11501_;
  assign new_n11503_ = ~new_n11291_ & ~new_n11502_;
  assign new_n11504_ = \b[17]  & ~new_n11280_;
  assign new_n11505_ = ~new_n11278_ & new_n11504_;
  assign new_n11506_ = ~new_n11282_ & ~new_n11505_;
  assign new_n11507_ = ~new_n11503_ & new_n11506_;
  assign new_n11508_ = ~new_n11282_ & ~new_n11507_;
  assign new_n11509_ = \b[18]  & ~new_n11271_;
  assign new_n11510_ = ~new_n11269_ & new_n11509_;
  assign new_n11511_ = ~new_n11273_ & ~new_n11510_;
  assign new_n11512_ = ~new_n11508_ & new_n11511_;
  assign new_n11513_ = ~new_n11273_ & ~new_n11512_;
  assign new_n11514_ = \b[19]  & ~new_n11262_;
  assign new_n11515_ = ~new_n11260_ & new_n11514_;
  assign new_n11516_ = ~new_n11264_ & ~new_n11515_;
  assign new_n11517_ = ~new_n11513_ & new_n11516_;
  assign new_n11518_ = ~new_n11264_ & ~new_n11517_;
  assign new_n11519_ = \b[20]  & ~new_n11253_;
  assign new_n11520_ = ~new_n11251_ & new_n11519_;
  assign new_n11521_ = ~new_n11255_ & ~new_n11520_;
  assign new_n11522_ = ~new_n11518_ & new_n11521_;
  assign new_n11523_ = ~new_n11255_ & ~new_n11522_;
  assign new_n11524_ = \b[21]  & ~new_n11244_;
  assign new_n11525_ = ~new_n11242_ & new_n11524_;
  assign new_n11526_ = ~new_n11246_ & ~new_n11525_;
  assign new_n11527_ = ~new_n11523_ & new_n11526_;
  assign new_n11528_ = ~new_n11246_ & ~new_n11527_;
  assign new_n11529_ = \b[22]  & ~new_n11235_;
  assign new_n11530_ = ~new_n11233_ & new_n11529_;
  assign new_n11531_ = ~new_n11237_ & ~new_n11530_;
  assign new_n11532_ = ~new_n11528_ & new_n11531_;
  assign new_n11533_ = ~new_n11237_ & ~new_n11532_;
  assign new_n11534_ = \b[23]  & ~new_n11226_;
  assign new_n11535_ = ~new_n11224_ & new_n11534_;
  assign new_n11536_ = ~new_n11228_ & ~new_n11535_;
  assign new_n11537_ = ~new_n11533_ & new_n11536_;
  assign new_n11538_ = ~new_n11228_ & ~new_n11537_;
  assign new_n11539_ = \b[24]  & ~new_n11217_;
  assign new_n11540_ = ~new_n11215_ & new_n11539_;
  assign new_n11541_ = ~new_n11219_ & ~new_n11540_;
  assign new_n11542_ = ~new_n11538_ & new_n11541_;
  assign new_n11543_ = ~new_n11219_ & ~new_n11542_;
  assign new_n11544_ = \b[25]  & ~new_n11208_;
  assign new_n11545_ = ~new_n11206_ & new_n11544_;
  assign new_n11546_ = ~new_n11210_ & ~new_n11545_;
  assign new_n11547_ = ~new_n11543_ & new_n11546_;
  assign new_n11548_ = ~new_n11210_ & ~new_n11547_;
  assign new_n11549_ = \b[26]  & ~new_n11199_;
  assign new_n11550_ = ~new_n11197_ & new_n11549_;
  assign new_n11551_ = ~new_n11201_ & ~new_n11550_;
  assign new_n11552_ = ~new_n11548_ & new_n11551_;
  assign new_n11553_ = ~new_n11201_ & ~new_n11552_;
  assign new_n11554_ = \b[27]  & ~new_n11190_;
  assign new_n11555_ = ~new_n11188_ & new_n11554_;
  assign new_n11556_ = ~new_n11192_ & ~new_n11555_;
  assign new_n11557_ = ~new_n11553_ & new_n11556_;
  assign new_n11558_ = ~new_n11192_ & ~new_n11557_;
  assign new_n11559_ = \b[28]  & ~new_n11181_;
  assign new_n11560_ = ~new_n11179_ & new_n11559_;
  assign new_n11561_ = ~new_n11183_ & ~new_n11560_;
  assign new_n11562_ = ~new_n11558_ & new_n11561_;
  assign new_n11563_ = ~new_n11183_ & ~new_n11562_;
  assign new_n11564_ = \b[29]  & ~new_n11172_;
  assign new_n11565_ = ~new_n11170_ & new_n11564_;
  assign new_n11566_ = ~new_n11174_ & ~new_n11565_;
  assign new_n11567_ = ~new_n11563_ & new_n11566_;
  assign new_n11568_ = ~new_n11174_ & ~new_n11567_;
  assign new_n11569_ = \b[30]  & ~new_n11163_;
  assign new_n11570_ = ~new_n11161_ & new_n11569_;
  assign new_n11571_ = ~new_n11165_ & ~new_n11570_;
  assign new_n11572_ = ~new_n11568_ & new_n11571_;
  assign new_n11573_ = ~new_n11165_ & ~new_n11572_;
  assign new_n11574_ = \b[31]  & ~new_n11154_;
  assign new_n11575_ = ~new_n11152_ & new_n11574_;
  assign new_n11576_ = ~new_n11156_ & ~new_n11575_;
  assign new_n11577_ = ~new_n11573_ & new_n11576_;
  assign new_n11578_ = ~new_n11156_ & ~new_n11577_;
  assign new_n11579_ = \b[32]  & ~new_n11145_;
  assign new_n11580_ = ~new_n11143_ & new_n11579_;
  assign new_n11581_ = ~new_n11147_ & ~new_n11580_;
  assign new_n11582_ = ~new_n11578_ & new_n11581_;
  assign new_n11583_ = ~new_n11147_ & ~new_n11582_;
  assign new_n11584_ = \b[33]  & ~new_n11136_;
  assign new_n11585_ = ~new_n11134_ & new_n11584_;
  assign new_n11586_ = ~new_n11138_ & ~new_n11585_;
  assign new_n11587_ = ~new_n11583_ & new_n11586_;
  assign new_n11588_ = ~new_n11138_ & ~new_n11587_;
  assign new_n11589_ = \b[34]  & ~new_n11127_;
  assign new_n11590_ = ~new_n11125_ & new_n11589_;
  assign new_n11591_ = ~new_n11129_ & ~new_n11590_;
  assign new_n11592_ = ~new_n11588_ & new_n11591_;
  assign new_n11593_ = ~new_n11129_ & ~new_n11592_;
  assign new_n11594_ = \b[35]  & ~new_n11118_;
  assign new_n11595_ = ~new_n11116_ & new_n11594_;
  assign new_n11596_ = ~new_n11120_ & ~new_n11595_;
  assign new_n11597_ = ~new_n11593_ & new_n11596_;
  assign new_n11598_ = ~new_n11120_ & ~new_n11597_;
  assign new_n11599_ = \b[36]  & ~new_n11109_;
  assign new_n11600_ = ~new_n11107_ & new_n11599_;
  assign new_n11601_ = ~new_n11111_ & ~new_n11600_;
  assign new_n11602_ = ~new_n11598_ & new_n11601_;
  assign new_n11603_ = ~new_n11111_ & ~new_n11602_;
  assign new_n11604_ = \b[37]  & ~new_n11100_;
  assign new_n11605_ = ~new_n11098_ & new_n11604_;
  assign new_n11606_ = ~new_n11102_ & ~new_n11605_;
  assign new_n11607_ = ~new_n11603_ & new_n11606_;
  assign new_n11608_ = ~new_n11102_ & ~new_n11607_;
  assign new_n11609_ = \b[38]  & ~new_n11080_;
  assign new_n11610_ = ~new_n11078_ & new_n11609_;
  assign new_n11611_ = ~new_n11093_ & ~new_n11610_;
  assign new_n11612_ = ~new_n11608_ & new_n11611_;
  assign new_n11613_ = ~new_n11093_ & ~new_n11612_;
  assign new_n11614_ = \b[39]  & ~new_n11090_;
  assign new_n11615_ = ~new_n11088_ & new_n11614_;
  assign new_n11616_ = ~new_n11092_ & ~new_n11615_;
  assign new_n11617_ = ~new_n11613_ & new_n11616_;
  assign new_n11618_ = ~new_n11092_ & ~new_n11617_;
  assign new_n11619_ = new_n338_ & new_n340_;
  assign \quotient[24]  = ~new_n11618_ & new_n11619_;
  assign new_n11621_ = ~new_n11081_ & ~\quotient[24] ;
  assign new_n11622_ = ~new_n11102_ & new_n11611_;
  assign new_n11623_ = ~new_n11607_ & new_n11622_;
  assign new_n11624_ = ~new_n11608_ & ~new_n11611_;
  assign new_n11625_ = ~new_n11623_ & ~new_n11624_;
  assign new_n11626_ = new_n11619_ & ~new_n11625_;
  assign new_n11627_ = ~new_n11618_ & new_n11626_;
  assign new_n11628_ = ~new_n11621_ & ~new_n11627_;
  assign new_n11629_ = ~new_n11091_ & ~\quotient[24] ;
  assign new_n11630_ = ~new_n11093_ & new_n11616_;
  assign new_n11631_ = ~new_n11612_ & new_n11630_;
  assign new_n11632_ = ~new_n11613_ & ~new_n11616_;
  assign new_n11633_ = ~new_n11631_ & ~new_n11632_;
  assign new_n11634_ = \quotient[24]  & ~new_n11633_;
  assign new_n11635_ = ~new_n11629_ & ~new_n11634_;
  assign new_n11636_ = ~\b[40]  & ~new_n11635_;
  assign new_n11637_ = ~\b[39]  & ~new_n11628_;
  assign new_n11638_ = ~new_n11101_ & ~\quotient[24] ;
  assign new_n11639_ = ~new_n11111_ & new_n11606_;
  assign new_n11640_ = ~new_n11602_ & new_n11639_;
  assign new_n11641_ = ~new_n11603_ & ~new_n11606_;
  assign new_n11642_ = ~new_n11640_ & ~new_n11641_;
  assign new_n11643_ = new_n11619_ & ~new_n11642_;
  assign new_n11644_ = ~new_n11618_ & new_n11643_;
  assign new_n11645_ = ~new_n11638_ & ~new_n11644_;
  assign new_n11646_ = ~\b[38]  & ~new_n11645_;
  assign new_n11647_ = ~new_n11110_ & ~\quotient[24] ;
  assign new_n11648_ = ~new_n11120_ & new_n11601_;
  assign new_n11649_ = ~new_n11597_ & new_n11648_;
  assign new_n11650_ = ~new_n11598_ & ~new_n11601_;
  assign new_n11651_ = ~new_n11649_ & ~new_n11650_;
  assign new_n11652_ = new_n11619_ & ~new_n11651_;
  assign new_n11653_ = ~new_n11618_ & new_n11652_;
  assign new_n11654_ = ~new_n11647_ & ~new_n11653_;
  assign new_n11655_ = ~\b[37]  & ~new_n11654_;
  assign new_n11656_ = ~new_n11119_ & ~\quotient[24] ;
  assign new_n11657_ = ~new_n11129_ & new_n11596_;
  assign new_n11658_ = ~new_n11592_ & new_n11657_;
  assign new_n11659_ = ~new_n11593_ & ~new_n11596_;
  assign new_n11660_ = ~new_n11658_ & ~new_n11659_;
  assign new_n11661_ = new_n11619_ & ~new_n11660_;
  assign new_n11662_ = ~new_n11618_ & new_n11661_;
  assign new_n11663_ = ~new_n11656_ & ~new_n11662_;
  assign new_n11664_ = ~\b[36]  & ~new_n11663_;
  assign new_n11665_ = ~new_n11128_ & ~\quotient[24] ;
  assign new_n11666_ = ~new_n11138_ & new_n11591_;
  assign new_n11667_ = ~new_n11587_ & new_n11666_;
  assign new_n11668_ = ~new_n11588_ & ~new_n11591_;
  assign new_n11669_ = ~new_n11667_ & ~new_n11668_;
  assign new_n11670_ = new_n11619_ & ~new_n11669_;
  assign new_n11671_ = ~new_n11618_ & new_n11670_;
  assign new_n11672_ = ~new_n11665_ & ~new_n11671_;
  assign new_n11673_ = ~\b[35]  & ~new_n11672_;
  assign new_n11674_ = ~new_n11137_ & ~\quotient[24] ;
  assign new_n11675_ = ~new_n11147_ & new_n11586_;
  assign new_n11676_ = ~new_n11582_ & new_n11675_;
  assign new_n11677_ = ~new_n11583_ & ~new_n11586_;
  assign new_n11678_ = ~new_n11676_ & ~new_n11677_;
  assign new_n11679_ = new_n11619_ & ~new_n11678_;
  assign new_n11680_ = ~new_n11618_ & new_n11679_;
  assign new_n11681_ = ~new_n11674_ & ~new_n11680_;
  assign new_n11682_ = ~\b[34]  & ~new_n11681_;
  assign new_n11683_ = ~new_n11146_ & ~\quotient[24] ;
  assign new_n11684_ = ~new_n11156_ & new_n11581_;
  assign new_n11685_ = ~new_n11577_ & new_n11684_;
  assign new_n11686_ = ~new_n11578_ & ~new_n11581_;
  assign new_n11687_ = ~new_n11685_ & ~new_n11686_;
  assign new_n11688_ = new_n11619_ & ~new_n11687_;
  assign new_n11689_ = ~new_n11618_ & new_n11688_;
  assign new_n11690_ = ~new_n11683_ & ~new_n11689_;
  assign new_n11691_ = ~\b[33]  & ~new_n11690_;
  assign new_n11692_ = ~new_n11155_ & ~\quotient[24] ;
  assign new_n11693_ = ~new_n11165_ & new_n11576_;
  assign new_n11694_ = ~new_n11572_ & new_n11693_;
  assign new_n11695_ = ~new_n11573_ & ~new_n11576_;
  assign new_n11696_ = ~new_n11694_ & ~new_n11695_;
  assign new_n11697_ = new_n11619_ & ~new_n11696_;
  assign new_n11698_ = ~new_n11618_ & new_n11697_;
  assign new_n11699_ = ~new_n11692_ & ~new_n11698_;
  assign new_n11700_ = ~\b[32]  & ~new_n11699_;
  assign new_n11701_ = ~new_n11164_ & ~\quotient[24] ;
  assign new_n11702_ = ~new_n11174_ & new_n11571_;
  assign new_n11703_ = ~new_n11567_ & new_n11702_;
  assign new_n11704_ = ~new_n11568_ & ~new_n11571_;
  assign new_n11705_ = ~new_n11703_ & ~new_n11704_;
  assign new_n11706_ = new_n11619_ & ~new_n11705_;
  assign new_n11707_ = ~new_n11618_ & new_n11706_;
  assign new_n11708_ = ~new_n11701_ & ~new_n11707_;
  assign new_n11709_ = ~\b[31]  & ~new_n11708_;
  assign new_n11710_ = ~new_n11173_ & ~\quotient[24] ;
  assign new_n11711_ = ~new_n11183_ & new_n11566_;
  assign new_n11712_ = ~new_n11562_ & new_n11711_;
  assign new_n11713_ = ~new_n11563_ & ~new_n11566_;
  assign new_n11714_ = ~new_n11712_ & ~new_n11713_;
  assign new_n11715_ = new_n11619_ & ~new_n11714_;
  assign new_n11716_ = ~new_n11618_ & new_n11715_;
  assign new_n11717_ = ~new_n11710_ & ~new_n11716_;
  assign new_n11718_ = ~\b[30]  & ~new_n11717_;
  assign new_n11719_ = ~new_n11182_ & ~\quotient[24] ;
  assign new_n11720_ = ~new_n11192_ & new_n11561_;
  assign new_n11721_ = ~new_n11557_ & new_n11720_;
  assign new_n11722_ = ~new_n11558_ & ~new_n11561_;
  assign new_n11723_ = ~new_n11721_ & ~new_n11722_;
  assign new_n11724_ = new_n11619_ & ~new_n11723_;
  assign new_n11725_ = ~new_n11618_ & new_n11724_;
  assign new_n11726_ = ~new_n11719_ & ~new_n11725_;
  assign new_n11727_ = ~\b[29]  & ~new_n11726_;
  assign new_n11728_ = ~new_n11191_ & ~\quotient[24] ;
  assign new_n11729_ = ~new_n11201_ & new_n11556_;
  assign new_n11730_ = ~new_n11552_ & new_n11729_;
  assign new_n11731_ = ~new_n11553_ & ~new_n11556_;
  assign new_n11732_ = ~new_n11730_ & ~new_n11731_;
  assign new_n11733_ = new_n11619_ & ~new_n11732_;
  assign new_n11734_ = ~new_n11618_ & new_n11733_;
  assign new_n11735_ = ~new_n11728_ & ~new_n11734_;
  assign new_n11736_ = ~\b[28]  & ~new_n11735_;
  assign new_n11737_ = ~new_n11200_ & ~\quotient[24] ;
  assign new_n11738_ = ~new_n11210_ & new_n11551_;
  assign new_n11739_ = ~new_n11547_ & new_n11738_;
  assign new_n11740_ = ~new_n11548_ & ~new_n11551_;
  assign new_n11741_ = ~new_n11739_ & ~new_n11740_;
  assign new_n11742_ = new_n11619_ & ~new_n11741_;
  assign new_n11743_ = ~new_n11618_ & new_n11742_;
  assign new_n11744_ = ~new_n11737_ & ~new_n11743_;
  assign new_n11745_ = ~\b[27]  & ~new_n11744_;
  assign new_n11746_ = ~new_n11209_ & ~\quotient[24] ;
  assign new_n11747_ = ~new_n11219_ & new_n11546_;
  assign new_n11748_ = ~new_n11542_ & new_n11747_;
  assign new_n11749_ = ~new_n11543_ & ~new_n11546_;
  assign new_n11750_ = ~new_n11748_ & ~new_n11749_;
  assign new_n11751_ = new_n11619_ & ~new_n11750_;
  assign new_n11752_ = ~new_n11618_ & new_n11751_;
  assign new_n11753_ = ~new_n11746_ & ~new_n11752_;
  assign new_n11754_ = ~\b[26]  & ~new_n11753_;
  assign new_n11755_ = ~new_n11218_ & ~\quotient[24] ;
  assign new_n11756_ = ~new_n11228_ & new_n11541_;
  assign new_n11757_ = ~new_n11537_ & new_n11756_;
  assign new_n11758_ = ~new_n11538_ & ~new_n11541_;
  assign new_n11759_ = ~new_n11757_ & ~new_n11758_;
  assign new_n11760_ = new_n11619_ & ~new_n11759_;
  assign new_n11761_ = ~new_n11618_ & new_n11760_;
  assign new_n11762_ = ~new_n11755_ & ~new_n11761_;
  assign new_n11763_ = ~\b[25]  & ~new_n11762_;
  assign new_n11764_ = ~new_n11227_ & ~\quotient[24] ;
  assign new_n11765_ = ~new_n11237_ & new_n11536_;
  assign new_n11766_ = ~new_n11532_ & new_n11765_;
  assign new_n11767_ = ~new_n11533_ & ~new_n11536_;
  assign new_n11768_ = ~new_n11766_ & ~new_n11767_;
  assign new_n11769_ = new_n11619_ & ~new_n11768_;
  assign new_n11770_ = ~new_n11618_ & new_n11769_;
  assign new_n11771_ = ~new_n11764_ & ~new_n11770_;
  assign new_n11772_ = ~\b[24]  & ~new_n11771_;
  assign new_n11773_ = ~new_n11236_ & ~\quotient[24] ;
  assign new_n11774_ = ~new_n11246_ & new_n11531_;
  assign new_n11775_ = ~new_n11527_ & new_n11774_;
  assign new_n11776_ = ~new_n11528_ & ~new_n11531_;
  assign new_n11777_ = ~new_n11775_ & ~new_n11776_;
  assign new_n11778_ = new_n11619_ & ~new_n11777_;
  assign new_n11779_ = ~new_n11618_ & new_n11778_;
  assign new_n11780_ = ~new_n11773_ & ~new_n11779_;
  assign new_n11781_ = ~\b[23]  & ~new_n11780_;
  assign new_n11782_ = ~new_n11245_ & ~\quotient[24] ;
  assign new_n11783_ = ~new_n11255_ & new_n11526_;
  assign new_n11784_ = ~new_n11522_ & new_n11783_;
  assign new_n11785_ = ~new_n11523_ & ~new_n11526_;
  assign new_n11786_ = ~new_n11784_ & ~new_n11785_;
  assign new_n11787_ = new_n11619_ & ~new_n11786_;
  assign new_n11788_ = ~new_n11618_ & new_n11787_;
  assign new_n11789_ = ~new_n11782_ & ~new_n11788_;
  assign new_n11790_ = ~\b[22]  & ~new_n11789_;
  assign new_n11791_ = ~new_n11254_ & ~\quotient[24] ;
  assign new_n11792_ = ~new_n11264_ & new_n11521_;
  assign new_n11793_ = ~new_n11517_ & new_n11792_;
  assign new_n11794_ = ~new_n11518_ & ~new_n11521_;
  assign new_n11795_ = ~new_n11793_ & ~new_n11794_;
  assign new_n11796_ = new_n11619_ & ~new_n11795_;
  assign new_n11797_ = ~new_n11618_ & new_n11796_;
  assign new_n11798_ = ~new_n11791_ & ~new_n11797_;
  assign new_n11799_ = ~\b[21]  & ~new_n11798_;
  assign new_n11800_ = ~new_n11263_ & ~\quotient[24] ;
  assign new_n11801_ = ~new_n11273_ & new_n11516_;
  assign new_n11802_ = ~new_n11512_ & new_n11801_;
  assign new_n11803_ = ~new_n11513_ & ~new_n11516_;
  assign new_n11804_ = ~new_n11802_ & ~new_n11803_;
  assign new_n11805_ = new_n11619_ & ~new_n11804_;
  assign new_n11806_ = ~new_n11618_ & new_n11805_;
  assign new_n11807_ = ~new_n11800_ & ~new_n11806_;
  assign new_n11808_ = ~\b[20]  & ~new_n11807_;
  assign new_n11809_ = ~new_n11272_ & ~\quotient[24] ;
  assign new_n11810_ = ~new_n11282_ & new_n11511_;
  assign new_n11811_ = ~new_n11507_ & new_n11810_;
  assign new_n11812_ = ~new_n11508_ & ~new_n11511_;
  assign new_n11813_ = ~new_n11811_ & ~new_n11812_;
  assign new_n11814_ = new_n11619_ & ~new_n11813_;
  assign new_n11815_ = ~new_n11618_ & new_n11814_;
  assign new_n11816_ = ~new_n11809_ & ~new_n11815_;
  assign new_n11817_ = ~\b[19]  & ~new_n11816_;
  assign new_n11818_ = ~new_n11281_ & ~\quotient[24] ;
  assign new_n11819_ = ~new_n11291_ & new_n11506_;
  assign new_n11820_ = ~new_n11502_ & new_n11819_;
  assign new_n11821_ = ~new_n11503_ & ~new_n11506_;
  assign new_n11822_ = ~new_n11820_ & ~new_n11821_;
  assign new_n11823_ = new_n11619_ & ~new_n11822_;
  assign new_n11824_ = ~new_n11618_ & new_n11823_;
  assign new_n11825_ = ~new_n11818_ & ~new_n11824_;
  assign new_n11826_ = ~\b[18]  & ~new_n11825_;
  assign new_n11827_ = ~new_n11290_ & ~\quotient[24] ;
  assign new_n11828_ = ~new_n11300_ & new_n11501_;
  assign new_n11829_ = ~new_n11497_ & new_n11828_;
  assign new_n11830_ = ~new_n11498_ & ~new_n11501_;
  assign new_n11831_ = ~new_n11829_ & ~new_n11830_;
  assign new_n11832_ = new_n11619_ & ~new_n11831_;
  assign new_n11833_ = ~new_n11618_ & new_n11832_;
  assign new_n11834_ = ~new_n11827_ & ~new_n11833_;
  assign new_n11835_ = ~\b[17]  & ~new_n11834_;
  assign new_n11836_ = ~new_n11299_ & ~\quotient[24] ;
  assign new_n11837_ = ~new_n11309_ & new_n11496_;
  assign new_n11838_ = ~new_n11492_ & new_n11837_;
  assign new_n11839_ = ~new_n11493_ & ~new_n11496_;
  assign new_n11840_ = ~new_n11838_ & ~new_n11839_;
  assign new_n11841_ = new_n11619_ & ~new_n11840_;
  assign new_n11842_ = ~new_n11618_ & new_n11841_;
  assign new_n11843_ = ~new_n11836_ & ~new_n11842_;
  assign new_n11844_ = ~\b[16]  & ~new_n11843_;
  assign new_n11845_ = ~new_n11308_ & ~\quotient[24] ;
  assign new_n11846_ = ~new_n11318_ & new_n11491_;
  assign new_n11847_ = ~new_n11487_ & new_n11846_;
  assign new_n11848_ = ~new_n11488_ & ~new_n11491_;
  assign new_n11849_ = ~new_n11847_ & ~new_n11848_;
  assign new_n11850_ = new_n11619_ & ~new_n11849_;
  assign new_n11851_ = ~new_n11618_ & new_n11850_;
  assign new_n11852_ = ~new_n11845_ & ~new_n11851_;
  assign new_n11853_ = ~\b[15]  & ~new_n11852_;
  assign new_n11854_ = ~new_n11317_ & ~\quotient[24] ;
  assign new_n11855_ = ~new_n11327_ & new_n11486_;
  assign new_n11856_ = ~new_n11482_ & new_n11855_;
  assign new_n11857_ = ~new_n11483_ & ~new_n11486_;
  assign new_n11858_ = ~new_n11856_ & ~new_n11857_;
  assign new_n11859_ = new_n11619_ & ~new_n11858_;
  assign new_n11860_ = ~new_n11618_ & new_n11859_;
  assign new_n11861_ = ~new_n11854_ & ~new_n11860_;
  assign new_n11862_ = ~\b[14]  & ~new_n11861_;
  assign new_n11863_ = ~new_n11326_ & ~\quotient[24] ;
  assign new_n11864_ = ~new_n11336_ & new_n11481_;
  assign new_n11865_ = ~new_n11477_ & new_n11864_;
  assign new_n11866_ = ~new_n11478_ & ~new_n11481_;
  assign new_n11867_ = ~new_n11865_ & ~new_n11866_;
  assign new_n11868_ = new_n11619_ & ~new_n11867_;
  assign new_n11869_ = ~new_n11618_ & new_n11868_;
  assign new_n11870_ = ~new_n11863_ & ~new_n11869_;
  assign new_n11871_ = ~\b[13]  & ~new_n11870_;
  assign new_n11872_ = ~new_n11335_ & ~\quotient[24] ;
  assign new_n11873_ = ~new_n11345_ & new_n11476_;
  assign new_n11874_ = ~new_n11472_ & new_n11873_;
  assign new_n11875_ = ~new_n11473_ & ~new_n11476_;
  assign new_n11876_ = ~new_n11874_ & ~new_n11875_;
  assign new_n11877_ = new_n11619_ & ~new_n11876_;
  assign new_n11878_ = ~new_n11618_ & new_n11877_;
  assign new_n11879_ = ~new_n11872_ & ~new_n11878_;
  assign new_n11880_ = ~\b[12]  & ~new_n11879_;
  assign new_n11881_ = ~new_n11344_ & ~\quotient[24] ;
  assign new_n11882_ = ~new_n11354_ & new_n11471_;
  assign new_n11883_ = ~new_n11467_ & new_n11882_;
  assign new_n11884_ = ~new_n11468_ & ~new_n11471_;
  assign new_n11885_ = ~new_n11883_ & ~new_n11884_;
  assign new_n11886_ = new_n11619_ & ~new_n11885_;
  assign new_n11887_ = ~new_n11618_ & new_n11886_;
  assign new_n11888_ = ~new_n11881_ & ~new_n11887_;
  assign new_n11889_ = ~\b[11]  & ~new_n11888_;
  assign new_n11890_ = ~new_n11353_ & ~\quotient[24] ;
  assign new_n11891_ = ~new_n11363_ & new_n11466_;
  assign new_n11892_ = ~new_n11462_ & new_n11891_;
  assign new_n11893_ = ~new_n11463_ & ~new_n11466_;
  assign new_n11894_ = ~new_n11892_ & ~new_n11893_;
  assign new_n11895_ = new_n11619_ & ~new_n11894_;
  assign new_n11896_ = ~new_n11618_ & new_n11895_;
  assign new_n11897_ = ~new_n11890_ & ~new_n11896_;
  assign new_n11898_ = ~\b[10]  & ~new_n11897_;
  assign new_n11899_ = ~new_n11362_ & ~\quotient[24] ;
  assign new_n11900_ = ~new_n11372_ & new_n11461_;
  assign new_n11901_ = ~new_n11457_ & new_n11900_;
  assign new_n11902_ = ~new_n11458_ & ~new_n11461_;
  assign new_n11903_ = ~new_n11901_ & ~new_n11902_;
  assign new_n11904_ = new_n11619_ & ~new_n11903_;
  assign new_n11905_ = ~new_n11618_ & new_n11904_;
  assign new_n11906_ = ~new_n11899_ & ~new_n11905_;
  assign new_n11907_ = ~\b[9]  & ~new_n11906_;
  assign new_n11908_ = ~new_n11371_ & ~\quotient[24] ;
  assign new_n11909_ = ~new_n11381_ & new_n11456_;
  assign new_n11910_ = ~new_n11452_ & new_n11909_;
  assign new_n11911_ = ~new_n11453_ & ~new_n11456_;
  assign new_n11912_ = ~new_n11910_ & ~new_n11911_;
  assign new_n11913_ = new_n11619_ & ~new_n11912_;
  assign new_n11914_ = ~new_n11618_ & new_n11913_;
  assign new_n11915_ = ~new_n11908_ & ~new_n11914_;
  assign new_n11916_ = ~\b[8]  & ~new_n11915_;
  assign new_n11917_ = ~new_n11380_ & ~\quotient[24] ;
  assign new_n11918_ = ~new_n11390_ & new_n11451_;
  assign new_n11919_ = ~new_n11447_ & new_n11918_;
  assign new_n11920_ = ~new_n11448_ & ~new_n11451_;
  assign new_n11921_ = ~new_n11919_ & ~new_n11920_;
  assign new_n11922_ = new_n11619_ & ~new_n11921_;
  assign new_n11923_ = ~new_n11618_ & new_n11922_;
  assign new_n11924_ = ~new_n11917_ & ~new_n11923_;
  assign new_n11925_ = ~\b[7]  & ~new_n11924_;
  assign new_n11926_ = ~new_n11389_ & ~\quotient[24] ;
  assign new_n11927_ = ~new_n11399_ & new_n11446_;
  assign new_n11928_ = ~new_n11442_ & new_n11927_;
  assign new_n11929_ = ~new_n11443_ & ~new_n11446_;
  assign new_n11930_ = ~new_n11928_ & ~new_n11929_;
  assign new_n11931_ = new_n11619_ & ~new_n11930_;
  assign new_n11932_ = ~new_n11618_ & new_n11931_;
  assign new_n11933_ = ~new_n11926_ & ~new_n11932_;
  assign new_n11934_ = ~\b[6]  & ~new_n11933_;
  assign new_n11935_ = ~new_n11398_ & ~\quotient[24] ;
  assign new_n11936_ = ~new_n11408_ & new_n11441_;
  assign new_n11937_ = ~new_n11437_ & new_n11936_;
  assign new_n11938_ = ~new_n11438_ & ~new_n11441_;
  assign new_n11939_ = ~new_n11937_ & ~new_n11938_;
  assign new_n11940_ = new_n11619_ & ~new_n11939_;
  assign new_n11941_ = ~new_n11618_ & new_n11940_;
  assign new_n11942_ = ~new_n11935_ & ~new_n11941_;
  assign new_n11943_ = ~\b[5]  & ~new_n11942_;
  assign new_n11944_ = ~new_n11407_ & ~\quotient[24] ;
  assign new_n11945_ = ~new_n11416_ & new_n11436_;
  assign new_n11946_ = ~new_n11432_ & new_n11945_;
  assign new_n11947_ = ~new_n11433_ & ~new_n11436_;
  assign new_n11948_ = ~new_n11946_ & ~new_n11947_;
  assign new_n11949_ = new_n11619_ & ~new_n11948_;
  assign new_n11950_ = ~new_n11618_ & new_n11949_;
  assign new_n11951_ = ~new_n11944_ & ~new_n11950_;
  assign new_n11952_ = ~\b[4]  & ~new_n11951_;
  assign new_n11953_ = ~new_n11415_ & ~\quotient[24] ;
  assign new_n11954_ = ~new_n11427_ & new_n11431_;
  assign new_n11955_ = ~new_n11426_ & new_n11954_;
  assign new_n11956_ = ~new_n11428_ & ~new_n11431_;
  assign new_n11957_ = ~new_n11955_ & ~new_n11956_;
  assign new_n11958_ = new_n11619_ & ~new_n11957_;
  assign new_n11959_ = ~new_n11618_ & new_n11958_;
  assign new_n11960_ = ~new_n11953_ & ~new_n11959_;
  assign new_n11961_ = ~\b[3]  & ~new_n11960_;
  assign new_n11962_ = ~new_n11420_ & ~\quotient[24] ;
  assign new_n11963_ = ~new_n11423_ & new_n11425_;
  assign new_n11964_ = ~new_n11421_ & new_n11963_;
  assign new_n11965_ = new_n11619_ & ~new_n11964_;
  assign new_n11966_ = ~new_n11426_ & new_n11965_;
  assign new_n11967_ = ~new_n11618_ & new_n11966_;
  assign new_n11968_ = ~new_n11962_ & ~new_n11967_;
  assign new_n11969_ = ~\b[2]  & ~new_n11968_;
  assign new_n11970_ = \b[0]  & ~\b[40] ;
  assign new_n11971_ = new_n421_ & new_n11970_;
  assign new_n11972_ = new_n597_ & new_n11971_;
  assign new_n11973_ = new_n595_ & new_n11972_;
  assign new_n11974_ = ~new_n11618_ & new_n11973_;
  assign new_n11975_ = \a[24]  & ~new_n11974_;
  assign new_n11976_ = new_n291_ & new_n11425_;
  assign new_n11977_ = new_n302_ & new_n11976_;
  assign new_n11978_ = new_n288_ & new_n11977_;
  assign new_n11979_ = ~new_n11618_ & new_n11978_;
  assign new_n11980_ = ~new_n11975_ & ~new_n11979_;
  assign new_n11981_ = \b[1]  & ~new_n11980_;
  assign new_n11982_ = ~\b[1]  & ~new_n11979_;
  assign new_n11983_ = ~new_n11975_ & new_n11982_;
  assign new_n11984_ = ~new_n11981_ & ~new_n11983_;
  assign new_n11985_ = ~\a[23]  & \b[0] ;
  assign new_n11986_ = ~new_n11984_ & ~new_n11985_;
  assign new_n11987_ = ~\b[1]  & ~new_n11980_;
  assign new_n11988_ = ~new_n11986_ & ~new_n11987_;
  assign new_n11989_ = \b[2]  & ~new_n11967_;
  assign new_n11990_ = ~new_n11962_ & new_n11989_;
  assign new_n11991_ = ~new_n11969_ & ~new_n11990_;
  assign new_n11992_ = ~new_n11988_ & new_n11991_;
  assign new_n11993_ = ~new_n11969_ & ~new_n11992_;
  assign new_n11994_ = \b[3]  & ~new_n11959_;
  assign new_n11995_ = ~new_n11953_ & new_n11994_;
  assign new_n11996_ = ~new_n11961_ & ~new_n11995_;
  assign new_n11997_ = ~new_n11993_ & new_n11996_;
  assign new_n11998_ = ~new_n11961_ & ~new_n11997_;
  assign new_n11999_ = \b[4]  & ~new_n11950_;
  assign new_n12000_ = ~new_n11944_ & new_n11999_;
  assign new_n12001_ = ~new_n11952_ & ~new_n12000_;
  assign new_n12002_ = ~new_n11998_ & new_n12001_;
  assign new_n12003_ = ~new_n11952_ & ~new_n12002_;
  assign new_n12004_ = \b[5]  & ~new_n11941_;
  assign new_n12005_ = ~new_n11935_ & new_n12004_;
  assign new_n12006_ = ~new_n11943_ & ~new_n12005_;
  assign new_n12007_ = ~new_n12003_ & new_n12006_;
  assign new_n12008_ = ~new_n11943_ & ~new_n12007_;
  assign new_n12009_ = \b[6]  & ~new_n11932_;
  assign new_n12010_ = ~new_n11926_ & new_n12009_;
  assign new_n12011_ = ~new_n11934_ & ~new_n12010_;
  assign new_n12012_ = ~new_n12008_ & new_n12011_;
  assign new_n12013_ = ~new_n11934_ & ~new_n12012_;
  assign new_n12014_ = \b[7]  & ~new_n11923_;
  assign new_n12015_ = ~new_n11917_ & new_n12014_;
  assign new_n12016_ = ~new_n11925_ & ~new_n12015_;
  assign new_n12017_ = ~new_n12013_ & new_n12016_;
  assign new_n12018_ = ~new_n11925_ & ~new_n12017_;
  assign new_n12019_ = \b[8]  & ~new_n11914_;
  assign new_n12020_ = ~new_n11908_ & new_n12019_;
  assign new_n12021_ = ~new_n11916_ & ~new_n12020_;
  assign new_n12022_ = ~new_n12018_ & new_n12021_;
  assign new_n12023_ = ~new_n11916_ & ~new_n12022_;
  assign new_n12024_ = \b[9]  & ~new_n11905_;
  assign new_n12025_ = ~new_n11899_ & new_n12024_;
  assign new_n12026_ = ~new_n11907_ & ~new_n12025_;
  assign new_n12027_ = ~new_n12023_ & new_n12026_;
  assign new_n12028_ = ~new_n11907_ & ~new_n12027_;
  assign new_n12029_ = \b[10]  & ~new_n11896_;
  assign new_n12030_ = ~new_n11890_ & new_n12029_;
  assign new_n12031_ = ~new_n11898_ & ~new_n12030_;
  assign new_n12032_ = ~new_n12028_ & new_n12031_;
  assign new_n12033_ = ~new_n11898_ & ~new_n12032_;
  assign new_n12034_ = \b[11]  & ~new_n11887_;
  assign new_n12035_ = ~new_n11881_ & new_n12034_;
  assign new_n12036_ = ~new_n11889_ & ~new_n12035_;
  assign new_n12037_ = ~new_n12033_ & new_n12036_;
  assign new_n12038_ = ~new_n11889_ & ~new_n12037_;
  assign new_n12039_ = \b[12]  & ~new_n11878_;
  assign new_n12040_ = ~new_n11872_ & new_n12039_;
  assign new_n12041_ = ~new_n11880_ & ~new_n12040_;
  assign new_n12042_ = ~new_n12038_ & new_n12041_;
  assign new_n12043_ = ~new_n11880_ & ~new_n12042_;
  assign new_n12044_ = \b[13]  & ~new_n11869_;
  assign new_n12045_ = ~new_n11863_ & new_n12044_;
  assign new_n12046_ = ~new_n11871_ & ~new_n12045_;
  assign new_n12047_ = ~new_n12043_ & new_n12046_;
  assign new_n12048_ = ~new_n11871_ & ~new_n12047_;
  assign new_n12049_ = \b[14]  & ~new_n11860_;
  assign new_n12050_ = ~new_n11854_ & new_n12049_;
  assign new_n12051_ = ~new_n11862_ & ~new_n12050_;
  assign new_n12052_ = ~new_n12048_ & new_n12051_;
  assign new_n12053_ = ~new_n11862_ & ~new_n12052_;
  assign new_n12054_ = \b[15]  & ~new_n11851_;
  assign new_n12055_ = ~new_n11845_ & new_n12054_;
  assign new_n12056_ = ~new_n11853_ & ~new_n12055_;
  assign new_n12057_ = ~new_n12053_ & new_n12056_;
  assign new_n12058_ = ~new_n11853_ & ~new_n12057_;
  assign new_n12059_ = \b[16]  & ~new_n11842_;
  assign new_n12060_ = ~new_n11836_ & new_n12059_;
  assign new_n12061_ = ~new_n11844_ & ~new_n12060_;
  assign new_n12062_ = ~new_n12058_ & new_n12061_;
  assign new_n12063_ = ~new_n11844_ & ~new_n12062_;
  assign new_n12064_ = \b[17]  & ~new_n11833_;
  assign new_n12065_ = ~new_n11827_ & new_n12064_;
  assign new_n12066_ = ~new_n11835_ & ~new_n12065_;
  assign new_n12067_ = ~new_n12063_ & new_n12066_;
  assign new_n12068_ = ~new_n11835_ & ~new_n12067_;
  assign new_n12069_ = \b[18]  & ~new_n11824_;
  assign new_n12070_ = ~new_n11818_ & new_n12069_;
  assign new_n12071_ = ~new_n11826_ & ~new_n12070_;
  assign new_n12072_ = ~new_n12068_ & new_n12071_;
  assign new_n12073_ = ~new_n11826_ & ~new_n12072_;
  assign new_n12074_ = \b[19]  & ~new_n11815_;
  assign new_n12075_ = ~new_n11809_ & new_n12074_;
  assign new_n12076_ = ~new_n11817_ & ~new_n12075_;
  assign new_n12077_ = ~new_n12073_ & new_n12076_;
  assign new_n12078_ = ~new_n11817_ & ~new_n12077_;
  assign new_n12079_ = \b[20]  & ~new_n11806_;
  assign new_n12080_ = ~new_n11800_ & new_n12079_;
  assign new_n12081_ = ~new_n11808_ & ~new_n12080_;
  assign new_n12082_ = ~new_n12078_ & new_n12081_;
  assign new_n12083_ = ~new_n11808_ & ~new_n12082_;
  assign new_n12084_ = \b[21]  & ~new_n11797_;
  assign new_n12085_ = ~new_n11791_ & new_n12084_;
  assign new_n12086_ = ~new_n11799_ & ~new_n12085_;
  assign new_n12087_ = ~new_n12083_ & new_n12086_;
  assign new_n12088_ = ~new_n11799_ & ~new_n12087_;
  assign new_n12089_ = \b[22]  & ~new_n11788_;
  assign new_n12090_ = ~new_n11782_ & new_n12089_;
  assign new_n12091_ = ~new_n11790_ & ~new_n12090_;
  assign new_n12092_ = ~new_n12088_ & new_n12091_;
  assign new_n12093_ = ~new_n11790_ & ~new_n12092_;
  assign new_n12094_ = \b[23]  & ~new_n11779_;
  assign new_n12095_ = ~new_n11773_ & new_n12094_;
  assign new_n12096_ = ~new_n11781_ & ~new_n12095_;
  assign new_n12097_ = ~new_n12093_ & new_n12096_;
  assign new_n12098_ = ~new_n11781_ & ~new_n12097_;
  assign new_n12099_ = \b[24]  & ~new_n11770_;
  assign new_n12100_ = ~new_n11764_ & new_n12099_;
  assign new_n12101_ = ~new_n11772_ & ~new_n12100_;
  assign new_n12102_ = ~new_n12098_ & new_n12101_;
  assign new_n12103_ = ~new_n11772_ & ~new_n12102_;
  assign new_n12104_ = \b[25]  & ~new_n11761_;
  assign new_n12105_ = ~new_n11755_ & new_n12104_;
  assign new_n12106_ = ~new_n11763_ & ~new_n12105_;
  assign new_n12107_ = ~new_n12103_ & new_n12106_;
  assign new_n12108_ = ~new_n11763_ & ~new_n12107_;
  assign new_n12109_ = \b[26]  & ~new_n11752_;
  assign new_n12110_ = ~new_n11746_ & new_n12109_;
  assign new_n12111_ = ~new_n11754_ & ~new_n12110_;
  assign new_n12112_ = ~new_n12108_ & new_n12111_;
  assign new_n12113_ = ~new_n11754_ & ~new_n12112_;
  assign new_n12114_ = \b[27]  & ~new_n11743_;
  assign new_n12115_ = ~new_n11737_ & new_n12114_;
  assign new_n12116_ = ~new_n11745_ & ~new_n12115_;
  assign new_n12117_ = ~new_n12113_ & new_n12116_;
  assign new_n12118_ = ~new_n11745_ & ~new_n12117_;
  assign new_n12119_ = \b[28]  & ~new_n11734_;
  assign new_n12120_ = ~new_n11728_ & new_n12119_;
  assign new_n12121_ = ~new_n11736_ & ~new_n12120_;
  assign new_n12122_ = ~new_n12118_ & new_n12121_;
  assign new_n12123_ = ~new_n11736_ & ~new_n12122_;
  assign new_n12124_ = \b[29]  & ~new_n11725_;
  assign new_n12125_ = ~new_n11719_ & new_n12124_;
  assign new_n12126_ = ~new_n11727_ & ~new_n12125_;
  assign new_n12127_ = ~new_n12123_ & new_n12126_;
  assign new_n12128_ = ~new_n11727_ & ~new_n12127_;
  assign new_n12129_ = \b[30]  & ~new_n11716_;
  assign new_n12130_ = ~new_n11710_ & new_n12129_;
  assign new_n12131_ = ~new_n11718_ & ~new_n12130_;
  assign new_n12132_ = ~new_n12128_ & new_n12131_;
  assign new_n12133_ = ~new_n11718_ & ~new_n12132_;
  assign new_n12134_ = \b[31]  & ~new_n11707_;
  assign new_n12135_ = ~new_n11701_ & new_n12134_;
  assign new_n12136_ = ~new_n11709_ & ~new_n12135_;
  assign new_n12137_ = ~new_n12133_ & new_n12136_;
  assign new_n12138_ = ~new_n11709_ & ~new_n12137_;
  assign new_n12139_ = \b[32]  & ~new_n11698_;
  assign new_n12140_ = ~new_n11692_ & new_n12139_;
  assign new_n12141_ = ~new_n11700_ & ~new_n12140_;
  assign new_n12142_ = ~new_n12138_ & new_n12141_;
  assign new_n12143_ = ~new_n11700_ & ~new_n12142_;
  assign new_n12144_ = \b[33]  & ~new_n11689_;
  assign new_n12145_ = ~new_n11683_ & new_n12144_;
  assign new_n12146_ = ~new_n11691_ & ~new_n12145_;
  assign new_n12147_ = ~new_n12143_ & new_n12146_;
  assign new_n12148_ = ~new_n11691_ & ~new_n12147_;
  assign new_n12149_ = \b[34]  & ~new_n11680_;
  assign new_n12150_ = ~new_n11674_ & new_n12149_;
  assign new_n12151_ = ~new_n11682_ & ~new_n12150_;
  assign new_n12152_ = ~new_n12148_ & new_n12151_;
  assign new_n12153_ = ~new_n11682_ & ~new_n12152_;
  assign new_n12154_ = \b[35]  & ~new_n11671_;
  assign new_n12155_ = ~new_n11665_ & new_n12154_;
  assign new_n12156_ = ~new_n11673_ & ~new_n12155_;
  assign new_n12157_ = ~new_n12153_ & new_n12156_;
  assign new_n12158_ = ~new_n11673_ & ~new_n12157_;
  assign new_n12159_ = \b[36]  & ~new_n11662_;
  assign new_n12160_ = ~new_n11656_ & new_n12159_;
  assign new_n12161_ = ~new_n11664_ & ~new_n12160_;
  assign new_n12162_ = ~new_n12158_ & new_n12161_;
  assign new_n12163_ = ~new_n11664_ & ~new_n12162_;
  assign new_n12164_ = \b[37]  & ~new_n11653_;
  assign new_n12165_ = ~new_n11647_ & new_n12164_;
  assign new_n12166_ = ~new_n11655_ & ~new_n12165_;
  assign new_n12167_ = ~new_n12163_ & new_n12166_;
  assign new_n12168_ = ~new_n11655_ & ~new_n12167_;
  assign new_n12169_ = \b[38]  & ~new_n11644_;
  assign new_n12170_ = ~new_n11638_ & new_n12169_;
  assign new_n12171_ = ~new_n11646_ & ~new_n12170_;
  assign new_n12172_ = ~new_n12168_ & new_n12171_;
  assign new_n12173_ = ~new_n11646_ & ~new_n12172_;
  assign new_n12174_ = \b[39]  & ~new_n11627_;
  assign new_n12175_ = ~new_n11621_ & new_n12174_;
  assign new_n12176_ = ~new_n11637_ & ~new_n12175_;
  assign new_n12177_ = ~new_n12173_ & new_n12176_;
  assign new_n12178_ = ~new_n11637_ & ~new_n12177_;
  assign new_n12179_ = \b[40]  & ~new_n11629_;
  assign new_n12180_ = ~new_n11634_ & new_n12179_;
  assign new_n12181_ = ~new_n11636_ & ~new_n12180_;
  assign new_n12182_ = ~new_n12178_ & new_n12181_;
  assign new_n12183_ = ~new_n11636_ & ~new_n12182_;
  assign new_n12184_ = new_n408_ & new_n422_;
  assign \quotient[23]  = ~new_n12183_ & new_n12184_;
  assign new_n12186_ = ~new_n11628_ & ~\quotient[23] ;
  assign new_n12187_ = ~new_n11646_ & new_n12176_;
  assign new_n12188_ = ~new_n12172_ & new_n12187_;
  assign new_n12189_ = ~new_n12173_ & ~new_n12176_;
  assign new_n12190_ = ~new_n12188_ & ~new_n12189_;
  assign new_n12191_ = new_n12184_ & ~new_n12190_;
  assign new_n12192_ = ~new_n12183_ & new_n12191_;
  assign new_n12193_ = ~new_n12186_ & ~new_n12192_;
  assign new_n12194_ = ~\b[40]  & ~new_n12193_;
  assign new_n12195_ = ~new_n11645_ & ~\quotient[23] ;
  assign new_n12196_ = ~new_n11655_ & new_n12171_;
  assign new_n12197_ = ~new_n12167_ & new_n12196_;
  assign new_n12198_ = ~new_n12168_ & ~new_n12171_;
  assign new_n12199_ = ~new_n12197_ & ~new_n12198_;
  assign new_n12200_ = new_n12184_ & ~new_n12199_;
  assign new_n12201_ = ~new_n12183_ & new_n12200_;
  assign new_n12202_ = ~new_n12195_ & ~new_n12201_;
  assign new_n12203_ = ~\b[39]  & ~new_n12202_;
  assign new_n12204_ = ~new_n11654_ & ~\quotient[23] ;
  assign new_n12205_ = ~new_n11664_ & new_n12166_;
  assign new_n12206_ = ~new_n12162_ & new_n12205_;
  assign new_n12207_ = ~new_n12163_ & ~new_n12166_;
  assign new_n12208_ = ~new_n12206_ & ~new_n12207_;
  assign new_n12209_ = new_n12184_ & ~new_n12208_;
  assign new_n12210_ = ~new_n12183_ & new_n12209_;
  assign new_n12211_ = ~new_n12204_ & ~new_n12210_;
  assign new_n12212_ = ~\b[38]  & ~new_n12211_;
  assign new_n12213_ = ~new_n11663_ & ~\quotient[23] ;
  assign new_n12214_ = ~new_n11673_ & new_n12161_;
  assign new_n12215_ = ~new_n12157_ & new_n12214_;
  assign new_n12216_ = ~new_n12158_ & ~new_n12161_;
  assign new_n12217_ = ~new_n12215_ & ~new_n12216_;
  assign new_n12218_ = new_n12184_ & ~new_n12217_;
  assign new_n12219_ = ~new_n12183_ & new_n12218_;
  assign new_n12220_ = ~new_n12213_ & ~new_n12219_;
  assign new_n12221_ = ~\b[37]  & ~new_n12220_;
  assign new_n12222_ = ~new_n11672_ & ~\quotient[23] ;
  assign new_n12223_ = ~new_n11682_ & new_n12156_;
  assign new_n12224_ = ~new_n12152_ & new_n12223_;
  assign new_n12225_ = ~new_n12153_ & ~new_n12156_;
  assign new_n12226_ = ~new_n12224_ & ~new_n12225_;
  assign new_n12227_ = new_n12184_ & ~new_n12226_;
  assign new_n12228_ = ~new_n12183_ & new_n12227_;
  assign new_n12229_ = ~new_n12222_ & ~new_n12228_;
  assign new_n12230_ = ~\b[36]  & ~new_n12229_;
  assign new_n12231_ = ~new_n11681_ & ~\quotient[23] ;
  assign new_n12232_ = ~new_n11691_ & new_n12151_;
  assign new_n12233_ = ~new_n12147_ & new_n12232_;
  assign new_n12234_ = ~new_n12148_ & ~new_n12151_;
  assign new_n12235_ = ~new_n12233_ & ~new_n12234_;
  assign new_n12236_ = new_n12184_ & ~new_n12235_;
  assign new_n12237_ = ~new_n12183_ & new_n12236_;
  assign new_n12238_ = ~new_n12231_ & ~new_n12237_;
  assign new_n12239_ = ~\b[35]  & ~new_n12238_;
  assign new_n12240_ = ~new_n11690_ & ~\quotient[23] ;
  assign new_n12241_ = ~new_n11700_ & new_n12146_;
  assign new_n12242_ = ~new_n12142_ & new_n12241_;
  assign new_n12243_ = ~new_n12143_ & ~new_n12146_;
  assign new_n12244_ = ~new_n12242_ & ~new_n12243_;
  assign new_n12245_ = new_n12184_ & ~new_n12244_;
  assign new_n12246_ = ~new_n12183_ & new_n12245_;
  assign new_n12247_ = ~new_n12240_ & ~new_n12246_;
  assign new_n12248_ = ~\b[34]  & ~new_n12247_;
  assign new_n12249_ = ~new_n11699_ & ~\quotient[23] ;
  assign new_n12250_ = ~new_n11709_ & new_n12141_;
  assign new_n12251_ = ~new_n12137_ & new_n12250_;
  assign new_n12252_ = ~new_n12138_ & ~new_n12141_;
  assign new_n12253_ = ~new_n12251_ & ~new_n12252_;
  assign new_n12254_ = new_n12184_ & ~new_n12253_;
  assign new_n12255_ = ~new_n12183_ & new_n12254_;
  assign new_n12256_ = ~new_n12249_ & ~new_n12255_;
  assign new_n12257_ = ~\b[33]  & ~new_n12256_;
  assign new_n12258_ = ~new_n11708_ & ~\quotient[23] ;
  assign new_n12259_ = ~new_n11718_ & new_n12136_;
  assign new_n12260_ = ~new_n12132_ & new_n12259_;
  assign new_n12261_ = ~new_n12133_ & ~new_n12136_;
  assign new_n12262_ = ~new_n12260_ & ~new_n12261_;
  assign new_n12263_ = new_n12184_ & ~new_n12262_;
  assign new_n12264_ = ~new_n12183_ & new_n12263_;
  assign new_n12265_ = ~new_n12258_ & ~new_n12264_;
  assign new_n12266_ = ~\b[32]  & ~new_n12265_;
  assign new_n12267_ = ~new_n11717_ & ~\quotient[23] ;
  assign new_n12268_ = ~new_n11727_ & new_n12131_;
  assign new_n12269_ = ~new_n12127_ & new_n12268_;
  assign new_n12270_ = ~new_n12128_ & ~new_n12131_;
  assign new_n12271_ = ~new_n12269_ & ~new_n12270_;
  assign new_n12272_ = new_n12184_ & ~new_n12271_;
  assign new_n12273_ = ~new_n12183_ & new_n12272_;
  assign new_n12274_ = ~new_n12267_ & ~new_n12273_;
  assign new_n12275_ = ~\b[31]  & ~new_n12274_;
  assign new_n12276_ = ~new_n11726_ & ~\quotient[23] ;
  assign new_n12277_ = ~new_n11736_ & new_n12126_;
  assign new_n12278_ = ~new_n12122_ & new_n12277_;
  assign new_n12279_ = ~new_n12123_ & ~new_n12126_;
  assign new_n12280_ = ~new_n12278_ & ~new_n12279_;
  assign new_n12281_ = new_n12184_ & ~new_n12280_;
  assign new_n12282_ = ~new_n12183_ & new_n12281_;
  assign new_n12283_ = ~new_n12276_ & ~new_n12282_;
  assign new_n12284_ = ~\b[30]  & ~new_n12283_;
  assign new_n12285_ = ~new_n11735_ & ~\quotient[23] ;
  assign new_n12286_ = ~new_n11745_ & new_n12121_;
  assign new_n12287_ = ~new_n12117_ & new_n12286_;
  assign new_n12288_ = ~new_n12118_ & ~new_n12121_;
  assign new_n12289_ = ~new_n12287_ & ~new_n12288_;
  assign new_n12290_ = new_n12184_ & ~new_n12289_;
  assign new_n12291_ = ~new_n12183_ & new_n12290_;
  assign new_n12292_ = ~new_n12285_ & ~new_n12291_;
  assign new_n12293_ = ~\b[29]  & ~new_n12292_;
  assign new_n12294_ = ~new_n11744_ & ~\quotient[23] ;
  assign new_n12295_ = ~new_n11754_ & new_n12116_;
  assign new_n12296_ = ~new_n12112_ & new_n12295_;
  assign new_n12297_ = ~new_n12113_ & ~new_n12116_;
  assign new_n12298_ = ~new_n12296_ & ~new_n12297_;
  assign new_n12299_ = new_n12184_ & ~new_n12298_;
  assign new_n12300_ = ~new_n12183_ & new_n12299_;
  assign new_n12301_ = ~new_n12294_ & ~new_n12300_;
  assign new_n12302_ = ~\b[28]  & ~new_n12301_;
  assign new_n12303_ = ~new_n11753_ & ~\quotient[23] ;
  assign new_n12304_ = ~new_n11763_ & new_n12111_;
  assign new_n12305_ = ~new_n12107_ & new_n12304_;
  assign new_n12306_ = ~new_n12108_ & ~new_n12111_;
  assign new_n12307_ = ~new_n12305_ & ~new_n12306_;
  assign new_n12308_ = new_n12184_ & ~new_n12307_;
  assign new_n12309_ = ~new_n12183_ & new_n12308_;
  assign new_n12310_ = ~new_n12303_ & ~new_n12309_;
  assign new_n12311_ = ~\b[27]  & ~new_n12310_;
  assign new_n12312_ = ~new_n11762_ & ~\quotient[23] ;
  assign new_n12313_ = ~new_n11772_ & new_n12106_;
  assign new_n12314_ = ~new_n12102_ & new_n12313_;
  assign new_n12315_ = ~new_n12103_ & ~new_n12106_;
  assign new_n12316_ = ~new_n12314_ & ~new_n12315_;
  assign new_n12317_ = new_n12184_ & ~new_n12316_;
  assign new_n12318_ = ~new_n12183_ & new_n12317_;
  assign new_n12319_ = ~new_n12312_ & ~new_n12318_;
  assign new_n12320_ = ~\b[26]  & ~new_n12319_;
  assign new_n12321_ = ~new_n11771_ & ~\quotient[23] ;
  assign new_n12322_ = ~new_n11781_ & new_n12101_;
  assign new_n12323_ = ~new_n12097_ & new_n12322_;
  assign new_n12324_ = ~new_n12098_ & ~new_n12101_;
  assign new_n12325_ = ~new_n12323_ & ~new_n12324_;
  assign new_n12326_ = new_n12184_ & ~new_n12325_;
  assign new_n12327_ = ~new_n12183_ & new_n12326_;
  assign new_n12328_ = ~new_n12321_ & ~new_n12327_;
  assign new_n12329_ = ~\b[25]  & ~new_n12328_;
  assign new_n12330_ = ~new_n11780_ & ~\quotient[23] ;
  assign new_n12331_ = ~new_n11790_ & new_n12096_;
  assign new_n12332_ = ~new_n12092_ & new_n12331_;
  assign new_n12333_ = ~new_n12093_ & ~new_n12096_;
  assign new_n12334_ = ~new_n12332_ & ~new_n12333_;
  assign new_n12335_ = new_n12184_ & ~new_n12334_;
  assign new_n12336_ = ~new_n12183_ & new_n12335_;
  assign new_n12337_ = ~new_n12330_ & ~new_n12336_;
  assign new_n12338_ = ~\b[24]  & ~new_n12337_;
  assign new_n12339_ = ~new_n11789_ & ~\quotient[23] ;
  assign new_n12340_ = ~new_n11799_ & new_n12091_;
  assign new_n12341_ = ~new_n12087_ & new_n12340_;
  assign new_n12342_ = ~new_n12088_ & ~new_n12091_;
  assign new_n12343_ = ~new_n12341_ & ~new_n12342_;
  assign new_n12344_ = new_n12184_ & ~new_n12343_;
  assign new_n12345_ = ~new_n12183_ & new_n12344_;
  assign new_n12346_ = ~new_n12339_ & ~new_n12345_;
  assign new_n12347_ = ~\b[23]  & ~new_n12346_;
  assign new_n12348_ = ~new_n11798_ & ~\quotient[23] ;
  assign new_n12349_ = ~new_n11808_ & new_n12086_;
  assign new_n12350_ = ~new_n12082_ & new_n12349_;
  assign new_n12351_ = ~new_n12083_ & ~new_n12086_;
  assign new_n12352_ = ~new_n12350_ & ~new_n12351_;
  assign new_n12353_ = new_n12184_ & ~new_n12352_;
  assign new_n12354_ = ~new_n12183_ & new_n12353_;
  assign new_n12355_ = ~new_n12348_ & ~new_n12354_;
  assign new_n12356_ = ~\b[22]  & ~new_n12355_;
  assign new_n12357_ = ~new_n11807_ & ~\quotient[23] ;
  assign new_n12358_ = ~new_n11817_ & new_n12081_;
  assign new_n12359_ = ~new_n12077_ & new_n12358_;
  assign new_n12360_ = ~new_n12078_ & ~new_n12081_;
  assign new_n12361_ = ~new_n12359_ & ~new_n12360_;
  assign new_n12362_ = new_n12184_ & ~new_n12361_;
  assign new_n12363_ = ~new_n12183_ & new_n12362_;
  assign new_n12364_ = ~new_n12357_ & ~new_n12363_;
  assign new_n12365_ = ~\b[21]  & ~new_n12364_;
  assign new_n12366_ = ~new_n11816_ & ~\quotient[23] ;
  assign new_n12367_ = ~new_n11826_ & new_n12076_;
  assign new_n12368_ = ~new_n12072_ & new_n12367_;
  assign new_n12369_ = ~new_n12073_ & ~new_n12076_;
  assign new_n12370_ = ~new_n12368_ & ~new_n12369_;
  assign new_n12371_ = new_n12184_ & ~new_n12370_;
  assign new_n12372_ = ~new_n12183_ & new_n12371_;
  assign new_n12373_ = ~new_n12366_ & ~new_n12372_;
  assign new_n12374_ = ~\b[20]  & ~new_n12373_;
  assign new_n12375_ = ~new_n11825_ & ~\quotient[23] ;
  assign new_n12376_ = ~new_n11835_ & new_n12071_;
  assign new_n12377_ = ~new_n12067_ & new_n12376_;
  assign new_n12378_ = ~new_n12068_ & ~new_n12071_;
  assign new_n12379_ = ~new_n12377_ & ~new_n12378_;
  assign new_n12380_ = new_n12184_ & ~new_n12379_;
  assign new_n12381_ = ~new_n12183_ & new_n12380_;
  assign new_n12382_ = ~new_n12375_ & ~new_n12381_;
  assign new_n12383_ = ~\b[19]  & ~new_n12382_;
  assign new_n12384_ = ~new_n11834_ & ~\quotient[23] ;
  assign new_n12385_ = ~new_n11844_ & new_n12066_;
  assign new_n12386_ = ~new_n12062_ & new_n12385_;
  assign new_n12387_ = ~new_n12063_ & ~new_n12066_;
  assign new_n12388_ = ~new_n12386_ & ~new_n12387_;
  assign new_n12389_ = new_n12184_ & ~new_n12388_;
  assign new_n12390_ = ~new_n12183_ & new_n12389_;
  assign new_n12391_ = ~new_n12384_ & ~new_n12390_;
  assign new_n12392_ = ~\b[18]  & ~new_n12391_;
  assign new_n12393_ = ~new_n11843_ & ~\quotient[23] ;
  assign new_n12394_ = ~new_n11853_ & new_n12061_;
  assign new_n12395_ = ~new_n12057_ & new_n12394_;
  assign new_n12396_ = ~new_n12058_ & ~new_n12061_;
  assign new_n12397_ = ~new_n12395_ & ~new_n12396_;
  assign new_n12398_ = new_n12184_ & ~new_n12397_;
  assign new_n12399_ = ~new_n12183_ & new_n12398_;
  assign new_n12400_ = ~new_n12393_ & ~new_n12399_;
  assign new_n12401_ = ~\b[17]  & ~new_n12400_;
  assign new_n12402_ = ~new_n11852_ & ~\quotient[23] ;
  assign new_n12403_ = ~new_n11862_ & new_n12056_;
  assign new_n12404_ = ~new_n12052_ & new_n12403_;
  assign new_n12405_ = ~new_n12053_ & ~new_n12056_;
  assign new_n12406_ = ~new_n12404_ & ~new_n12405_;
  assign new_n12407_ = new_n12184_ & ~new_n12406_;
  assign new_n12408_ = ~new_n12183_ & new_n12407_;
  assign new_n12409_ = ~new_n12402_ & ~new_n12408_;
  assign new_n12410_ = ~\b[16]  & ~new_n12409_;
  assign new_n12411_ = ~new_n11861_ & ~\quotient[23] ;
  assign new_n12412_ = ~new_n11871_ & new_n12051_;
  assign new_n12413_ = ~new_n12047_ & new_n12412_;
  assign new_n12414_ = ~new_n12048_ & ~new_n12051_;
  assign new_n12415_ = ~new_n12413_ & ~new_n12414_;
  assign new_n12416_ = new_n12184_ & ~new_n12415_;
  assign new_n12417_ = ~new_n12183_ & new_n12416_;
  assign new_n12418_ = ~new_n12411_ & ~new_n12417_;
  assign new_n12419_ = ~\b[15]  & ~new_n12418_;
  assign new_n12420_ = ~new_n11870_ & ~\quotient[23] ;
  assign new_n12421_ = ~new_n11880_ & new_n12046_;
  assign new_n12422_ = ~new_n12042_ & new_n12421_;
  assign new_n12423_ = ~new_n12043_ & ~new_n12046_;
  assign new_n12424_ = ~new_n12422_ & ~new_n12423_;
  assign new_n12425_ = new_n12184_ & ~new_n12424_;
  assign new_n12426_ = ~new_n12183_ & new_n12425_;
  assign new_n12427_ = ~new_n12420_ & ~new_n12426_;
  assign new_n12428_ = ~\b[14]  & ~new_n12427_;
  assign new_n12429_ = ~new_n11879_ & ~\quotient[23] ;
  assign new_n12430_ = ~new_n11889_ & new_n12041_;
  assign new_n12431_ = ~new_n12037_ & new_n12430_;
  assign new_n12432_ = ~new_n12038_ & ~new_n12041_;
  assign new_n12433_ = ~new_n12431_ & ~new_n12432_;
  assign new_n12434_ = new_n12184_ & ~new_n12433_;
  assign new_n12435_ = ~new_n12183_ & new_n12434_;
  assign new_n12436_ = ~new_n12429_ & ~new_n12435_;
  assign new_n12437_ = ~\b[13]  & ~new_n12436_;
  assign new_n12438_ = ~new_n11888_ & ~\quotient[23] ;
  assign new_n12439_ = ~new_n11898_ & new_n12036_;
  assign new_n12440_ = ~new_n12032_ & new_n12439_;
  assign new_n12441_ = ~new_n12033_ & ~new_n12036_;
  assign new_n12442_ = ~new_n12440_ & ~new_n12441_;
  assign new_n12443_ = new_n12184_ & ~new_n12442_;
  assign new_n12444_ = ~new_n12183_ & new_n12443_;
  assign new_n12445_ = ~new_n12438_ & ~new_n12444_;
  assign new_n12446_ = ~\b[12]  & ~new_n12445_;
  assign new_n12447_ = ~new_n11897_ & ~\quotient[23] ;
  assign new_n12448_ = ~new_n11907_ & new_n12031_;
  assign new_n12449_ = ~new_n12027_ & new_n12448_;
  assign new_n12450_ = ~new_n12028_ & ~new_n12031_;
  assign new_n12451_ = ~new_n12449_ & ~new_n12450_;
  assign new_n12452_ = new_n12184_ & ~new_n12451_;
  assign new_n12453_ = ~new_n12183_ & new_n12452_;
  assign new_n12454_ = ~new_n12447_ & ~new_n12453_;
  assign new_n12455_ = ~\b[11]  & ~new_n12454_;
  assign new_n12456_ = ~new_n11906_ & ~\quotient[23] ;
  assign new_n12457_ = ~new_n11916_ & new_n12026_;
  assign new_n12458_ = ~new_n12022_ & new_n12457_;
  assign new_n12459_ = ~new_n12023_ & ~new_n12026_;
  assign new_n12460_ = ~new_n12458_ & ~new_n12459_;
  assign new_n12461_ = new_n12184_ & ~new_n12460_;
  assign new_n12462_ = ~new_n12183_ & new_n12461_;
  assign new_n12463_ = ~new_n12456_ & ~new_n12462_;
  assign new_n12464_ = ~\b[10]  & ~new_n12463_;
  assign new_n12465_ = ~new_n11915_ & ~\quotient[23] ;
  assign new_n12466_ = ~new_n11925_ & new_n12021_;
  assign new_n12467_ = ~new_n12017_ & new_n12466_;
  assign new_n12468_ = ~new_n12018_ & ~new_n12021_;
  assign new_n12469_ = ~new_n12467_ & ~new_n12468_;
  assign new_n12470_ = new_n12184_ & ~new_n12469_;
  assign new_n12471_ = ~new_n12183_ & new_n12470_;
  assign new_n12472_ = ~new_n12465_ & ~new_n12471_;
  assign new_n12473_ = ~\b[9]  & ~new_n12472_;
  assign new_n12474_ = ~new_n11924_ & ~\quotient[23] ;
  assign new_n12475_ = ~new_n11934_ & new_n12016_;
  assign new_n12476_ = ~new_n12012_ & new_n12475_;
  assign new_n12477_ = ~new_n12013_ & ~new_n12016_;
  assign new_n12478_ = ~new_n12476_ & ~new_n12477_;
  assign new_n12479_ = new_n12184_ & ~new_n12478_;
  assign new_n12480_ = ~new_n12183_ & new_n12479_;
  assign new_n12481_ = ~new_n12474_ & ~new_n12480_;
  assign new_n12482_ = ~\b[8]  & ~new_n12481_;
  assign new_n12483_ = ~new_n11933_ & ~\quotient[23] ;
  assign new_n12484_ = ~new_n11943_ & new_n12011_;
  assign new_n12485_ = ~new_n12007_ & new_n12484_;
  assign new_n12486_ = ~new_n12008_ & ~new_n12011_;
  assign new_n12487_ = ~new_n12485_ & ~new_n12486_;
  assign new_n12488_ = new_n12184_ & ~new_n12487_;
  assign new_n12489_ = ~new_n12183_ & new_n12488_;
  assign new_n12490_ = ~new_n12483_ & ~new_n12489_;
  assign new_n12491_ = ~\b[7]  & ~new_n12490_;
  assign new_n12492_ = ~new_n11942_ & ~\quotient[23] ;
  assign new_n12493_ = ~new_n11952_ & new_n12006_;
  assign new_n12494_ = ~new_n12002_ & new_n12493_;
  assign new_n12495_ = ~new_n12003_ & ~new_n12006_;
  assign new_n12496_ = ~new_n12494_ & ~new_n12495_;
  assign new_n12497_ = new_n12184_ & ~new_n12496_;
  assign new_n12498_ = ~new_n12183_ & new_n12497_;
  assign new_n12499_ = ~new_n12492_ & ~new_n12498_;
  assign new_n12500_ = ~\b[6]  & ~new_n12499_;
  assign new_n12501_ = ~new_n11951_ & ~\quotient[23] ;
  assign new_n12502_ = ~new_n11961_ & new_n12001_;
  assign new_n12503_ = ~new_n11997_ & new_n12502_;
  assign new_n12504_ = ~new_n11998_ & ~new_n12001_;
  assign new_n12505_ = ~new_n12503_ & ~new_n12504_;
  assign new_n12506_ = new_n12184_ & ~new_n12505_;
  assign new_n12507_ = ~new_n12183_ & new_n12506_;
  assign new_n12508_ = ~new_n12501_ & ~new_n12507_;
  assign new_n12509_ = ~\b[5]  & ~new_n12508_;
  assign new_n12510_ = ~new_n11960_ & ~\quotient[23] ;
  assign new_n12511_ = ~new_n11969_ & new_n11996_;
  assign new_n12512_ = ~new_n11992_ & new_n12511_;
  assign new_n12513_ = ~new_n11993_ & ~new_n11996_;
  assign new_n12514_ = ~new_n12512_ & ~new_n12513_;
  assign new_n12515_ = new_n12184_ & ~new_n12514_;
  assign new_n12516_ = ~new_n12183_ & new_n12515_;
  assign new_n12517_ = ~new_n12510_ & ~new_n12516_;
  assign new_n12518_ = ~\b[4]  & ~new_n12517_;
  assign new_n12519_ = ~new_n11968_ & ~\quotient[23] ;
  assign new_n12520_ = ~new_n11987_ & new_n11991_;
  assign new_n12521_ = ~new_n11986_ & new_n12520_;
  assign new_n12522_ = ~new_n11988_ & ~new_n11991_;
  assign new_n12523_ = ~new_n12521_ & ~new_n12522_;
  assign new_n12524_ = new_n12184_ & ~new_n12523_;
  assign new_n12525_ = ~new_n12183_ & new_n12524_;
  assign new_n12526_ = ~new_n12519_ & ~new_n12525_;
  assign new_n12527_ = ~\b[3]  & ~new_n12526_;
  assign new_n12528_ = ~new_n11980_ & ~\quotient[23] ;
  assign new_n12529_ = ~new_n11983_ & new_n11985_;
  assign new_n12530_ = ~new_n11981_ & new_n12529_;
  assign new_n12531_ = new_n12184_ & ~new_n12530_;
  assign new_n12532_ = ~new_n11986_ & new_n12531_;
  assign new_n12533_ = ~new_n12183_ & new_n12532_;
  assign new_n12534_ = ~new_n12528_ & ~new_n12533_;
  assign new_n12535_ = ~\b[2]  & ~new_n12534_;
  assign new_n12536_ = \b[0]  & ~\b[41] ;
  assign new_n12537_ = new_n290_ & new_n12536_;
  assign new_n12538_ = new_n301_ & new_n12537_;
  assign new_n12539_ = new_n338_ & new_n12538_;
  assign new_n12540_ = ~new_n12183_ & new_n12539_;
  assign new_n12541_ = \a[23]  & ~new_n12540_;
  assign new_n12542_ = new_n421_ & new_n11985_;
  assign new_n12543_ = new_n597_ & new_n12542_;
  assign new_n12544_ = new_n595_ & new_n12543_;
  assign new_n12545_ = ~new_n12183_ & new_n12544_;
  assign new_n12546_ = ~new_n12541_ & ~new_n12545_;
  assign new_n12547_ = \b[1]  & ~new_n12546_;
  assign new_n12548_ = ~\b[1]  & ~new_n12545_;
  assign new_n12549_ = ~new_n12541_ & new_n12548_;
  assign new_n12550_ = ~new_n12547_ & ~new_n12549_;
  assign new_n12551_ = ~\a[22]  & \b[0] ;
  assign new_n12552_ = ~new_n12550_ & ~new_n12551_;
  assign new_n12553_ = ~\b[1]  & ~new_n12546_;
  assign new_n12554_ = ~new_n12552_ & ~new_n12553_;
  assign new_n12555_ = \b[2]  & ~new_n12533_;
  assign new_n12556_ = ~new_n12528_ & new_n12555_;
  assign new_n12557_ = ~new_n12535_ & ~new_n12556_;
  assign new_n12558_ = ~new_n12554_ & new_n12557_;
  assign new_n12559_ = ~new_n12535_ & ~new_n12558_;
  assign new_n12560_ = \b[3]  & ~new_n12525_;
  assign new_n12561_ = ~new_n12519_ & new_n12560_;
  assign new_n12562_ = ~new_n12527_ & ~new_n12561_;
  assign new_n12563_ = ~new_n12559_ & new_n12562_;
  assign new_n12564_ = ~new_n12527_ & ~new_n12563_;
  assign new_n12565_ = \b[4]  & ~new_n12516_;
  assign new_n12566_ = ~new_n12510_ & new_n12565_;
  assign new_n12567_ = ~new_n12518_ & ~new_n12566_;
  assign new_n12568_ = ~new_n12564_ & new_n12567_;
  assign new_n12569_ = ~new_n12518_ & ~new_n12568_;
  assign new_n12570_ = \b[5]  & ~new_n12507_;
  assign new_n12571_ = ~new_n12501_ & new_n12570_;
  assign new_n12572_ = ~new_n12509_ & ~new_n12571_;
  assign new_n12573_ = ~new_n12569_ & new_n12572_;
  assign new_n12574_ = ~new_n12509_ & ~new_n12573_;
  assign new_n12575_ = \b[6]  & ~new_n12498_;
  assign new_n12576_ = ~new_n12492_ & new_n12575_;
  assign new_n12577_ = ~new_n12500_ & ~new_n12576_;
  assign new_n12578_ = ~new_n12574_ & new_n12577_;
  assign new_n12579_ = ~new_n12500_ & ~new_n12578_;
  assign new_n12580_ = \b[7]  & ~new_n12489_;
  assign new_n12581_ = ~new_n12483_ & new_n12580_;
  assign new_n12582_ = ~new_n12491_ & ~new_n12581_;
  assign new_n12583_ = ~new_n12579_ & new_n12582_;
  assign new_n12584_ = ~new_n12491_ & ~new_n12583_;
  assign new_n12585_ = \b[8]  & ~new_n12480_;
  assign new_n12586_ = ~new_n12474_ & new_n12585_;
  assign new_n12587_ = ~new_n12482_ & ~new_n12586_;
  assign new_n12588_ = ~new_n12584_ & new_n12587_;
  assign new_n12589_ = ~new_n12482_ & ~new_n12588_;
  assign new_n12590_ = \b[9]  & ~new_n12471_;
  assign new_n12591_ = ~new_n12465_ & new_n12590_;
  assign new_n12592_ = ~new_n12473_ & ~new_n12591_;
  assign new_n12593_ = ~new_n12589_ & new_n12592_;
  assign new_n12594_ = ~new_n12473_ & ~new_n12593_;
  assign new_n12595_ = \b[10]  & ~new_n12462_;
  assign new_n12596_ = ~new_n12456_ & new_n12595_;
  assign new_n12597_ = ~new_n12464_ & ~new_n12596_;
  assign new_n12598_ = ~new_n12594_ & new_n12597_;
  assign new_n12599_ = ~new_n12464_ & ~new_n12598_;
  assign new_n12600_ = \b[11]  & ~new_n12453_;
  assign new_n12601_ = ~new_n12447_ & new_n12600_;
  assign new_n12602_ = ~new_n12455_ & ~new_n12601_;
  assign new_n12603_ = ~new_n12599_ & new_n12602_;
  assign new_n12604_ = ~new_n12455_ & ~new_n12603_;
  assign new_n12605_ = \b[12]  & ~new_n12444_;
  assign new_n12606_ = ~new_n12438_ & new_n12605_;
  assign new_n12607_ = ~new_n12446_ & ~new_n12606_;
  assign new_n12608_ = ~new_n12604_ & new_n12607_;
  assign new_n12609_ = ~new_n12446_ & ~new_n12608_;
  assign new_n12610_ = \b[13]  & ~new_n12435_;
  assign new_n12611_ = ~new_n12429_ & new_n12610_;
  assign new_n12612_ = ~new_n12437_ & ~new_n12611_;
  assign new_n12613_ = ~new_n12609_ & new_n12612_;
  assign new_n12614_ = ~new_n12437_ & ~new_n12613_;
  assign new_n12615_ = \b[14]  & ~new_n12426_;
  assign new_n12616_ = ~new_n12420_ & new_n12615_;
  assign new_n12617_ = ~new_n12428_ & ~new_n12616_;
  assign new_n12618_ = ~new_n12614_ & new_n12617_;
  assign new_n12619_ = ~new_n12428_ & ~new_n12618_;
  assign new_n12620_ = \b[15]  & ~new_n12417_;
  assign new_n12621_ = ~new_n12411_ & new_n12620_;
  assign new_n12622_ = ~new_n12419_ & ~new_n12621_;
  assign new_n12623_ = ~new_n12619_ & new_n12622_;
  assign new_n12624_ = ~new_n12419_ & ~new_n12623_;
  assign new_n12625_ = \b[16]  & ~new_n12408_;
  assign new_n12626_ = ~new_n12402_ & new_n12625_;
  assign new_n12627_ = ~new_n12410_ & ~new_n12626_;
  assign new_n12628_ = ~new_n12624_ & new_n12627_;
  assign new_n12629_ = ~new_n12410_ & ~new_n12628_;
  assign new_n12630_ = \b[17]  & ~new_n12399_;
  assign new_n12631_ = ~new_n12393_ & new_n12630_;
  assign new_n12632_ = ~new_n12401_ & ~new_n12631_;
  assign new_n12633_ = ~new_n12629_ & new_n12632_;
  assign new_n12634_ = ~new_n12401_ & ~new_n12633_;
  assign new_n12635_ = \b[18]  & ~new_n12390_;
  assign new_n12636_ = ~new_n12384_ & new_n12635_;
  assign new_n12637_ = ~new_n12392_ & ~new_n12636_;
  assign new_n12638_ = ~new_n12634_ & new_n12637_;
  assign new_n12639_ = ~new_n12392_ & ~new_n12638_;
  assign new_n12640_ = \b[19]  & ~new_n12381_;
  assign new_n12641_ = ~new_n12375_ & new_n12640_;
  assign new_n12642_ = ~new_n12383_ & ~new_n12641_;
  assign new_n12643_ = ~new_n12639_ & new_n12642_;
  assign new_n12644_ = ~new_n12383_ & ~new_n12643_;
  assign new_n12645_ = \b[20]  & ~new_n12372_;
  assign new_n12646_ = ~new_n12366_ & new_n12645_;
  assign new_n12647_ = ~new_n12374_ & ~new_n12646_;
  assign new_n12648_ = ~new_n12644_ & new_n12647_;
  assign new_n12649_ = ~new_n12374_ & ~new_n12648_;
  assign new_n12650_ = \b[21]  & ~new_n12363_;
  assign new_n12651_ = ~new_n12357_ & new_n12650_;
  assign new_n12652_ = ~new_n12365_ & ~new_n12651_;
  assign new_n12653_ = ~new_n12649_ & new_n12652_;
  assign new_n12654_ = ~new_n12365_ & ~new_n12653_;
  assign new_n12655_ = \b[22]  & ~new_n12354_;
  assign new_n12656_ = ~new_n12348_ & new_n12655_;
  assign new_n12657_ = ~new_n12356_ & ~new_n12656_;
  assign new_n12658_ = ~new_n12654_ & new_n12657_;
  assign new_n12659_ = ~new_n12356_ & ~new_n12658_;
  assign new_n12660_ = \b[23]  & ~new_n12345_;
  assign new_n12661_ = ~new_n12339_ & new_n12660_;
  assign new_n12662_ = ~new_n12347_ & ~new_n12661_;
  assign new_n12663_ = ~new_n12659_ & new_n12662_;
  assign new_n12664_ = ~new_n12347_ & ~new_n12663_;
  assign new_n12665_ = \b[24]  & ~new_n12336_;
  assign new_n12666_ = ~new_n12330_ & new_n12665_;
  assign new_n12667_ = ~new_n12338_ & ~new_n12666_;
  assign new_n12668_ = ~new_n12664_ & new_n12667_;
  assign new_n12669_ = ~new_n12338_ & ~new_n12668_;
  assign new_n12670_ = \b[25]  & ~new_n12327_;
  assign new_n12671_ = ~new_n12321_ & new_n12670_;
  assign new_n12672_ = ~new_n12329_ & ~new_n12671_;
  assign new_n12673_ = ~new_n12669_ & new_n12672_;
  assign new_n12674_ = ~new_n12329_ & ~new_n12673_;
  assign new_n12675_ = \b[26]  & ~new_n12318_;
  assign new_n12676_ = ~new_n12312_ & new_n12675_;
  assign new_n12677_ = ~new_n12320_ & ~new_n12676_;
  assign new_n12678_ = ~new_n12674_ & new_n12677_;
  assign new_n12679_ = ~new_n12320_ & ~new_n12678_;
  assign new_n12680_ = \b[27]  & ~new_n12309_;
  assign new_n12681_ = ~new_n12303_ & new_n12680_;
  assign new_n12682_ = ~new_n12311_ & ~new_n12681_;
  assign new_n12683_ = ~new_n12679_ & new_n12682_;
  assign new_n12684_ = ~new_n12311_ & ~new_n12683_;
  assign new_n12685_ = \b[28]  & ~new_n12300_;
  assign new_n12686_ = ~new_n12294_ & new_n12685_;
  assign new_n12687_ = ~new_n12302_ & ~new_n12686_;
  assign new_n12688_ = ~new_n12684_ & new_n12687_;
  assign new_n12689_ = ~new_n12302_ & ~new_n12688_;
  assign new_n12690_ = \b[29]  & ~new_n12291_;
  assign new_n12691_ = ~new_n12285_ & new_n12690_;
  assign new_n12692_ = ~new_n12293_ & ~new_n12691_;
  assign new_n12693_ = ~new_n12689_ & new_n12692_;
  assign new_n12694_ = ~new_n12293_ & ~new_n12693_;
  assign new_n12695_ = \b[30]  & ~new_n12282_;
  assign new_n12696_ = ~new_n12276_ & new_n12695_;
  assign new_n12697_ = ~new_n12284_ & ~new_n12696_;
  assign new_n12698_ = ~new_n12694_ & new_n12697_;
  assign new_n12699_ = ~new_n12284_ & ~new_n12698_;
  assign new_n12700_ = \b[31]  & ~new_n12273_;
  assign new_n12701_ = ~new_n12267_ & new_n12700_;
  assign new_n12702_ = ~new_n12275_ & ~new_n12701_;
  assign new_n12703_ = ~new_n12699_ & new_n12702_;
  assign new_n12704_ = ~new_n12275_ & ~new_n12703_;
  assign new_n12705_ = \b[32]  & ~new_n12264_;
  assign new_n12706_ = ~new_n12258_ & new_n12705_;
  assign new_n12707_ = ~new_n12266_ & ~new_n12706_;
  assign new_n12708_ = ~new_n12704_ & new_n12707_;
  assign new_n12709_ = ~new_n12266_ & ~new_n12708_;
  assign new_n12710_ = \b[33]  & ~new_n12255_;
  assign new_n12711_ = ~new_n12249_ & new_n12710_;
  assign new_n12712_ = ~new_n12257_ & ~new_n12711_;
  assign new_n12713_ = ~new_n12709_ & new_n12712_;
  assign new_n12714_ = ~new_n12257_ & ~new_n12713_;
  assign new_n12715_ = \b[34]  & ~new_n12246_;
  assign new_n12716_ = ~new_n12240_ & new_n12715_;
  assign new_n12717_ = ~new_n12248_ & ~new_n12716_;
  assign new_n12718_ = ~new_n12714_ & new_n12717_;
  assign new_n12719_ = ~new_n12248_ & ~new_n12718_;
  assign new_n12720_ = \b[35]  & ~new_n12237_;
  assign new_n12721_ = ~new_n12231_ & new_n12720_;
  assign new_n12722_ = ~new_n12239_ & ~new_n12721_;
  assign new_n12723_ = ~new_n12719_ & new_n12722_;
  assign new_n12724_ = ~new_n12239_ & ~new_n12723_;
  assign new_n12725_ = \b[36]  & ~new_n12228_;
  assign new_n12726_ = ~new_n12222_ & new_n12725_;
  assign new_n12727_ = ~new_n12230_ & ~new_n12726_;
  assign new_n12728_ = ~new_n12724_ & new_n12727_;
  assign new_n12729_ = ~new_n12230_ & ~new_n12728_;
  assign new_n12730_ = \b[37]  & ~new_n12219_;
  assign new_n12731_ = ~new_n12213_ & new_n12730_;
  assign new_n12732_ = ~new_n12221_ & ~new_n12731_;
  assign new_n12733_ = ~new_n12729_ & new_n12732_;
  assign new_n12734_ = ~new_n12221_ & ~new_n12733_;
  assign new_n12735_ = \b[38]  & ~new_n12210_;
  assign new_n12736_ = ~new_n12204_ & new_n12735_;
  assign new_n12737_ = ~new_n12212_ & ~new_n12736_;
  assign new_n12738_ = ~new_n12734_ & new_n12737_;
  assign new_n12739_ = ~new_n12212_ & ~new_n12738_;
  assign new_n12740_ = \b[39]  & ~new_n12201_;
  assign new_n12741_ = ~new_n12195_ & new_n12740_;
  assign new_n12742_ = ~new_n12203_ & ~new_n12741_;
  assign new_n12743_ = ~new_n12739_ & new_n12742_;
  assign new_n12744_ = ~new_n12203_ & ~new_n12743_;
  assign new_n12745_ = \b[40]  & ~new_n12192_;
  assign new_n12746_ = ~new_n12186_ & new_n12745_;
  assign new_n12747_ = ~new_n12194_ & ~new_n12746_;
  assign new_n12748_ = ~new_n12744_ & new_n12747_;
  assign new_n12749_ = ~new_n12194_ & ~new_n12748_;
  assign new_n12750_ = ~new_n11635_ & ~\quotient[23] ;
  assign new_n12751_ = ~new_n11637_ & new_n12181_;
  assign new_n12752_ = ~new_n12177_ & new_n12751_;
  assign new_n12753_ = ~new_n12178_ & ~new_n12181_;
  assign new_n12754_ = ~new_n12752_ & ~new_n12753_;
  assign new_n12755_ = \quotient[23]  & ~new_n12754_;
  assign new_n12756_ = ~new_n12750_ & ~new_n12755_;
  assign new_n12757_ = ~\b[41]  & ~new_n12756_;
  assign new_n12758_ = \b[41]  & ~new_n12750_;
  assign new_n12759_ = ~new_n12755_ & new_n12758_;
  assign new_n12760_ = new_n290_ & new_n301_;
  assign new_n12761_ = new_n338_ & new_n12760_;
  assign new_n12762_ = ~new_n12759_ & new_n12761_;
  assign new_n12763_ = ~new_n12757_ & new_n12762_;
  assign new_n12764_ = ~new_n12749_ & new_n12763_;
  assign new_n12765_ = new_n12184_ & ~new_n12756_;
  assign \quotient[22]  = new_n12764_ | new_n12765_;
  assign new_n12767_ = ~new_n12203_ & new_n12747_;
  assign new_n12768_ = ~new_n12743_ & new_n12767_;
  assign new_n12769_ = ~new_n12744_ & ~new_n12747_;
  assign new_n12770_ = ~new_n12768_ & ~new_n12769_;
  assign new_n12771_ = \quotient[22]  & ~new_n12770_;
  assign new_n12772_ = ~new_n12193_ & ~new_n12765_;
  assign new_n12773_ = ~new_n12764_ & new_n12772_;
  assign new_n12774_ = ~new_n12771_ & ~new_n12773_;
  assign new_n12775_ = ~new_n12194_ & ~new_n12759_;
  assign new_n12776_ = ~new_n12757_ & new_n12775_;
  assign new_n12777_ = ~new_n12748_ & new_n12776_;
  assign new_n12778_ = ~new_n12757_ & ~new_n12759_;
  assign new_n12779_ = ~new_n12749_ & ~new_n12778_;
  assign new_n12780_ = ~new_n12777_ & ~new_n12779_;
  assign new_n12781_ = \quotient[22]  & ~new_n12780_;
  assign new_n12782_ = ~new_n12756_ & ~new_n12765_;
  assign new_n12783_ = ~new_n12764_ & new_n12782_;
  assign new_n12784_ = ~new_n12781_ & ~new_n12783_;
  assign new_n12785_ = ~\b[42]  & ~new_n12784_;
  assign new_n12786_ = ~\b[41]  & ~new_n12774_;
  assign new_n12787_ = ~new_n12212_ & new_n12742_;
  assign new_n12788_ = ~new_n12738_ & new_n12787_;
  assign new_n12789_ = ~new_n12739_ & ~new_n12742_;
  assign new_n12790_ = ~new_n12788_ & ~new_n12789_;
  assign new_n12791_ = \quotient[22]  & ~new_n12790_;
  assign new_n12792_ = ~new_n12202_ & ~new_n12765_;
  assign new_n12793_ = ~new_n12764_ & new_n12792_;
  assign new_n12794_ = ~new_n12791_ & ~new_n12793_;
  assign new_n12795_ = ~\b[40]  & ~new_n12794_;
  assign new_n12796_ = ~new_n12221_ & new_n12737_;
  assign new_n12797_ = ~new_n12733_ & new_n12796_;
  assign new_n12798_ = ~new_n12734_ & ~new_n12737_;
  assign new_n12799_ = ~new_n12797_ & ~new_n12798_;
  assign new_n12800_ = \quotient[22]  & ~new_n12799_;
  assign new_n12801_ = ~new_n12211_ & ~new_n12765_;
  assign new_n12802_ = ~new_n12764_ & new_n12801_;
  assign new_n12803_ = ~new_n12800_ & ~new_n12802_;
  assign new_n12804_ = ~\b[39]  & ~new_n12803_;
  assign new_n12805_ = ~new_n12230_ & new_n12732_;
  assign new_n12806_ = ~new_n12728_ & new_n12805_;
  assign new_n12807_ = ~new_n12729_ & ~new_n12732_;
  assign new_n12808_ = ~new_n12806_ & ~new_n12807_;
  assign new_n12809_ = \quotient[22]  & ~new_n12808_;
  assign new_n12810_ = ~new_n12220_ & ~new_n12765_;
  assign new_n12811_ = ~new_n12764_ & new_n12810_;
  assign new_n12812_ = ~new_n12809_ & ~new_n12811_;
  assign new_n12813_ = ~\b[38]  & ~new_n12812_;
  assign new_n12814_ = ~new_n12239_ & new_n12727_;
  assign new_n12815_ = ~new_n12723_ & new_n12814_;
  assign new_n12816_ = ~new_n12724_ & ~new_n12727_;
  assign new_n12817_ = ~new_n12815_ & ~new_n12816_;
  assign new_n12818_ = \quotient[22]  & ~new_n12817_;
  assign new_n12819_ = ~new_n12229_ & ~new_n12765_;
  assign new_n12820_ = ~new_n12764_ & new_n12819_;
  assign new_n12821_ = ~new_n12818_ & ~new_n12820_;
  assign new_n12822_ = ~\b[37]  & ~new_n12821_;
  assign new_n12823_ = ~new_n12248_ & new_n12722_;
  assign new_n12824_ = ~new_n12718_ & new_n12823_;
  assign new_n12825_ = ~new_n12719_ & ~new_n12722_;
  assign new_n12826_ = ~new_n12824_ & ~new_n12825_;
  assign new_n12827_ = \quotient[22]  & ~new_n12826_;
  assign new_n12828_ = ~new_n12238_ & ~new_n12765_;
  assign new_n12829_ = ~new_n12764_ & new_n12828_;
  assign new_n12830_ = ~new_n12827_ & ~new_n12829_;
  assign new_n12831_ = ~\b[36]  & ~new_n12830_;
  assign new_n12832_ = ~new_n12257_ & new_n12717_;
  assign new_n12833_ = ~new_n12713_ & new_n12832_;
  assign new_n12834_ = ~new_n12714_ & ~new_n12717_;
  assign new_n12835_ = ~new_n12833_ & ~new_n12834_;
  assign new_n12836_ = \quotient[22]  & ~new_n12835_;
  assign new_n12837_ = ~new_n12247_ & ~new_n12765_;
  assign new_n12838_ = ~new_n12764_ & new_n12837_;
  assign new_n12839_ = ~new_n12836_ & ~new_n12838_;
  assign new_n12840_ = ~\b[35]  & ~new_n12839_;
  assign new_n12841_ = ~new_n12266_ & new_n12712_;
  assign new_n12842_ = ~new_n12708_ & new_n12841_;
  assign new_n12843_ = ~new_n12709_ & ~new_n12712_;
  assign new_n12844_ = ~new_n12842_ & ~new_n12843_;
  assign new_n12845_ = \quotient[22]  & ~new_n12844_;
  assign new_n12846_ = ~new_n12256_ & ~new_n12765_;
  assign new_n12847_ = ~new_n12764_ & new_n12846_;
  assign new_n12848_ = ~new_n12845_ & ~new_n12847_;
  assign new_n12849_ = ~\b[34]  & ~new_n12848_;
  assign new_n12850_ = ~new_n12275_ & new_n12707_;
  assign new_n12851_ = ~new_n12703_ & new_n12850_;
  assign new_n12852_ = ~new_n12704_ & ~new_n12707_;
  assign new_n12853_ = ~new_n12851_ & ~new_n12852_;
  assign new_n12854_ = \quotient[22]  & ~new_n12853_;
  assign new_n12855_ = ~new_n12265_ & ~new_n12765_;
  assign new_n12856_ = ~new_n12764_ & new_n12855_;
  assign new_n12857_ = ~new_n12854_ & ~new_n12856_;
  assign new_n12858_ = ~\b[33]  & ~new_n12857_;
  assign new_n12859_ = ~new_n12284_ & new_n12702_;
  assign new_n12860_ = ~new_n12698_ & new_n12859_;
  assign new_n12861_ = ~new_n12699_ & ~new_n12702_;
  assign new_n12862_ = ~new_n12860_ & ~new_n12861_;
  assign new_n12863_ = \quotient[22]  & ~new_n12862_;
  assign new_n12864_ = ~new_n12274_ & ~new_n12765_;
  assign new_n12865_ = ~new_n12764_ & new_n12864_;
  assign new_n12866_ = ~new_n12863_ & ~new_n12865_;
  assign new_n12867_ = ~\b[32]  & ~new_n12866_;
  assign new_n12868_ = ~new_n12293_ & new_n12697_;
  assign new_n12869_ = ~new_n12693_ & new_n12868_;
  assign new_n12870_ = ~new_n12694_ & ~new_n12697_;
  assign new_n12871_ = ~new_n12869_ & ~new_n12870_;
  assign new_n12872_ = \quotient[22]  & ~new_n12871_;
  assign new_n12873_ = ~new_n12283_ & ~new_n12765_;
  assign new_n12874_ = ~new_n12764_ & new_n12873_;
  assign new_n12875_ = ~new_n12872_ & ~new_n12874_;
  assign new_n12876_ = ~\b[31]  & ~new_n12875_;
  assign new_n12877_ = ~new_n12302_ & new_n12692_;
  assign new_n12878_ = ~new_n12688_ & new_n12877_;
  assign new_n12879_ = ~new_n12689_ & ~new_n12692_;
  assign new_n12880_ = ~new_n12878_ & ~new_n12879_;
  assign new_n12881_ = \quotient[22]  & ~new_n12880_;
  assign new_n12882_ = ~new_n12292_ & ~new_n12765_;
  assign new_n12883_ = ~new_n12764_ & new_n12882_;
  assign new_n12884_ = ~new_n12881_ & ~new_n12883_;
  assign new_n12885_ = ~\b[30]  & ~new_n12884_;
  assign new_n12886_ = ~new_n12311_ & new_n12687_;
  assign new_n12887_ = ~new_n12683_ & new_n12886_;
  assign new_n12888_ = ~new_n12684_ & ~new_n12687_;
  assign new_n12889_ = ~new_n12887_ & ~new_n12888_;
  assign new_n12890_ = \quotient[22]  & ~new_n12889_;
  assign new_n12891_ = ~new_n12301_ & ~new_n12765_;
  assign new_n12892_ = ~new_n12764_ & new_n12891_;
  assign new_n12893_ = ~new_n12890_ & ~new_n12892_;
  assign new_n12894_ = ~\b[29]  & ~new_n12893_;
  assign new_n12895_ = ~new_n12320_ & new_n12682_;
  assign new_n12896_ = ~new_n12678_ & new_n12895_;
  assign new_n12897_ = ~new_n12679_ & ~new_n12682_;
  assign new_n12898_ = ~new_n12896_ & ~new_n12897_;
  assign new_n12899_ = \quotient[22]  & ~new_n12898_;
  assign new_n12900_ = ~new_n12310_ & ~new_n12765_;
  assign new_n12901_ = ~new_n12764_ & new_n12900_;
  assign new_n12902_ = ~new_n12899_ & ~new_n12901_;
  assign new_n12903_ = ~\b[28]  & ~new_n12902_;
  assign new_n12904_ = ~new_n12329_ & new_n12677_;
  assign new_n12905_ = ~new_n12673_ & new_n12904_;
  assign new_n12906_ = ~new_n12674_ & ~new_n12677_;
  assign new_n12907_ = ~new_n12905_ & ~new_n12906_;
  assign new_n12908_ = \quotient[22]  & ~new_n12907_;
  assign new_n12909_ = ~new_n12319_ & ~new_n12765_;
  assign new_n12910_ = ~new_n12764_ & new_n12909_;
  assign new_n12911_ = ~new_n12908_ & ~new_n12910_;
  assign new_n12912_ = ~\b[27]  & ~new_n12911_;
  assign new_n12913_ = ~new_n12338_ & new_n12672_;
  assign new_n12914_ = ~new_n12668_ & new_n12913_;
  assign new_n12915_ = ~new_n12669_ & ~new_n12672_;
  assign new_n12916_ = ~new_n12914_ & ~new_n12915_;
  assign new_n12917_ = \quotient[22]  & ~new_n12916_;
  assign new_n12918_ = ~new_n12328_ & ~new_n12765_;
  assign new_n12919_ = ~new_n12764_ & new_n12918_;
  assign new_n12920_ = ~new_n12917_ & ~new_n12919_;
  assign new_n12921_ = ~\b[26]  & ~new_n12920_;
  assign new_n12922_ = ~new_n12347_ & new_n12667_;
  assign new_n12923_ = ~new_n12663_ & new_n12922_;
  assign new_n12924_ = ~new_n12664_ & ~new_n12667_;
  assign new_n12925_ = ~new_n12923_ & ~new_n12924_;
  assign new_n12926_ = \quotient[22]  & ~new_n12925_;
  assign new_n12927_ = ~new_n12337_ & ~new_n12765_;
  assign new_n12928_ = ~new_n12764_ & new_n12927_;
  assign new_n12929_ = ~new_n12926_ & ~new_n12928_;
  assign new_n12930_ = ~\b[25]  & ~new_n12929_;
  assign new_n12931_ = ~new_n12356_ & new_n12662_;
  assign new_n12932_ = ~new_n12658_ & new_n12931_;
  assign new_n12933_ = ~new_n12659_ & ~new_n12662_;
  assign new_n12934_ = ~new_n12932_ & ~new_n12933_;
  assign new_n12935_ = \quotient[22]  & ~new_n12934_;
  assign new_n12936_ = ~new_n12346_ & ~new_n12765_;
  assign new_n12937_ = ~new_n12764_ & new_n12936_;
  assign new_n12938_ = ~new_n12935_ & ~new_n12937_;
  assign new_n12939_ = ~\b[24]  & ~new_n12938_;
  assign new_n12940_ = ~new_n12365_ & new_n12657_;
  assign new_n12941_ = ~new_n12653_ & new_n12940_;
  assign new_n12942_ = ~new_n12654_ & ~new_n12657_;
  assign new_n12943_ = ~new_n12941_ & ~new_n12942_;
  assign new_n12944_ = \quotient[22]  & ~new_n12943_;
  assign new_n12945_ = ~new_n12355_ & ~new_n12765_;
  assign new_n12946_ = ~new_n12764_ & new_n12945_;
  assign new_n12947_ = ~new_n12944_ & ~new_n12946_;
  assign new_n12948_ = ~\b[23]  & ~new_n12947_;
  assign new_n12949_ = ~new_n12374_ & new_n12652_;
  assign new_n12950_ = ~new_n12648_ & new_n12949_;
  assign new_n12951_ = ~new_n12649_ & ~new_n12652_;
  assign new_n12952_ = ~new_n12950_ & ~new_n12951_;
  assign new_n12953_ = \quotient[22]  & ~new_n12952_;
  assign new_n12954_ = ~new_n12364_ & ~new_n12765_;
  assign new_n12955_ = ~new_n12764_ & new_n12954_;
  assign new_n12956_ = ~new_n12953_ & ~new_n12955_;
  assign new_n12957_ = ~\b[22]  & ~new_n12956_;
  assign new_n12958_ = ~new_n12383_ & new_n12647_;
  assign new_n12959_ = ~new_n12643_ & new_n12958_;
  assign new_n12960_ = ~new_n12644_ & ~new_n12647_;
  assign new_n12961_ = ~new_n12959_ & ~new_n12960_;
  assign new_n12962_ = \quotient[22]  & ~new_n12961_;
  assign new_n12963_ = ~new_n12373_ & ~new_n12765_;
  assign new_n12964_ = ~new_n12764_ & new_n12963_;
  assign new_n12965_ = ~new_n12962_ & ~new_n12964_;
  assign new_n12966_ = ~\b[21]  & ~new_n12965_;
  assign new_n12967_ = ~new_n12392_ & new_n12642_;
  assign new_n12968_ = ~new_n12638_ & new_n12967_;
  assign new_n12969_ = ~new_n12639_ & ~new_n12642_;
  assign new_n12970_ = ~new_n12968_ & ~new_n12969_;
  assign new_n12971_ = \quotient[22]  & ~new_n12970_;
  assign new_n12972_ = ~new_n12382_ & ~new_n12765_;
  assign new_n12973_ = ~new_n12764_ & new_n12972_;
  assign new_n12974_ = ~new_n12971_ & ~new_n12973_;
  assign new_n12975_ = ~\b[20]  & ~new_n12974_;
  assign new_n12976_ = ~new_n12401_ & new_n12637_;
  assign new_n12977_ = ~new_n12633_ & new_n12976_;
  assign new_n12978_ = ~new_n12634_ & ~new_n12637_;
  assign new_n12979_ = ~new_n12977_ & ~new_n12978_;
  assign new_n12980_ = \quotient[22]  & ~new_n12979_;
  assign new_n12981_ = ~new_n12391_ & ~new_n12765_;
  assign new_n12982_ = ~new_n12764_ & new_n12981_;
  assign new_n12983_ = ~new_n12980_ & ~new_n12982_;
  assign new_n12984_ = ~\b[19]  & ~new_n12983_;
  assign new_n12985_ = ~new_n12410_ & new_n12632_;
  assign new_n12986_ = ~new_n12628_ & new_n12985_;
  assign new_n12987_ = ~new_n12629_ & ~new_n12632_;
  assign new_n12988_ = ~new_n12986_ & ~new_n12987_;
  assign new_n12989_ = \quotient[22]  & ~new_n12988_;
  assign new_n12990_ = ~new_n12400_ & ~new_n12765_;
  assign new_n12991_ = ~new_n12764_ & new_n12990_;
  assign new_n12992_ = ~new_n12989_ & ~new_n12991_;
  assign new_n12993_ = ~\b[18]  & ~new_n12992_;
  assign new_n12994_ = ~new_n12419_ & new_n12627_;
  assign new_n12995_ = ~new_n12623_ & new_n12994_;
  assign new_n12996_ = ~new_n12624_ & ~new_n12627_;
  assign new_n12997_ = ~new_n12995_ & ~new_n12996_;
  assign new_n12998_ = \quotient[22]  & ~new_n12997_;
  assign new_n12999_ = ~new_n12409_ & ~new_n12765_;
  assign new_n13000_ = ~new_n12764_ & new_n12999_;
  assign new_n13001_ = ~new_n12998_ & ~new_n13000_;
  assign new_n13002_ = ~\b[17]  & ~new_n13001_;
  assign new_n13003_ = ~new_n12428_ & new_n12622_;
  assign new_n13004_ = ~new_n12618_ & new_n13003_;
  assign new_n13005_ = ~new_n12619_ & ~new_n12622_;
  assign new_n13006_ = ~new_n13004_ & ~new_n13005_;
  assign new_n13007_ = \quotient[22]  & ~new_n13006_;
  assign new_n13008_ = ~new_n12418_ & ~new_n12765_;
  assign new_n13009_ = ~new_n12764_ & new_n13008_;
  assign new_n13010_ = ~new_n13007_ & ~new_n13009_;
  assign new_n13011_ = ~\b[16]  & ~new_n13010_;
  assign new_n13012_ = ~new_n12437_ & new_n12617_;
  assign new_n13013_ = ~new_n12613_ & new_n13012_;
  assign new_n13014_ = ~new_n12614_ & ~new_n12617_;
  assign new_n13015_ = ~new_n13013_ & ~new_n13014_;
  assign new_n13016_ = \quotient[22]  & ~new_n13015_;
  assign new_n13017_ = ~new_n12427_ & ~new_n12765_;
  assign new_n13018_ = ~new_n12764_ & new_n13017_;
  assign new_n13019_ = ~new_n13016_ & ~new_n13018_;
  assign new_n13020_ = ~\b[15]  & ~new_n13019_;
  assign new_n13021_ = ~new_n12446_ & new_n12612_;
  assign new_n13022_ = ~new_n12608_ & new_n13021_;
  assign new_n13023_ = ~new_n12609_ & ~new_n12612_;
  assign new_n13024_ = ~new_n13022_ & ~new_n13023_;
  assign new_n13025_ = \quotient[22]  & ~new_n13024_;
  assign new_n13026_ = ~new_n12436_ & ~new_n12765_;
  assign new_n13027_ = ~new_n12764_ & new_n13026_;
  assign new_n13028_ = ~new_n13025_ & ~new_n13027_;
  assign new_n13029_ = ~\b[14]  & ~new_n13028_;
  assign new_n13030_ = ~new_n12455_ & new_n12607_;
  assign new_n13031_ = ~new_n12603_ & new_n13030_;
  assign new_n13032_ = ~new_n12604_ & ~new_n12607_;
  assign new_n13033_ = ~new_n13031_ & ~new_n13032_;
  assign new_n13034_ = \quotient[22]  & ~new_n13033_;
  assign new_n13035_ = ~new_n12445_ & ~new_n12765_;
  assign new_n13036_ = ~new_n12764_ & new_n13035_;
  assign new_n13037_ = ~new_n13034_ & ~new_n13036_;
  assign new_n13038_ = ~\b[13]  & ~new_n13037_;
  assign new_n13039_ = ~new_n12464_ & new_n12602_;
  assign new_n13040_ = ~new_n12598_ & new_n13039_;
  assign new_n13041_ = ~new_n12599_ & ~new_n12602_;
  assign new_n13042_ = ~new_n13040_ & ~new_n13041_;
  assign new_n13043_ = \quotient[22]  & ~new_n13042_;
  assign new_n13044_ = ~new_n12454_ & ~new_n12765_;
  assign new_n13045_ = ~new_n12764_ & new_n13044_;
  assign new_n13046_ = ~new_n13043_ & ~new_n13045_;
  assign new_n13047_ = ~\b[12]  & ~new_n13046_;
  assign new_n13048_ = ~new_n12473_ & new_n12597_;
  assign new_n13049_ = ~new_n12593_ & new_n13048_;
  assign new_n13050_ = ~new_n12594_ & ~new_n12597_;
  assign new_n13051_ = ~new_n13049_ & ~new_n13050_;
  assign new_n13052_ = \quotient[22]  & ~new_n13051_;
  assign new_n13053_ = ~new_n12463_ & ~new_n12765_;
  assign new_n13054_ = ~new_n12764_ & new_n13053_;
  assign new_n13055_ = ~new_n13052_ & ~new_n13054_;
  assign new_n13056_ = ~\b[11]  & ~new_n13055_;
  assign new_n13057_ = ~new_n12482_ & new_n12592_;
  assign new_n13058_ = ~new_n12588_ & new_n13057_;
  assign new_n13059_ = ~new_n12589_ & ~new_n12592_;
  assign new_n13060_ = ~new_n13058_ & ~new_n13059_;
  assign new_n13061_ = \quotient[22]  & ~new_n13060_;
  assign new_n13062_ = ~new_n12472_ & ~new_n12765_;
  assign new_n13063_ = ~new_n12764_ & new_n13062_;
  assign new_n13064_ = ~new_n13061_ & ~new_n13063_;
  assign new_n13065_ = ~\b[10]  & ~new_n13064_;
  assign new_n13066_ = ~new_n12491_ & new_n12587_;
  assign new_n13067_ = ~new_n12583_ & new_n13066_;
  assign new_n13068_ = ~new_n12584_ & ~new_n12587_;
  assign new_n13069_ = ~new_n13067_ & ~new_n13068_;
  assign new_n13070_ = \quotient[22]  & ~new_n13069_;
  assign new_n13071_ = ~new_n12481_ & ~new_n12765_;
  assign new_n13072_ = ~new_n12764_ & new_n13071_;
  assign new_n13073_ = ~new_n13070_ & ~new_n13072_;
  assign new_n13074_ = ~\b[9]  & ~new_n13073_;
  assign new_n13075_ = ~new_n12500_ & new_n12582_;
  assign new_n13076_ = ~new_n12578_ & new_n13075_;
  assign new_n13077_ = ~new_n12579_ & ~new_n12582_;
  assign new_n13078_ = ~new_n13076_ & ~new_n13077_;
  assign new_n13079_ = \quotient[22]  & ~new_n13078_;
  assign new_n13080_ = ~new_n12490_ & ~new_n12765_;
  assign new_n13081_ = ~new_n12764_ & new_n13080_;
  assign new_n13082_ = ~new_n13079_ & ~new_n13081_;
  assign new_n13083_ = ~\b[8]  & ~new_n13082_;
  assign new_n13084_ = ~new_n12509_ & new_n12577_;
  assign new_n13085_ = ~new_n12573_ & new_n13084_;
  assign new_n13086_ = ~new_n12574_ & ~new_n12577_;
  assign new_n13087_ = ~new_n13085_ & ~new_n13086_;
  assign new_n13088_ = \quotient[22]  & ~new_n13087_;
  assign new_n13089_ = ~new_n12499_ & ~new_n12765_;
  assign new_n13090_ = ~new_n12764_ & new_n13089_;
  assign new_n13091_ = ~new_n13088_ & ~new_n13090_;
  assign new_n13092_ = ~\b[7]  & ~new_n13091_;
  assign new_n13093_ = ~new_n12518_ & new_n12572_;
  assign new_n13094_ = ~new_n12568_ & new_n13093_;
  assign new_n13095_ = ~new_n12569_ & ~new_n12572_;
  assign new_n13096_ = ~new_n13094_ & ~new_n13095_;
  assign new_n13097_ = \quotient[22]  & ~new_n13096_;
  assign new_n13098_ = ~new_n12508_ & ~new_n12765_;
  assign new_n13099_ = ~new_n12764_ & new_n13098_;
  assign new_n13100_ = ~new_n13097_ & ~new_n13099_;
  assign new_n13101_ = ~\b[6]  & ~new_n13100_;
  assign new_n13102_ = ~new_n12527_ & new_n12567_;
  assign new_n13103_ = ~new_n12563_ & new_n13102_;
  assign new_n13104_ = ~new_n12564_ & ~new_n12567_;
  assign new_n13105_ = ~new_n13103_ & ~new_n13104_;
  assign new_n13106_ = \quotient[22]  & ~new_n13105_;
  assign new_n13107_ = ~new_n12517_ & ~new_n12765_;
  assign new_n13108_ = ~new_n12764_ & new_n13107_;
  assign new_n13109_ = ~new_n13106_ & ~new_n13108_;
  assign new_n13110_ = ~\b[5]  & ~new_n13109_;
  assign new_n13111_ = ~new_n12535_ & new_n12562_;
  assign new_n13112_ = ~new_n12558_ & new_n13111_;
  assign new_n13113_ = ~new_n12559_ & ~new_n12562_;
  assign new_n13114_ = ~new_n13112_ & ~new_n13113_;
  assign new_n13115_ = \quotient[22]  & ~new_n13114_;
  assign new_n13116_ = ~new_n12526_ & ~new_n12765_;
  assign new_n13117_ = ~new_n12764_ & new_n13116_;
  assign new_n13118_ = ~new_n13115_ & ~new_n13117_;
  assign new_n13119_ = ~\b[4]  & ~new_n13118_;
  assign new_n13120_ = ~new_n12553_ & new_n12557_;
  assign new_n13121_ = ~new_n12552_ & new_n13120_;
  assign new_n13122_ = ~new_n12554_ & ~new_n12557_;
  assign new_n13123_ = ~new_n13121_ & ~new_n13122_;
  assign new_n13124_ = \quotient[22]  & ~new_n13123_;
  assign new_n13125_ = ~new_n12534_ & ~new_n12765_;
  assign new_n13126_ = ~new_n12764_ & new_n13125_;
  assign new_n13127_ = ~new_n13124_ & ~new_n13126_;
  assign new_n13128_ = ~\b[3]  & ~new_n13127_;
  assign new_n13129_ = ~new_n12549_ & new_n12551_;
  assign new_n13130_ = ~new_n12547_ & new_n13129_;
  assign new_n13131_ = ~new_n12552_ & ~new_n13130_;
  assign new_n13132_ = \quotient[22]  & new_n13131_;
  assign new_n13133_ = ~new_n12546_ & ~new_n12765_;
  assign new_n13134_ = ~new_n12764_ & new_n13133_;
  assign new_n13135_ = ~new_n13132_ & ~new_n13134_;
  assign new_n13136_ = ~\b[2]  & ~new_n13135_;
  assign new_n13137_ = \b[0]  & \quotient[22] ;
  assign new_n13138_ = \a[22]  & ~new_n13137_;
  assign new_n13139_ = new_n12551_ & \quotient[22] ;
  assign new_n13140_ = ~new_n13138_ & ~new_n13139_;
  assign new_n13141_ = \b[1]  & ~new_n13140_;
  assign new_n13142_ = ~\b[1]  & ~new_n13139_;
  assign new_n13143_ = ~new_n13138_ & new_n13142_;
  assign new_n13144_ = ~new_n13141_ & ~new_n13143_;
  assign new_n13145_ = ~\a[21]  & \b[0] ;
  assign new_n13146_ = ~new_n13144_ & ~new_n13145_;
  assign new_n13147_ = ~\b[1]  & ~new_n13140_;
  assign new_n13148_ = ~new_n13146_ & ~new_n13147_;
  assign new_n13149_ = \b[2]  & ~new_n13134_;
  assign new_n13150_ = ~new_n13132_ & new_n13149_;
  assign new_n13151_ = ~new_n13136_ & ~new_n13150_;
  assign new_n13152_ = ~new_n13148_ & new_n13151_;
  assign new_n13153_ = ~new_n13136_ & ~new_n13152_;
  assign new_n13154_ = \b[3]  & ~new_n13126_;
  assign new_n13155_ = ~new_n13124_ & new_n13154_;
  assign new_n13156_ = ~new_n13128_ & ~new_n13155_;
  assign new_n13157_ = ~new_n13153_ & new_n13156_;
  assign new_n13158_ = ~new_n13128_ & ~new_n13157_;
  assign new_n13159_ = \b[4]  & ~new_n13117_;
  assign new_n13160_ = ~new_n13115_ & new_n13159_;
  assign new_n13161_ = ~new_n13119_ & ~new_n13160_;
  assign new_n13162_ = ~new_n13158_ & new_n13161_;
  assign new_n13163_ = ~new_n13119_ & ~new_n13162_;
  assign new_n13164_ = \b[5]  & ~new_n13108_;
  assign new_n13165_ = ~new_n13106_ & new_n13164_;
  assign new_n13166_ = ~new_n13110_ & ~new_n13165_;
  assign new_n13167_ = ~new_n13163_ & new_n13166_;
  assign new_n13168_ = ~new_n13110_ & ~new_n13167_;
  assign new_n13169_ = \b[6]  & ~new_n13099_;
  assign new_n13170_ = ~new_n13097_ & new_n13169_;
  assign new_n13171_ = ~new_n13101_ & ~new_n13170_;
  assign new_n13172_ = ~new_n13168_ & new_n13171_;
  assign new_n13173_ = ~new_n13101_ & ~new_n13172_;
  assign new_n13174_ = \b[7]  & ~new_n13090_;
  assign new_n13175_ = ~new_n13088_ & new_n13174_;
  assign new_n13176_ = ~new_n13092_ & ~new_n13175_;
  assign new_n13177_ = ~new_n13173_ & new_n13176_;
  assign new_n13178_ = ~new_n13092_ & ~new_n13177_;
  assign new_n13179_ = \b[8]  & ~new_n13081_;
  assign new_n13180_ = ~new_n13079_ & new_n13179_;
  assign new_n13181_ = ~new_n13083_ & ~new_n13180_;
  assign new_n13182_ = ~new_n13178_ & new_n13181_;
  assign new_n13183_ = ~new_n13083_ & ~new_n13182_;
  assign new_n13184_ = \b[9]  & ~new_n13072_;
  assign new_n13185_ = ~new_n13070_ & new_n13184_;
  assign new_n13186_ = ~new_n13074_ & ~new_n13185_;
  assign new_n13187_ = ~new_n13183_ & new_n13186_;
  assign new_n13188_ = ~new_n13074_ & ~new_n13187_;
  assign new_n13189_ = \b[10]  & ~new_n13063_;
  assign new_n13190_ = ~new_n13061_ & new_n13189_;
  assign new_n13191_ = ~new_n13065_ & ~new_n13190_;
  assign new_n13192_ = ~new_n13188_ & new_n13191_;
  assign new_n13193_ = ~new_n13065_ & ~new_n13192_;
  assign new_n13194_ = \b[11]  & ~new_n13054_;
  assign new_n13195_ = ~new_n13052_ & new_n13194_;
  assign new_n13196_ = ~new_n13056_ & ~new_n13195_;
  assign new_n13197_ = ~new_n13193_ & new_n13196_;
  assign new_n13198_ = ~new_n13056_ & ~new_n13197_;
  assign new_n13199_ = \b[12]  & ~new_n13045_;
  assign new_n13200_ = ~new_n13043_ & new_n13199_;
  assign new_n13201_ = ~new_n13047_ & ~new_n13200_;
  assign new_n13202_ = ~new_n13198_ & new_n13201_;
  assign new_n13203_ = ~new_n13047_ & ~new_n13202_;
  assign new_n13204_ = \b[13]  & ~new_n13036_;
  assign new_n13205_ = ~new_n13034_ & new_n13204_;
  assign new_n13206_ = ~new_n13038_ & ~new_n13205_;
  assign new_n13207_ = ~new_n13203_ & new_n13206_;
  assign new_n13208_ = ~new_n13038_ & ~new_n13207_;
  assign new_n13209_ = \b[14]  & ~new_n13027_;
  assign new_n13210_ = ~new_n13025_ & new_n13209_;
  assign new_n13211_ = ~new_n13029_ & ~new_n13210_;
  assign new_n13212_ = ~new_n13208_ & new_n13211_;
  assign new_n13213_ = ~new_n13029_ & ~new_n13212_;
  assign new_n13214_ = \b[15]  & ~new_n13018_;
  assign new_n13215_ = ~new_n13016_ & new_n13214_;
  assign new_n13216_ = ~new_n13020_ & ~new_n13215_;
  assign new_n13217_ = ~new_n13213_ & new_n13216_;
  assign new_n13218_ = ~new_n13020_ & ~new_n13217_;
  assign new_n13219_ = \b[16]  & ~new_n13009_;
  assign new_n13220_ = ~new_n13007_ & new_n13219_;
  assign new_n13221_ = ~new_n13011_ & ~new_n13220_;
  assign new_n13222_ = ~new_n13218_ & new_n13221_;
  assign new_n13223_ = ~new_n13011_ & ~new_n13222_;
  assign new_n13224_ = \b[17]  & ~new_n13000_;
  assign new_n13225_ = ~new_n12998_ & new_n13224_;
  assign new_n13226_ = ~new_n13002_ & ~new_n13225_;
  assign new_n13227_ = ~new_n13223_ & new_n13226_;
  assign new_n13228_ = ~new_n13002_ & ~new_n13227_;
  assign new_n13229_ = \b[18]  & ~new_n12991_;
  assign new_n13230_ = ~new_n12989_ & new_n13229_;
  assign new_n13231_ = ~new_n12993_ & ~new_n13230_;
  assign new_n13232_ = ~new_n13228_ & new_n13231_;
  assign new_n13233_ = ~new_n12993_ & ~new_n13232_;
  assign new_n13234_ = \b[19]  & ~new_n12982_;
  assign new_n13235_ = ~new_n12980_ & new_n13234_;
  assign new_n13236_ = ~new_n12984_ & ~new_n13235_;
  assign new_n13237_ = ~new_n13233_ & new_n13236_;
  assign new_n13238_ = ~new_n12984_ & ~new_n13237_;
  assign new_n13239_ = \b[20]  & ~new_n12973_;
  assign new_n13240_ = ~new_n12971_ & new_n13239_;
  assign new_n13241_ = ~new_n12975_ & ~new_n13240_;
  assign new_n13242_ = ~new_n13238_ & new_n13241_;
  assign new_n13243_ = ~new_n12975_ & ~new_n13242_;
  assign new_n13244_ = \b[21]  & ~new_n12964_;
  assign new_n13245_ = ~new_n12962_ & new_n13244_;
  assign new_n13246_ = ~new_n12966_ & ~new_n13245_;
  assign new_n13247_ = ~new_n13243_ & new_n13246_;
  assign new_n13248_ = ~new_n12966_ & ~new_n13247_;
  assign new_n13249_ = \b[22]  & ~new_n12955_;
  assign new_n13250_ = ~new_n12953_ & new_n13249_;
  assign new_n13251_ = ~new_n12957_ & ~new_n13250_;
  assign new_n13252_ = ~new_n13248_ & new_n13251_;
  assign new_n13253_ = ~new_n12957_ & ~new_n13252_;
  assign new_n13254_ = \b[23]  & ~new_n12946_;
  assign new_n13255_ = ~new_n12944_ & new_n13254_;
  assign new_n13256_ = ~new_n12948_ & ~new_n13255_;
  assign new_n13257_ = ~new_n13253_ & new_n13256_;
  assign new_n13258_ = ~new_n12948_ & ~new_n13257_;
  assign new_n13259_ = \b[24]  & ~new_n12937_;
  assign new_n13260_ = ~new_n12935_ & new_n13259_;
  assign new_n13261_ = ~new_n12939_ & ~new_n13260_;
  assign new_n13262_ = ~new_n13258_ & new_n13261_;
  assign new_n13263_ = ~new_n12939_ & ~new_n13262_;
  assign new_n13264_ = \b[25]  & ~new_n12928_;
  assign new_n13265_ = ~new_n12926_ & new_n13264_;
  assign new_n13266_ = ~new_n12930_ & ~new_n13265_;
  assign new_n13267_ = ~new_n13263_ & new_n13266_;
  assign new_n13268_ = ~new_n12930_ & ~new_n13267_;
  assign new_n13269_ = \b[26]  & ~new_n12919_;
  assign new_n13270_ = ~new_n12917_ & new_n13269_;
  assign new_n13271_ = ~new_n12921_ & ~new_n13270_;
  assign new_n13272_ = ~new_n13268_ & new_n13271_;
  assign new_n13273_ = ~new_n12921_ & ~new_n13272_;
  assign new_n13274_ = \b[27]  & ~new_n12910_;
  assign new_n13275_ = ~new_n12908_ & new_n13274_;
  assign new_n13276_ = ~new_n12912_ & ~new_n13275_;
  assign new_n13277_ = ~new_n13273_ & new_n13276_;
  assign new_n13278_ = ~new_n12912_ & ~new_n13277_;
  assign new_n13279_ = \b[28]  & ~new_n12901_;
  assign new_n13280_ = ~new_n12899_ & new_n13279_;
  assign new_n13281_ = ~new_n12903_ & ~new_n13280_;
  assign new_n13282_ = ~new_n13278_ & new_n13281_;
  assign new_n13283_ = ~new_n12903_ & ~new_n13282_;
  assign new_n13284_ = \b[29]  & ~new_n12892_;
  assign new_n13285_ = ~new_n12890_ & new_n13284_;
  assign new_n13286_ = ~new_n12894_ & ~new_n13285_;
  assign new_n13287_ = ~new_n13283_ & new_n13286_;
  assign new_n13288_ = ~new_n12894_ & ~new_n13287_;
  assign new_n13289_ = \b[30]  & ~new_n12883_;
  assign new_n13290_ = ~new_n12881_ & new_n13289_;
  assign new_n13291_ = ~new_n12885_ & ~new_n13290_;
  assign new_n13292_ = ~new_n13288_ & new_n13291_;
  assign new_n13293_ = ~new_n12885_ & ~new_n13292_;
  assign new_n13294_ = \b[31]  & ~new_n12874_;
  assign new_n13295_ = ~new_n12872_ & new_n13294_;
  assign new_n13296_ = ~new_n12876_ & ~new_n13295_;
  assign new_n13297_ = ~new_n13293_ & new_n13296_;
  assign new_n13298_ = ~new_n12876_ & ~new_n13297_;
  assign new_n13299_ = \b[32]  & ~new_n12865_;
  assign new_n13300_ = ~new_n12863_ & new_n13299_;
  assign new_n13301_ = ~new_n12867_ & ~new_n13300_;
  assign new_n13302_ = ~new_n13298_ & new_n13301_;
  assign new_n13303_ = ~new_n12867_ & ~new_n13302_;
  assign new_n13304_ = \b[33]  & ~new_n12856_;
  assign new_n13305_ = ~new_n12854_ & new_n13304_;
  assign new_n13306_ = ~new_n12858_ & ~new_n13305_;
  assign new_n13307_ = ~new_n13303_ & new_n13306_;
  assign new_n13308_ = ~new_n12858_ & ~new_n13307_;
  assign new_n13309_ = \b[34]  & ~new_n12847_;
  assign new_n13310_ = ~new_n12845_ & new_n13309_;
  assign new_n13311_ = ~new_n12849_ & ~new_n13310_;
  assign new_n13312_ = ~new_n13308_ & new_n13311_;
  assign new_n13313_ = ~new_n12849_ & ~new_n13312_;
  assign new_n13314_ = \b[35]  & ~new_n12838_;
  assign new_n13315_ = ~new_n12836_ & new_n13314_;
  assign new_n13316_ = ~new_n12840_ & ~new_n13315_;
  assign new_n13317_ = ~new_n13313_ & new_n13316_;
  assign new_n13318_ = ~new_n12840_ & ~new_n13317_;
  assign new_n13319_ = \b[36]  & ~new_n12829_;
  assign new_n13320_ = ~new_n12827_ & new_n13319_;
  assign new_n13321_ = ~new_n12831_ & ~new_n13320_;
  assign new_n13322_ = ~new_n13318_ & new_n13321_;
  assign new_n13323_ = ~new_n12831_ & ~new_n13322_;
  assign new_n13324_ = \b[37]  & ~new_n12820_;
  assign new_n13325_ = ~new_n12818_ & new_n13324_;
  assign new_n13326_ = ~new_n12822_ & ~new_n13325_;
  assign new_n13327_ = ~new_n13323_ & new_n13326_;
  assign new_n13328_ = ~new_n12822_ & ~new_n13327_;
  assign new_n13329_ = \b[38]  & ~new_n12811_;
  assign new_n13330_ = ~new_n12809_ & new_n13329_;
  assign new_n13331_ = ~new_n12813_ & ~new_n13330_;
  assign new_n13332_ = ~new_n13328_ & new_n13331_;
  assign new_n13333_ = ~new_n12813_ & ~new_n13332_;
  assign new_n13334_ = \b[39]  & ~new_n12802_;
  assign new_n13335_ = ~new_n12800_ & new_n13334_;
  assign new_n13336_ = ~new_n12804_ & ~new_n13335_;
  assign new_n13337_ = ~new_n13333_ & new_n13336_;
  assign new_n13338_ = ~new_n12804_ & ~new_n13337_;
  assign new_n13339_ = \b[40]  & ~new_n12793_;
  assign new_n13340_ = ~new_n12791_ & new_n13339_;
  assign new_n13341_ = ~new_n12795_ & ~new_n13340_;
  assign new_n13342_ = ~new_n13338_ & new_n13341_;
  assign new_n13343_ = ~new_n12795_ & ~new_n13342_;
  assign new_n13344_ = \b[41]  & ~new_n12773_;
  assign new_n13345_ = ~new_n12771_ & new_n13344_;
  assign new_n13346_ = ~new_n12786_ & ~new_n13345_;
  assign new_n13347_ = ~new_n13343_ & new_n13346_;
  assign new_n13348_ = ~new_n12786_ & ~new_n13347_;
  assign new_n13349_ = \b[42]  & ~new_n12783_;
  assign new_n13350_ = ~new_n12781_ & new_n13349_;
  assign new_n13351_ = ~new_n12785_ & ~new_n13350_;
  assign new_n13352_ = ~new_n13348_ & new_n13351_;
  assign new_n13353_ = ~new_n12785_ & ~new_n13352_;
  assign new_n13354_ = new_n418_ & new_n420_;
  assign new_n13355_ = new_n408_ & new_n13354_;
  assign \quotient[21]  = ~new_n13353_ & new_n13355_;
  assign new_n13357_ = ~new_n12774_ & ~\quotient[21] ;
  assign new_n13358_ = ~new_n12795_ & new_n13346_;
  assign new_n13359_ = ~new_n13342_ & new_n13358_;
  assign new_n13360_ = ~new_n13343_ & ~new_n13346_;
  assign new_n13361_ = ~new_n13359_ & ~new_n13360_;
  assign new_n13362_ = new_n13355_ & ~new_n13361_;
  assign new_n13363_ = ~new_n13353_ & new_n13362_;
  assign new_n13364_ = ~new_n13357_ & ~new_n13363_;
  assign new_n13365_ = ~\b[42]  & ~new_n13364_;
  assign new_n13366_ = ~new_n12794_ & ~\quotient[21] ;
  assign new_n13367_ = ~new_n12804_ & new_n13341_;
  assign new_n13368_ = ~new_n13337_ & new_n13367_;
  assign new_n13369_ = ~new_n13338_ & ~new_n13341_;
  assign new_n13370_ = ~new_n13368_ & ~new_n13369_;
  assign new_n13371_ = new_n13355_ & ~new_n13370_;
  assign new_n13372_ = ~new_n13353_ & new_n13371_;
  assign new_n13373_ = ~new_n13366_ & ~new_n13372_;
  assign new_n13374_ = ~\b[41]  & ~new_n13373_;
  assign new_n13375_ = ~new_n12803_ & ~\quotient[21] ;
  assign new_n13376_ = ~new_n12813_ & new_n13336_;
  assign new_n13377_ = ~new_n13332_ & new_n13376_;
  assign new_n13378_ = ~new_n13333_ & ~new_n13336_;
  assign new_n13379_ = ~new_n13377_ & ~new_n13378_;
  assign new_n13380_ = new_n13355_ & ~new_n13379_;
  assign new_n13381_ = ~new_n13353_ & new_n13380_;
  assign new_n13382_ = ~new_n13375_ & ~new_n13381_;
  assign new_n13383_ = ~\b[40]  & ~new_n13382_;
  assign new_n13384_ = ~new_n12812_ & ~\quotient[21] ;
  assign new_n13385_ = ~new_n12822_ & new_n13331_;
  assign new_n13386_ = ~new_n13327_ & new_n13385_;
  assign new_n13387_ = ~new_n13328_ & ~new_n13331_;
  assign new_n13388_ = ~new_n13386_ & ~new_n13387_;
  assign new_n13389_ = new_n13355_ & ~new_n13388_;
  assign new_n13390_ = ~new_n13353_ & new_n13389_;
  assign new_n13391_ = ~new_n13384_ & ~new_n13390_;
  assign new_n13392_ = ~\b[39]  & ~new_n13391_;
  assign new_n13393_ = ~new_n12821_ & ~\quotient[21] ;
  assign new_n13394_ = ~new_n12831_ & new_n13326_;
  assign new_n13395_ = ~new_n13322_ & new_n13394_;
  assign new_n13396_ = ~new_n13323_ & ~new_n13326_;
  assign new_n13397_ = ~new_n13395_ & ~new_n13396_;
  assign new_n13398_ = new_n13355_ & ~new_n13397_;
  assign new_n13399_ = ~new_n13353_ & new_n13398_;
  assign new_n13400_ = ~new_n13393_ & ~new_n13399_;
  assign new_n13401_ = ~\b[38]  & ~new_n13400_;
  assign new_n13402_ = ~new_n12830_ & ~\quotient[21] ;
  assign new_n13403_ = ~new_n12840_ & new_n13321_;
  assign new_n13404_ = ~new_n13317_ & new_n13403_;
  assign new_n13405_ = ~new_n13318_ & ~new_n13321_;
  assign new_n13406_ = ~new_n13404_ & ~new_n13405_;
  assign new_n13407_ = new_n13355_ & ~new_n13406_;
  assign new_n13408_ = ~new_n13353_ & new_n13407_;
  assign new_n13409_ = ~new_n13402_ & ~new_n13408_;
  assign new_n13410_ = ~\b[37]  & ~new_n13409_;
  assign new_n13411_ = ~new_n12839_ & ~\quotient[21] ;
  assign new_n13412_ = ~new_n12849_ & new_n13316_;
  assign new_n13413_ = ~new_n13312_ & new_n13412_;
  assign new_n13414_ = ~new_n13313_ & ~new_n13316_;
  assign new_n13415_ = ~new_n13413_ & ~new_n13414_;
  assign new_n13416_ = new_n13355_ & ~new_n13415_;
  assign new_n13417_ = ~new_n13353_ & new_n13416_;
  assign new_n13418_ = ~new_n13411_ & ~new_n13417_;
  assign new_n13419_ = ~\b[36]  & ~new_n13418_;
  assign new_n13420_ = ~new_n12848_ & ~\quotient[21] ;
  assign new_n13421_ = ~new_n12858_ & new_n13311_;
  assign new_n13422_ = ~new_n13307_ & new_n13421_;
  assign new_n13423_ = ~new_n13308_ & ~new_n13311_;
  assign new_n13424_ = ~new_n13422_ & ~new_n13423_;
  assign new_n13425_ = new_n13355_ & ~new_n13424_;
  assign new_n13426_ = ~new_n13353_ & new_n13425_;
  assign new_n13427_ = ~new_n13420_ & ~new_n13426_;
  assign new_n13428_ = ~\b[35]  & ~new_n13427_;
  assign new_n13429_ = ~new_n12857_ & ~\quotient[21] ;
  assign new_n13430_ = ~new_n12867_ & new_n13306_;
  assign new_n13431_ = ~new_n13302_ & new_n13430_;
  assign new_n13432_ = ~new_n13303_ & ~new_n13306_;
  assign new_n13433_ = ~new_n13431_ & ~new_n13432_;
  assign new_n13434_ = new_n13355_ & ~new_n13433_;
  assign new_n13435_ = ~new_n13353_ & new_n13434_;
  assign new_n13436_ = ~new_n13429_ & ~new_n13435_;
  assign new_n13437_ = ~\b[34]  & ~new_n13436_;
  assign new_n13438_ = ~new_n12866_ & ~\quotient[21] ;
  assign new_n13439_ = ~new_n12876_ & new_n13301_;
  assign new_n13440_ = ~new_n13297_ & new_n13439_;
  assign new_n13441_ = ~new_n13298_ & ~new_n13301_;
  assign new_n13442_ = ~new_n13440_ & ~new_n13441_;
  assign new_n13443_ = new_n13355_ & ~new_n13442_;
  assign new_n13444_ = ~new_n13353_ & new_n13443_;
  assign new_n13445_ = ~new_n13438_ & ~new_n13444_;
  assign new_n13446_ = ~\b[33]  & ~new_n13445_;
  assign new_n13447_ = ~new_n12875_ & ~\quotient[21] ;
  assign new_n13448_ = ~new_n12885_ & new_n13296_;
  assign new_n13449_ = ~new_n13292_ & new_n13448_;
  assign new_n13450_ = ~new_n13293_ & ~new_n13296_;
  assign new_n13451_ = ~new_n13449_ & ~new_n13450_;
  assign new_n13452_ = new_n13355_ & ~new_n13451_;
  assign new_n13453_ = ~new_n13353_ & new_n13452_;
  assign new_n13454_ = ~new_n13447_ & ~new_n13453_;
  assign new_n13455_ = ~\b[32]  & ~new_n13454_;
  assign new_n13456_ = ~new_n12884_ & ~\quotient[21] ;
  assign new_n13457_ = ~new_n12894_ & new_n13291_;
  assign new_n13458_ = ~new_n13287_ & new_n13457_;
  assign new_n13459_ = ~new_n13288_ & ~new_n13291_;
  assign new_n13460_ = ~new_n13458_ & ~new_n13459_;
  assign new_n13461_ = new_n13355_ & ~new_n13460_;
  assign new_n13462_ = ~new_n13353_ & new_n13461_;
  assign new_n13463_ = ~new_n13456_ & ~new_n13462_;
  assign new_n13464_ = ~\b[31]  & ~new_n13463_;
  assign new_n13465_ = ~new_n12893_ & ~\quotient[21] ;
  assign new_n13466_ = ~new_n12903_ & new_n13286_;
  assign new_n13467_ = ~new_n13282_ & new_n13466_;
  assign new_n13468_ = ~new_n13283_ & ~new_n13286_;
  assign new_n13469_ = ~new_n13467_ & ~new_n13468_;
  assign new_n13470_ = new_n13355_ & ~new_n13469_;
  assign new_n13471_ = ~new_n13353_ & new_n13470_;
  assign new_n13472_ = ~new_n13465_ & ~new_n13471_;
  assign new_n13473_ = ~\b[30]  & ~new_n13472_;
  assign new_n13474_ = ~new_n12902_ & ~\quotient[21] ;
  assign new_n13475_ = ~new_n12912_ & new_n13281_;
  assign new_n13476_ = ~new_n13277_ & new_n13475_;
  assign new_n13477_ = ~new_n13278_ & ~new_n13281_;
  assign new_n13478_ = ~new_n13476_ & ~new_n13477_;
  assign new_n13479_ = new_n13355_ & ~new_n13478_;
  assign new_n13480_ = ~new_n13353_ & new_n13479_;
  assign new_n13481_ = ~new_n13474_ & ~new_n13480_;
  assign new_n13482_ = ~\b[29]  & ~new_n13481_;
  assign new_n13483_ = ~new_n12911_ & ~\quotient[21] ;
  assign new_n13484_ = ~new_n12921_ & new_n13276_;
  assign new_n13485_ = ~new_n13272_ & new_n13484_;
  assign new_n13486_ = ~new_n13273_ & ~new_n13276_;
  assign new_n13487_ = ~new_n13485_ & ~new_n13486_;
  assign new_n13488_ = new_n13355_ & ~new_n13487_;
  assign new_n13489_ = ~new_n13353_ & new_n13488_;
  assign new_n13490_ = ~new_n13483_ & ~new_n13489_;
  assign new_n13491_ = ~\b[28]  & ~new_n13490_;
  assign new_n13492_ = ~new_n12920_ & ~\quotient[21] ;
  assign new_n13493_ = ~new_n12930_ & new_n13271_;
  assign new_n13494_ = ~new_n13267_ & new_n13493_;
  assign new_n13495_ = ~new_n13268_ & ~new_n13271_;
  assign new_n13496_ = ~new_n13494_ & ~new_n13495_;
  assign new_n13497_ = new_n13355_ & ~new_n13496_;
  assign new_n13498_ = ~new_n13353_ & new_n13497_;
  assign new_n13499_ = ~new_n13492_ & ~new_n13498_;
  assign new_n13500_ = ~\b[27]  & ~new_n13499_;
  assign new_n13501_ = ~new_n12929_ & ~\quotient[21] ;
  assign new_n13502_ = ~new_n12939_ & new_n13266_;
  assign new_n13503_ = ~new_n13262_ & new_n13502_;
  assign new_n13504_ = ~new_n13263_ & ~new_n13266_;
  assign new_n13505_ = ~new_n13503_ & ~new_n13504_;
  assign new_n13506_ = new_n13355_ & ~new_n13505_;
  assign new_n13507_ = ~new_n13353_ & new_n13506_;
  assign new_n13508_ = ~new_n13501_ & ~new_n13507_;
  assign new_n13509_ = ~\b[26]  & ~new_n13508_;
  assign new_n13510_ = ~new_n12938_ & ~\quotient[21] ;
  assign new_n13511_ = ~new_n12948_ & new_n13261_;
  assign new_n13512_ = ~new_n13257_ & new_n13511_;
  assign new_n13513_ = ~new_n13258_ & ~new_n13261_;
  assign new_n13514_ = ~new_n13512_ & ~new_n13513_;
  assign new_n13515_ = new_n13355_ & ~new_n13514_;
  assign new_n13516_ = ~new_n13353_ & new_n13515_;
  assign new_n13517_ = ~new_n13510_ & ~new_n13516_;
  assign new_n13518_ = ~\b[25]  & ~new_n13517_;
  assign new_n13519_ = ~new_n12947_ & ~\quotient[21] ;
  assign new_n13520_ = ~new_n12957_ & new_n13256_;
  assign new_n13521_ = ~new_n13252_ & new_n13520_;
  assign new_n13522_ = ~new_n13253_ & ~new_n13256_;
  assign new_n13523_ = ~new_n13521_ & ~new_n13522_;
  assign new_n13524_ = new_n13355_ & ~new_n13523_;
  assign new_n13525_ = ~new_n13353_ & new_n13524_;
  assign new_n13526_ = ~new_n13519_ & ~new_n13525_;
  assign new_n13527_ = ~\b[24]  & ~new_n13526_;
  assign new_n13528_ = ~new_n12956_ & ~\quotient[21] ;
  assign new_n13529_ = ~new_n12966_ & new_n13251_;
  assign new_n13530_ = ~new_n13247_ & new_n13529_;
  assign new_n13531_ = ~new_n13248_ & ~new_n13251_;
  assign new_n13532_ = ~new_n13530_ & ~new_n13531_;
  assign new_n13533_ = new_n13355_ & ~new_n13532_;
  assign new_n13534_ = ~new_n13353_ & new_n13533_;
  assign new_n13535_ = ~new_n13528_ & ~new_n13534_;
  assign new_n13536_ = ~\b[23]  & ~new_n13535_;
  assign new_n13537_ = ~new_n12965_ & ~\quotient[21] ;
  assign new_n13538_ = ~new_n12975_ & new_n13246_;
  assign new_n13539_ = ~new_n13242_ & new_n13538_;
  assign new_n13540_ = ~new_n13243_ & ~new_n13246_;
  assign new_n13541_ = ~new_n13539_ & ~new_n13540_;
  assign new_n13542_ = new_n13355_ & ~new_n13541_;
  assign new_n13543_ = ~new_n13353_ & new_n13542_;
  assign new_n13544_ = ~new_n13537_ & ~new_n13543_;
  assign new_n13545_ = ~\b[22]  & ~new_n13544_;
  assign new_n13546_ = ~new_n12974_ & ~\quotient[21] ;
  assign new_n13547_ = ~new_n12984_ & new_n13241_;
  assign new_n13548_ = ~new_n13237_ & new_n13547_;
  assign new_n13549_ = ~new_n13238_ & ~new_n13241_;
  assign new_n13550_ = ~new_n13548_ & ~new_n13549_;
  assign new_n13551_ = new_n13355_ & ~new_n13550_;
  assign new_n13552_ = ~new_n13353_ & new_n13551_;
  assign new_n13553_ = ~new_n13546_ & ~new_n13552_;
  assign new_n13554_ = ~\b[21]  & ~new_n13553_;
  assign new_n13555_ = ~new_n12983_ & ~\quotient[21] ;
  assign new_n13556_ = ~new_n12993_ & new_n13236_;
  assign new_n13557_ = ~new_n13232_ & new_n13556_;
  assign new_n13558_ = ~new_n13233_ & ~new_n13236_;
  assign new_n13559_ = ~new_n13557_ & ~new_n13558_;
  assign new_n13560_ = new_n13355_ & ~new_n13559_;
  assign new_n13561_ = ~new_n13353_ & new_n13560_;
  assign new_n13562_ = ~new_n13555_ & ~new_n13561_;
  assign new_n13563_ = ~\b[20]  & ~new_n13562_;
  assign new_n13564_ = ~new_n12992_ & ~\quotient[21] ;
  assign new_n13565_ = ~new_n13002_ & new_n13231_;
  assign new_n13566_ = ~new_n13227_ & new_n13565_;
  assign new_n13567_ = ~new_n13228_ & ~new_n13231_;
  assign new_n13568_ = ~new_n13566_ & ~new_n13567_;
  assign new_n13569_ = new_n13355_ & ~new_n13568_;
  assign new_n13570_ = ~new_n13353_ & new_n13569_;
  assign new_n13571_ = ~new_n13564_ & ~new_n13570_;
  assign new_n13572_ = ~\b[19]  & ~new_n13571_;
  assign new_n13573_ = ~new_n13001_ & ~\quotient[21] ;
  assign new_n13574_ = ~new_n13011_ & new_n13226_;
  assign new_n13575_ = ~new_n13222_ & new_n13574_;
  assign new_n13576_ = ~new_n13223_ & ~new_n13226_;
  assign new_n13577_ = ~new_n13575_ & ~new_n13576_;
  assign new_n13578_ = new_n13355_ & ~new_n13577_;
  assign new_n13579_ = ~new_n13353_ & new_n13578_;
  assign new_n13580_ = ~new_n13573_ & ~new_n13579_;
  assign new_n13581_ = ~\b[18]  & ~new_n13580_;
  assign new_n13582_ = ~new_n13010_ & ~\quotient[21] ;
  assign new_n13583_ = ~new_n13020_ & new_n13221_;
  assign new_n13584_ = ~new_n13217_ & new_n13583_;
  assign new_n13585_ = ~new_n13218_ & ~new_n13221_;
  assign new_n13586_ = ~new_n13584_ & ~new_n13585_;
  assign new_n13587_ = new_n13355_ & ~new_n13586_;
  assign new_n13588_ = ~new_n13353_ & new_n13587_;
  assign new_n13589_ = ~new_n13582_ & ~new_n13588_;
  assign new_n13590_ = ~\b[17]  & ~new_n13589_;
  assign new_n13591_ = ~new_n13019_ & ~\quotient[21] ;
  assign new_n13592_ = ~new_n13029_ & new_n13216_;
  assign new_n13593_ = ~new_n13212_ & new_n13592_;
  assign new_n13594_ = ~new_n13213_ & ~new_n13216_;
  assign new_n13595_ = ~new_n13593_ & ~new_n13594_;
  assign new_n13596_ = new_n13355_ & ~new_n13595_;
  assign new_n13597_ = ~new_n13353_ & new_n13596_;
  assign new_n13598_ = ~new_n13591_ & ~new_n13597_;
  assign new_n13599_ = ~\b[16]  & ~new_n13598_;
  assign new_n13600_ = ~new_n13028_ & ~\quotient[21] ;
  assign new_n13601_ = ~new_n13038_ & new_n13211_;
  assign new_n13602_ = ~new_n13207_ & new_n13601_;
  assign new_n13603_ = ~new_n13208_ & ~new_n13211_;
  assign new_n13604_ = ~new_n13602_ & ~new_n13603_;
  assign new_n13605_ = new_n13355_ & ~new_n13604_;
  assign new_n13606_ = ~new_n13353_ & new_n13605_;
  assign new_n13607_ = ~new_n13600_ & ~new_n13606_;
  assign new_n13608_ = ~\b[15]  & ~new_n13607_;
  assign new_n13609_ = ~new_n13037_ & ~\quotient[21] ;
  assign new_n13610_ = ~new_n13047_ & new_n13206_;
  assign new_n13611_ = ~new_n13202_ & new_n13610_;
  assign new_n13612_ = ~new_n13203_ & ~new_n13206_;
  assign new_n13613_ = ~new_n13611_ & ~new_n13612_;
  assign new_n13614_ = new_n13355_ & ~new_n13613_;
  assign new_n13615_ = ~new_n13353_ & new_n13614_;
  assign new_n13616_ = ~new_n13609_ & ~new_n13615_;
  assign new_n13617_ = ~\b[14]  & ~new_n13616_;
  assign new_n13618_ = ~new_n13046_ & ~\quotient[21] ;
  assign new_n13619_ = ~new_n13056_ & new_n13201_;
  assign new_n13620_ = ~new_n13197_ & new_n13619_;
  assign new_n13621_ = ~new_n13198_ & ~new_n13201_;
  assign new_n13622_ = ~new_n13620_ & ~new_n13621_;
  assign new_n13623_ = new_n13355_ & ~new_n13622_;
  assign new_n13624_ = ~new_n13353_ & new_n13623_;
  assign new_n13625_ = ~new_n13618_ & ~new_n13624_;
  assign new_n13626_ = ~\b[13]  & ~new_n13625_;
  assign new_n13627_ = ~new_n13055_ & ~\quotient[21] ;
  assign new_n13628_ = ~new_n13065_ & new_n13196_;
  assign new_n13629_ = ~new_n13192_ & new_n13628_;
  assign new_n13630_ = ~new_n13193_ & ~new_n13196_;
  assign new_n13631_ = ~new_n13629_ & ~new_n13630_;
  assign new_n13632_ = new_n13355_ & ~new_n13631_;
  assign new_n13633_ = ~new_n13353_ & new_n13632_;
  assign new_n13634_ = ~new_n13627_ & ~new_n13633_;
  assign new_n13635_ = ~\b[12]  & ~new_n13634_;
  assign new_n13636_ = ~new_n13064_ & ~\quotient[21] ;
  assign new_n13637_ = ~new_n13074_ & new_n13191_;
  assign new_n13638_ = ~new_n13187_ & new_n13637_;
  assign new_n13639_ = ~new_n13188_ & ~new_n13191_;
  assign new_n13640_ = ~new_n13638_ & ~new_n13639_;
  assign new_n13641_ = new_n13355_ & ~new_n13640_;
  assign new_n13642_ = ~new_n13353_ & new_n13641_;
  assign new_n13643_ = ~new_n13636_ & ~new_n13642_;
  assign new_n13644_ = ~\b[11]  & ~new_n13643_;
  assign new_n13645_ = ~new_n13073_ & ~\quotient[21] ;
  assign new_n13646_ = ~new_n13083_ & new_n13186_;
  assign new_n13647_ = ~new_n13182_ & new_n13646_;
  assign new_n13648_ = ~new_n13183_ & ~new_n13186_;
  assign new_n13649_ = ~new_n13647_ & ~new_n13648_;
  assign new_n13650_ = new_n13355_ & ~new_n13649_;
  assign new_n13651_ = ~new_n13353_ & new_n13650_;
  assign new_n13652_ = ~new_n13645_ & ~new_n13651_;
  assign new_n13653_ = ~\b[10]  & ~new_n13652_;
  assign new_n13654_ = ~new_n13082_ & ~\quotient[21] ;
  assign new_n13655_ = ~new_n13092_ & new_n13181_;
  assign new_n13656_ = ~new_n13177_ & new_n13655_;
  assign new_n13657_ = ~new_n13178_ & ~new_n13181_;
  assign new_n13658_ = ~new_n13656_ & ~new_n13657_;
  assign new_n13659_ = new_n13355_ & ~new_n13658_;
  assign new_n13660_ = ~new_n13353_ & new_n13659_;
  assign new_n13661_ = ~new_n13654_ & ~new_n13660_;
  assign new_n13662_ = ~\b[9]  & ~new_n13661_;
  assign new_n13663_ = ~new_n13091_ & ~\quotient[21] ;
  assign new_n13664_ = ~new_n13101_ & new_n13176_;
  assign new_n13665_ = ~new_n13172_ & new_n13664_;
  assign new_n13666_ = ~new_n13173_ & ~new_n13176_;
  assign new_n13667_ = ~new_n13665_ & ~new_n13666_;
  assign new_n13668_ = new_n13355_ & ~new_n13667_;
  assign new_n13669_ = ~new_n13353_ & new_n13668_;
  assign new_n13670_ = ~new_n13663_ & ~new_n13669_;
  assign new_n13671_ = ~\b[8]  & ~new_n13670_;
  assign new_n13672_ = ~new_n13100_ & ~\quotient[21] ;
  assign new_n13673_ = ~new_n13110_ & new_n13171_;
  assign new_n13674_ = ~new_n13167_ & new_n13673_;
  assign new_n13675_ = ~new_n13168_ & ~new_n13171_;
  assign new_n13676_ = ~new_n13674_ & ~new_n13675_;
  assign new_n13677_ = new_n13355_ & ~new_n13676_;
  assign new_n13678_ = ~new_n13353_ & new_n13677_;
  assign new_n13679_ = ~new_n13672_ & ~new_n13678_;
  assign new_n13680_ = ~\b[7]  & ~new_n13679_;
  assign new_n13681_ = ~new_n13109_ & ~\quotient[21] ;
  assign new_n13682_ = ~new_n13119_ & new_n13166_;
  assign new_n13683_ = ~new_n13162_ & new_n13682_;
  assign new_n13684_ = ~new_n13163_ & ~new_n13166_;
  assign new_n13685_ = ~new_n13683_ & ~new_n13684_;
  assign new_n13686_ = new_n13355_ & ~new_n13685_;
  assign new_n13687_ = ~new_n13353_ & new_n13686_;
  assign new_n13688_ = ~new_n13681_ & ~new_n13687_;
  assign new_n13689_ = ~\b[6]  & ~new_n13688_;
  assign new_n13690_ = ~new_n13118_ & ~\quotient[21] ;
  assign new_n13691_ = ~new_n13128_ & new_n13161_;
  assign new_n13692_ = ~new_n13157_ & new_n13691_;
  assign new_n13693_ = ~new_n13158_ & ~new_n13161_;
  assign new_n13694_ = ~new_n13692_ & ~new_n13693_;
  assign new_n13695_ = new_n13355_ & ~new_n13694_;
  assign new_n13696_ = ~new_n13353_ & new_n13695_;
  assign new_n13697_ = ~new_n13690_ & ~new_n13696_;
  assign new_n13698_ = ~\b[5]  & ~new_n13697_;
  assign new_n13699_ = ~new_n13127_ & ~\quotient[21] ;
  assign new_n13700_ = ~new_n13136_ & new_n13156_;
  assign new_n13701_ = ~new_n13152_ & new_n13700_;
  assign new_n13702_ = ~new_n13153_ & ~new_n13156_;
  assign new_n13703_ = ~new_n13701_ & ~new_n13702_;
  assign new_n13704_ = new_n13355_ & ~new_n13703_;
  assign new_n13705_ = ~new_n13353_ & new_n13704_;
  assign new_n13706_ = ~new_n13699_ & ~new_n13705_;
  assign new_n13707_ = ~\b[4]  & ~new_n13706_;
  assign new_n13708_ = ~new_n13135_ & ~\quotient[21] ;
  assign new_n13709_ = ~new_n13147_ & new_n13151_;
  assign new_n13710_ = ~new_n13146_ & new_n13709_;
  assign new_n13711_ = ~new_n13148_ & ~new_n13151_;
  assign new_n13712_ = ~new_n13710_ & ~new_n13711_;
  assign new_n13713_ = new_n13355_ & ~new_n13712_;
  assign new_n13714_ = ~new_n13353_ & new_n13713_;
  assign new_n13715_ = ~new_n13708_ & ~new_n13714_;
  assign new_n13716_ = ~\b[3]  & ~new_n13715_;
  assign new_n13717_ = ~new_n13140_ & ~\quotient[21] ;
  assign new_n13718_ = ~new_n13143_ & new_n13145_;
  assign new_n13719_ = ~new_n13141_ & new_n13718_;
  assign new_n13720_ = new_n13355_ & ~new_n13719_;
  assign new_n13721_ = ~new_n13146_ & new_n13720_;
  assign new_n13722_ = ~new_n13353_ & new_n13721_;
  assign new_n13723_ = ~new_n13717_ & ~new_n13722_;
  assign new_n13724_ = ~\b[2]  & ~new_n13723_;
  assign new_n13725_ = \b[0]  & ~\b[43] ;
  assign new_n13726_ = new_n301_ & new_n13725_;
  assign new_n13727_ = new_n338_ & new_n13726_;
  assign new_n13728_ = ~new_n13353_ & new_n13727_;
  assign new_n13729_ = \a[21]  & ~new_n13728_;
  assign new_n13730_ = new_n420_ & new_n13145_;
  assign new_n13731_ = new_n418_ & new_n13730_;
  assign new_n13732_ = new_n408_ & new_n13731_;
  assign new_n13733_ = ~new_n13353_ & new_n13732_;
  assign new_n13734_ = ~new_n13729_ & ~new_n13733_;
  assign new_n13735_ = \b[1]  & ~new_n13734_;
  assign new_n13736_ = ~\b[1]  & ~new_n13733_;
  assign new_n13737_ = ~new_n13729_ & new_n13736_;
  assign new_n13738_ = ~new_n13735_ & ~new_n13737_;
  assign new_n13739_ = ~\a[20]  & \b[0] ;
  assign new_n13740_ = ~new_n13738_ & ~new_n13739_;
  assign new_n13741_ = ~\b[1]  & ~new_n13734_;
  assign new_n13742_ = ~new_n13740_ & ~new_n13741_;
  assign new_n13743_ = \b[2]  & ~new_n13722_;
  assign new_n13744_ = ~new_n13717_ & new_n13743_;
  assign new_n13745_ = ~new_n13724_ & ~new_n13744_;
  assign new_n13746_ = ~new_n13742_ & new_n13745_;
  assign new_n13747_ = ~new_n13724_ & ~new_n13746_;
  assign new_n13748_ = \b[3]  & ~new_n13714_;
  assign new_n13749_ = ~new_n13708_ & new_n13748_;
  assign new_n13750_ = ~new_n13716_ & ~new_n13749_;
  assign new_n13751_ = ~new_n13747_ & new_n13750_;
  assign new_n13752_ = ~new_n13716_ & ~new_n13751_;
  assign new_n13753_ = \b[4]  & ~new_n13705_;
  assign new_n13754_ = ~new_n13699_ & new_n13753_;
  assign new_n13755_ = ~new_n13707_ & ~new_n13754_;
  assign new_n13756_ = ~new_n13752_ & new_n13755_;
  assign new_n13757_ = ~new_n13707_ & ~new_n13756_;
  assign new_n13758_ = \b[5]  & ~new_n13696_;
  assign new_n13759_ = ~new_n13690_ & new_n13758_;
  assign new_n13760_ = ~new_n13698_ & ~new_n13759_;
  assign new_n13761_ = ~new_n13757_ & new_n13760_;
  assign new_n13762_ = ~new_n13698_ & ~new_n13761_;
  assign new_n13763_ = \b[6]  & ~new_n13687_;
  assign new_n13764_ = ~new_n13681_ & new_n13763_;
  assign new_n13765_ = ~new_n13689_ & ~new_n13764_;
  assign new_n13766_ = ~new_n13762_ & new_n13765_;
  assign new_n13767_ = ~new_n13689_ & ~new_n13766_;
  assign new_n13768_ = \b[7]  & ~new_n13678_;
  assign new_n13769_ = ~new_n13672_ & new_n13768_;
  assign new_n13770_ = ~new_n13680_ & ~new_n13769_;
  assign new_n13771_ = ~new_n13767_ & new_n13770_;
  assign new_n13772_ = ~new_n13680_ & ~new_n13771_;
  assign new_n13773_ = \b[8]  & ~new_n13669_;
  assign new_n13774_ = ~new_n13663_ & new_n13773_;
  assign new_n13775_ = ~new_n13671_ & ~new_n13774_;
  assign new_n13776_ = ~new_n13772_ & new_n13775_;
  assign new_n13777_ = ~new_n13671_ & ~new_n13776_;
  assign new_n13778_ = \b[9]  & ~new_n13660_;
  assign new_n13779_ = ~new_n13654_ & new_n13778_;
  assign new_n13780_ = ~new_n13662_ & ~new_n13779_;
  assign new_n13781_ = ~new_n13777_ & new_n13780_;
  assign new_n13782_ = ~new_n13662_ & ~new_n13781_;
  assign new_n13783_ = \b[10]  & ~new_n13651_;
  assign new_n13784_ = ~new_n13645_ & new_n13783_;
  assign new_n13785_ = ~new_n13653_ & ~new_n13784_;
  assign new_n13786_ = ~new_n13782_ & new_n13785_;
  assign new_n13787_ = ~new_n13653_ & ~new_n13786_;
  assign new_n13788_ = \b[11]  & ~new_n13642_;
  assign new_n13789_ = ~new_n13636_ & new_n13788_;
  assign new_n13790_ = ~new_n13644_ & ~new_n13789_;
  assign new_n13791_ = ~new_n13787_ & new_n13790_;
  assign new_n13792_ = ~new_n13644_ & ~new_n13791_;
  assign new_n13793_ = \b[12]  & ~new_n13633_;
  assign new_n13794_ = ~new_n13627_ & new_n13793_;
  assign new_n13795_ = ~new_n13635_ & ~new_n13794_;
  assign new_n13796_ = ~new_n13792_ & new_n13795_;
  assign new_n13797_ = ~new_n13635_ & ~new_n13796_;
  assign new_n13798_ = \b[13]  & ~new_n13624_;
  assign new_n13799_ = ~new_n13618_ & new_n13798_;
  assign new_n13800_ = ~new_n13626_ & ~new_n13799_;
  assign new_n13801_ = ~new_n13797_ & new_n13800_;
  assign new_n13802_ = ~new_n13626_ & ~new_n13801_;
  assign new_n13803_ = \b[14]  & ~new_n13615_;
  assign new_n13804_ = ~new_n13609_ & new_n13803_;
  assign new_n13805_ = ~new_n13617_ & ~new_n13804_;
  assign new_n13806_ = ~new_n13802_ & new_n13805_;
  assign new_n13807_ = ~new_n13617_ & ~new_n13806_;
  assign new_n13808_ = \b[15]  & ~new_n13606_;
  assign new_n13809_ = ~new_n13600_ & new_n13808_;
  assign new_n13810_ = ~new_n13608_ & ~new_n13809_;
  assign new_n13811_ = ~new_n13807_ & new_n13810_;
  assign new_n13812_ = ~new_n13608_ & ~new_n13811_;
  assign new_n13813_ = \b[16]  & ~new_n13597_;
  assign new_n13814_ = ~new_n13591_ & new_n13813_;
  assign new_n13815_ = ~new_n13599_ & ~new_n13814_;
  assign new_n13816_ = ~new_n13812_ & new_n13815_;
  assign new_n13817_ = ~new_n13599_ & ~new_n13816_;
  assign new_n13818_ = \b[17]  & ~new_n13588_;
  assign new_n13819_ = ~new_n13582_ & new_n13818_;
  assign new_n13820_ = ~new_n13590_ & ~new_n13819_;
  assign new_n13821_ = ~new_n13817_ & new_n13820_;
  assign new_n13822_ = ~new_n13590_ & ~new_n13821_;
  assign new_n13823_ = \b[18]  & ~new_n13579_;
  assign new_n13824_ = ~new_n13573_ & new_n13823_;
  assign new_n13825_ = ~new_n13581_ & ~new_n13824_;
  assign new_n13826_ = ~new_n13822_ & new_n13825_;
  assign new_n13827_ = ~new_n13581_ & ~new_n13826_;
  assign new_n13828_ = \b[19]  & ~new_n13570_;
  assign new_n13829_ = ~new_n13564_ & new_n13828_;
  assign new_n13830_ = ~new_n13572_ & ~new_n13829_;
  assign new_n13831_ = ~new_n13827_ & new_n13830_;
  assign new_n13832_ = ~new_n13572_ & ~new_n13831_;
  assign new_n13833_ = \b[20]  & ~new_n13561_;
  assign new_n13834_ = ~new_n13555_ & new_n13833_;
  assign new_n13835_ = ~new_n13563_ & ~new_n13834_;
  assign new_n13836_ = ~new_n13832_ & new_n13835_;
  assign new_n13837_ = ~new_n13563_ & ~new_n13836_;
  assign new_n13838_ = \b[21]  & ~new_n13552_;
  assign new_n13839_ = ~new_n13546_ & new_n13838_;
  assign new_n13840_ = ~new_n13554_ & ~new_n13839_;
  assign new_n13841_ = ~new_n13837_ & new_n13840_;
  assign new_n13842_ = ~new_n13554_ & ~new_n13841_;
  assign new_n13843_ = \b[22]  & ~new_n13543_;
  assign new_n13844_ = ~new_n13537_ & new_n13843_;
  assign new_n13845_ = ~new_n13545_ & ~new_n13844_;
  assign new_n13846_ = ~new_n13842_ & new_n13845_;
  assign new_n13847_ = ~new_n13545_ & ~new_n13846_;
  assign new_n13848_ = \b[23]  & ~new_n13534_;
  assign new_n13849_ = ~new_n13528_ & new_n13848_;
  assign new_n13850_ = ~new_n13536_ & ~new_n13849_;
  assign new_n13851_ = ~new_n13847_ & new_n13850_;
  assign new_n13852_ = ~new_n13536_ & ~new_n13851_;
  assign new_n13853_ = \b[24]  & ~new_n13525_;
  assign new_n13854_ = ~new_n13519_ & new_n13853_;
  assign new_n13855_ = ~new_n13527_ & ~new_n13854_;
  assign new_n13856_ = ~new_n13852_ & new_n13855_;
  assign new_n13857_ = ~new_n13527_ & ~new_n13856_;
  assign new_n13858_ = \b[25]  & ~new_n13516_;
  assign new_n13859_ = ~new_n13510_ & new_n13858_;
  assign new_n13860_ = ~new_n13518_ & ~new_n13859_;
  assign new_n13861_ = ~new_n13857_ & new_n13860_;
  assign new_n13862_ = ~new_n13518_ & ~new_n13861_;
  assign new_n13863_ = \b[26]  & ~new_n13507_;
  assign new_n13864_ = ~new_n13501_ & new_n13863_;
  assign new_n13865_ = ~new_n13509_ & ~new_n13864_;
  assign new_n13866_ = ~new_n13862_ & new_n13865_;
  assign new_n13867_ = ~new_n13509_ & ~new_n13866_;
  assign new_n13868_ = \b[27]  & ~new_n13498_;
  assign new_n13869_ = ~new_n13492_ & new_n13868_;
  assign new_n13870_ = ~new_n13500_ & ~new_n13869_;
  assign new_n13871_ = ~new_n13867_ & new_n13870_;
  assign new_n13872_ = ~new_n13500_ & ~new_n13871_;
  assign new_n13873_ = \b[28]  & ~new_n13489_;
  assign new_n13874_ = ~new_n13483_ & new_n13873_;
  assign new_n13875_ = ~new_n13491_ & ~new_n13874_;
  assign new_n13876_ = ~new_n13872_ & new_n13875_;
  assign new_n13877_ = ~new_n13491_ & ~new_n13876_;
  assign new_n13878_ = \b[29]  & ~new_n13480_;
  assign new_n13879_ = ~new_n13474_ & new_n13878_;
  assign new_n13880_ = ~new_n13482_ & ~new_n13879_;
  assign new_n13881_ = ~new_n13877_ & new_n13880_;
  assign new_n13882_ = ~new_n13482_ & ~new_n13881_;
  assign new_n13883_ = \b[30]  & ~new_n13471_;
  assign new_n13884_ = ~new_n13465_ & new_n13883_;
  assign new_n13885_ = ~new_n13473_ & ~new_n13884_;
  assign new_n13886_ = ~new_n13882_ & new_n13885_;
  assign new_n13887_ = ~new_n13473_ & ~new_n13886_;
  assign new_n13888_ = \b[31]  & ~new_n13462_;
  assign new_n13889_ = ~new_n13456_ & new_n13888_;
  assign new_n13890_ = ~new_n13464_ & ~new_n13889_;
  assign new_n13891_ = ~new_n13887_ & new_n13890_;
  assign new_n13892_ = ~new_n13464_ & ~new_n13891_;
  assign new_n13893_ = \b[32]  & ~new_n13453_;
  assign new_n13894_ = ~new_n13447_ & new_n13893_;
  assign new_n13895_ = ~new_n13455_ & ~new_n13894_;
  assign new_n13896_ = ~new_n13892_ & new_n13895_;
  assign new_n13897_ = ~new_n13455_ & ~new_n13896_;
  assign new_n13898_ = \b[33]  & ~new_n13444_;
  assign new_n13899_ = ~new_n13438_ & new_n13898_;
  assign new_n13900_ = ~new_n13446_ & ~new_n13899_;
  assign new_n13901_ = ~new_n13897_ & new_n13900_;
  assign new_n13902_ = ~new_n13446_ & ~new_n13901_;
  assign new_n13903_ = \b[34]  & ~new_n13435_;
  assign new_n13904_ = ~new_n13429_ & new_n13903_;
  assign new_n13905_ = ~new_n13437_ & ~new_n13904_;
  assign new_n13906_ = ~new_n13902_ & new_n13905_;
  assign new_n13907_ = ~new_n13437_ & ~new_n13906_;
  assign new_n13908_ = \b[35]  & ~new_n13426_;
  assign new_n13909_ = ~new_n13420_ & new_n13908_;
  assign new_n13910_ = ~new_n13428_ & ~new_n13909_;
  assign new_n13911_ = ~new_n13907_ & new_n13910_;
  assign new_n13912_ = ~new_n13428_ & ~new_n13911_;
  assign new_n13913_ = \b[36]  & ~new_n13417_;
  assign new_n13914_ = ~new_n13411_ & new_n13913_;
  assign new_n13915_ = ~new_n13419_ & ~new_n13914_;
  assign new_n13916_ = ~new_n13912_ & new_n13915_;
  assign new_n13917_ = ~new_n13419_ & ~new_n13916_;
  assign new_n13918_ = \b[37]  & ~new_n13408_;
  assign new_n13919_ = ~new_n13402_ & new_n13918_;
  assign new_n13920_ = ~new_n13410_ & ~new_n13919_;
  assign new_n13921_ = ~new_n13917_ & new_n13920_;
  assign new_n13922_ = ~new_n13410_ & ~new_n13921_;
  assign new_n13923_ = \b[38]  & ~new_n13399_;
  assign new_n13924_ = ~new_n13393_ & new_n13923_;
  assign new_n13925_ = ~new_n13401_ & ~new_n13924_;
  assign new_n13926_ = ~new_n13922_ & new_n13925_;
  assign new_n13927_ = ~new_n13401_ & ~new_n13926_;
  assign new_n13928_ = \b[39]  & ~new_n13390_;
  assign new_n13929_ = ~new_n13384_ & new_n13928_;
  assign new_n13930_ = ~new_n13392_ & ~new_n13929_;
  assign new_n13931_ = ~new_n13927_ & new_n13930_;
  assign new_n13932_ = ~new_n13392_ & ~new_n13931_;
  assign new_n13933_ = \b[40]  & ~new_n13381_;
  assign new_n13934_ = ~new_n13375_ & new_n13933_;
  assign new_n13935_ = ~new_n13383_ & ~new_n13934_;
  assign new_n13936_ = ~new_n13932_ & new_n13935_;
  assign new_n13937_ = ~new_n13383_ & ~new_n13936_;
  assign new_n13938_ = \b[41]  & ~new_n13372_;
  assign new_n13939_ = ~new_n13366_ & new_n13938_;
  assign new_n13940_ = ~new_n13374_ & ~new_n13939_;
  assign new_n13941_ = ~new_n13937_ & new_n13940_;
  assign new_n13942_ = ~new_n13374_ & ~new_n13941_;
  assign new_n13943_ = \b[42]  & ~new_n13363_;
  assign new_n13944_ = ~new_n13357_ & new_n13943_;
  assign new_n13945_ = ~new_n13365_ & ~new_n13944_;
  assign new_n13946_ = ~new_n13942_ & new_n13945_;
  assign new_n13947_ = ~new_n13365_ & ~new_n13946_;
  assign new_n13948_ = ~new_n12784_ & ~\quotient[21] ;
  assign new_n13949_ = ~new_n12786_ & new_n13351_;
  assign new_n13950_ = ~new_n13347_ & new_n13949_;
  assign new_n13951_ = ~new_n13348_ & ~new_n13351_;
  assign new_n13952_ = ~new_n13950_ & ~new_n13951_;
  assign new_n13953_ = \quotient[21]  & ~new_n13952_;
  assign new_n13954_ = ~new_n13948_ & ~new_n13953_;
  assign new_n13955_ = ~\b[43]  & ~new_n13954_;
  assign new_n13956_ = \b[43]  & ~new_n13948_;
  assign new_n13957_ = ~new_n13953_ & new_n13956_;
  assign new_n13958_ = new_n288_ & new_n302_;
  assign new_n13959_ = ~new_n13957_ & new_n13958_;
  assign new_n13960_ = ~new_n13955_ & new_n13959_;
  assign new_n13961_ = ~new_n13947_ & new_n13960_;
  assign new_n13962_ = new_n13355_ & ~new_n13954_;
  assign \quotient[20]  = new_n13961_ | new_n13962_;
  assign new_n13964_ = ~new_n13374_ & new_n13945_;
  assign new_n13965_ = ~new_n13941_ & new_n13964_;
  assign new_n13966_ = ~new_n13942_ & ~new_n13945_;
  assign new_n13967_ = ~new_n13965_ & ~new_n13966_;
  assign new_n13968_ = \quotient[20]  & ~new_n13967_;
  assign new_n13969_ = ~new_n13364_ & ~new_n13962_;
  assign new_n13970_ = ~new_n13961_ & new_n13969_;
  assign new_n13971_ = ~new_n13968_ & ~new_n13970_;
  assign new_n13972_ = ~\b[43]  & ~new_n13971_;
  assign new_n13973_ = ~new_n13383_ & new_n13940_;
  assign new_n13974_ = ~new_n13936_ & new_n13973_;
  assign new_n13975_ = ~new_n13937_ & ~new_n13940_;
  assign new_n13976_ = ~new_n13974_ & ~new_n13975_;
  assign new_n13977_ = \quotient[20]  & ~new_n13976_;
  assign new_n13978_ = ~new_n13373_ & ~new_n13962_;
  assign new_n13979_ = ~new_n13961_ & new_n13978_;
  assign new_n13980_ = ~new_n13977_ & ~new_n13979_;
  assign new_n13981_ = ~\b[42]  & ~new_n13980_;
  assign new_n13982_ = ~new_n13392_ & new_n13935_;
  assign new_n13983_ = ~new_n13931_ & new_n13982_;
  assign new_n13984_ = ~new_n13932_ & ~new_n13935_;
  assign new_n13985_ = ~new_n13983_ & ~new_n13984_;
  assign new_n13986_ = \quotient[20]  & ~new_n13985_;
  assign new_n13987_ = ~new_n13382_ & ~new_n13962_;
  assign new_n13988_ = ~new_n13961_ & new_n13987_;
  assign new_n13989_ = ~new_n13986_ & ~new_n13988_;
  assign new_n13990_ = ~\b[41]  & ~new_n13989_;
  assign new_n13991_ = ~new_n13401_ & new_n13930_;
  assign new_n13992_ = ~new_n13926_ & new_n13991_;
  assign new_n13993_ = ~new_n13927_ & ~new_n13930_;
  assign new_n13994_ = ~new_n13992_ & ~new_n13993_;
  assign new_n13995_ = \quotient[20]  & ~new_n13994_;
  assign new_n13996_ = ~new_n13391_ & ~new_n13962_;
  assign new_n13997_ = ~new_n13961_ & new_n13996_;
  assign new_n13998_ = ~new_n13995_ & ~new_n13997_;
  assign new_n13999_ = ~\b[40]  & ~new_n13998_;
  assign new_n14000_ = ~new_n13410_ & new_n13925_;
  assign new_n14001_ = ~new_n13921_ & new_n14000_;
  assign new_n14002_ = ~new_n13922_ & ~new_n13925_;
  assign new_n14003_ = ~new_n14001_ & ~new_n14002_;
  assign new_n14004_ = \quotient[20]  & ~new_n14003_;
  assign new_n14005_ = ~new_n13400_ & ~new_n13962_;
  assign new_n14006_ = ~new_n13961_ & new_n14005_;
  assign new_n14007_ = ~new_n14004_ & ~new_n14006_;
  assign new_n14008_ = ~\b[39]  & ~new_n14007_;
  assign new_n14009_ = ~new_n13419_ & new_n13920_;
  assign new_n14010_ = ~new_n13916_ & new_n14009_;
  assign new_n14011_ = ~new_n13917_ & ~new_n13920_;
  assign new_n14012_ = ~new_n14010_ & ~new_n14011_;
  assign new_n14013_ = \quotient[20]  & ~new_n14012_;
  assign new_n14014_ = ~new_n13409_ & ~new_n13962_;
  assign new_n14015_ = ~new_n13961_ & new_n14014_;
  assign new_n14016_ = ~new_n14013_ & ~new_n14015_;
  assign new_n14017_ = ~\b[38]  & ~new_n14016_;
  assign new_n14018_ = ~new_n13428_ & new_n13915_;
  assign new_n14019_ = ~new_n13911_ & new_n14018_;
  assign new_n14020_ = ~new_n13912_ & ~new_n13915_;
  assign new_n14021_ = ~new_n14019_ & ~new_n14020_;
  assign new_n14022_ = \quotient[20]  & ~new_n14021_;
  assign new_n14023_ = ~new_n13418_ & ~new_n13962_;
  assign new_n14024_ = ~new_n13961_ & new_n14023_;
  assign new_n14025_ = ~new_n14022_ & ~new_n14024_;
  assign new_n14026_ = ~\b[37]  & ~new_n14025_;
  assign new_n14027_ = ~new_n13437_ & new_n13910_;
  assign new_n14028_ = ~new_n13906_ & new_n14027_;
  assign new_n14029_ = ~new_n13907_ & ~new_n13910_;
  assign new_n14030_ = ~new_n14028_ & ~new_n14029_;
  assign new_n14031_ = \quotient[20]  & ~new_n14030_;
  assign new_n14032_ = ~new_n13427_ & ~new_n13962_;
  assign new_n14033_ = ~new_n13961_ & new_n14032_;
  assign new_n14034_ = ~new_n14031_ & ~new_n14033_;
  assign new_n14035_ = ~\b[36]  & ~new_n14034_;
  assign new_n14036_ = ~new_n13446_ & new_n13905_;
  assign new_n14037_ = ~new_n13901_ & new_n14036_;
  assign new_n14038_ = ~new_n13902_ & ~new_n13905_;
  assign new_n14039_ = ~new_n14037_ & ~new_n14038_;
  assign new_n14040_ = \quotient[20]  & ~new_n14039_;
  assign new_n14041_ = ~new_n13436_ & ~new_n13962_;
  assign new_n14042_ = ~new_n13961_ & new_n14041_;
  assign new_n14043_ = ~new_n14040_ & ~new_n14042_;
  assign new_n14044_ = ~\b[35]  & ~new_n14043_;
  assign new_n14045_ = ~new_n13455_ & new_n13900_;
  assign new_n14046_ = ~new_n13896_ & new_n14045_;
  assign new_n14047_ = ~new_n13897_ & ~new_n13900_;
  assign new_n14048_ = ~new_n14046_ & ~new_n14047_;
  assign new_n14049_ = \quotient[20]  & ~new_n14048_;
  assign new_n14050_ = ~new_n13445_ & ~new_n13962_;
  assign new_n14051_ = ~new_n13961_ & new_n14050_;
  assign new_n14052_ = ~new_n14049_ & ~new_n14051_;
  assign new_n14053_ = ~\b[34]  & ~new_n14052_;
  assign new_n14054_ = ~new_n13464_ & new_n13895_;
  assign new_n14055_ = ~new_n13891_ & new_n14054_;
  assign new_n14056_ = ~new_n13892_ & ~new_n13895_;
  assign new_n14057_ = ~new_n14055_ & ~new_n14056_;
  assign new_n14058_ = \quotient[20]  & ~new_n14057_;
  assign new_n14059_ = ~new_n13454_ & ~new_n13962_;
  assign new_n14060_ = ~new_n13961_ & new_n14059_;
  assign new_n14061_ = ~new_n14058_ & ~new_n14060_;
  assign new_n14062_ = ~\b[33]  & ~new_n14061_;
  assign new_n14063_ = ~new_n13473_ & new_n13890_;
  assign new_n14064_ = ~new_n13886_ & new_n14063_;
  assign new_n14065_ = ~new_n13887_ & ~new_n13890_;
  assign new_n14066_ = ~new_n14064_ & ~new_n14065_;
  assign new_n14067_ = \quotient[20]  & ~new_n14066_;
  assign new_n14068_ = ~new_n13463_ & ~new_n13962_;
  assign new_n14069_ = ~new_n13961_ & new_n14068_;
  assign new_n14070_ = ~new_n14067_ & ~new_n14069_;
  assign new_n14071_ = ~\b[32]  & ~new_n14070_;
  assign new_n14072_ = ~new_n13482_ & new_n13885_;
  assign new_n14073_ = ~new_n13881_ & new_n14072_;
  assign new_n14074_ = ~new_n13882_ & ~new_n13885_;
  assign new_n14075_ = ~new_n14073_ & ~new_n14074_;
  assign new_n14076_ = \quotient[20]  & ~new_n14075_;
  assign new_n14077_ = ~new_n13472_ & ~new_n13962_;
  assign new_n14078_ = ~new_n13961_ & new_n14077_;
  assign new_n14079_ = ~new_n14076_ & ~new_n14078_;
  assign new_n14080_ = ~\b[31]  & ~new_n14079_;
  assign new_n14081_ = ~new_n13491_ & new_n13880_;
  assign new_n14082_ = ~new_n13876_ & new_n14081_;
  assign new_n14083_ = ~new_n13877_ & ~new_n13880_;
  assign new_n14084_ = ~new_n14082_ & ~new_n14083_;
  assign new_n14085_ = \quotient[20]  & ~new_n14084_;
  assign new_n14086_ = ~new_n13481_ & ~new_n13962_;
  assign new_n14087_ = ~new_n13961_ & new_n14086_;
  assign new_n14088_ = ~new_n14085_ & ~new_n14087_;
  assign new_n14089_ = ~\b[30]  & ~new_n14088_;
  assign new_n14090_ = ~new_n13500_ & new_n13875_;
  assign new_n14091_ = ~new_n13871_ & new_n14090_;
  assign new_n14092_ = ~new_n13872_ & ~new_n13875_;
  assign new_n14093_ = ~new_n14091_ & ~new_n14092_;
  assign new_n14094_ = \quotient[20]  & ~new_n14093_;
  assign new_n14095_ = ~new_n13490_ & ~new_n13962_;
  assign new_n14096_ = ~new_n13961_ & new_n14095_;
  assign new_n14097_ = ~new_n14094_ & ~new_n14096_;
  assign new_n14098_ = ~\b[29]  & ~new_n14097_;
  assign new_n14099_ = ~new_n13509_ & new_n13870_;
  assign new_n14100_ = ~new_n13866_ & new_n14099_;
  assign new_n14101_ = ~new_n13867_ & ~new_n13870_;
  assign new_n14102_ = ~new_n14100_ & ~new_n14101_;
  assign new_n14103_ = \quotient[20]  & ~new_n14102_;
  assign new_n14104_ = ~new_n13499_ & ~new_n13962_;
  assign new_n14105_ = ~new_n13961_ & new_n14104_;
  assign new_n14106_ = ~new_n14103_ & ~new_n14105_;
  assign new_n14107_ = ~\b[28]  & ~new_n14106_;
  assign new_n14108_ = ~new_n13518_ & new_n13865_;
  assign new_n14109_ = ~new_n13861_ & new_n14108_;
  assign new_n14110_ = ~new_n13862_ & ~new_n13865_;
  assign new_n14111_ = ~new_n14109_ & ~new_n14110_;
  assign new_n14112_ = \quotient[20]  & ~new_n14111_;
  assign new_n14113_ = ~new_n13508_ & ~new_n13962_;
  assign new_n14114_ = ~new_n13961_ & new_n14113_;
  assign new_n14115_ = ~new_n14112_ & ~new_n14114_;
  assign new_n14116_ = ~\b[27]  & ~new_n14115_;
  assign new_n14117_ = ~new_n13527_ & new_n13860_;
  assign new_n14118_ = ~new_n13856_ & new_n14117_;
  assign new_n14119_ = ~new_n13857_ & ~new_n13860_;
  assign new_n14120_ = ~new_n14118_ & ~new_n14119_;
  assign new_n14121_ = \quotient[20]  & ~new_n14120_;
  assign new_n14122_ = ~new_n13517_ & ~new_n13962_;
  assign new_n14123_ = ~new_n13961_ & new_n14122_;
  assign new_n14124_ = ~new_n14121_ & ~new_n14123_;
  assign new_n14125_ = ~\b[26]  & ~new_n14124_;
  assign new_n14126_ = ~new_n13536_ & new_n13855_;
  assign new_n14127_ = ~new_n13851_ & new_n14126_;
  assign new_n14128_ = ~new_n13852_ & ~new_n13855_;
  assign new_n14129_ = ~new_n14127_ & ~new_n14128_;
  assign new_n14130_ = \quotient[20]  & ~new_n14129_;
  assign new_n14131_ = ~new_n13526_ & ~new_n13962_;
  assign new_n14132_ = ~new_n13961_ & new_n14131_;
  assign new_n14133_ = ~new_n14130_ & ~new_n14132_;
  assign new_n14134_ = ~\b[25]  & ~new_n14133_;
  assign new_n14135_ = ~new_n13545_ & new_n13850_;
  assign new_n14136_ = ~new_n13846_ & new_n14135_;
  assign new_n14137_ = ~new_n13847_ & ~new_n13850_;
  assign new_n14138_ = ~new_n14136_ & ~new_n14137_;
  assign new_n14139_ = \quotient[20]  & ~new_n14138_;
  assign new_n14140_ = ~new_n13535_ & ~new_n13962_;
  assign new_n14141_ = ~new_n13961_ & new_n14140_;
  assign new_n14142_ = ~new_n14139_ & ~new_n14141_;
  assign new_n14143_ = ~\b[24]  & ~new_n14142_;
  assign new_n14144_ = ~new_n13554_ & new_n13845_;
  assign new_n14145_ = ~new_n13841_ & new_n14144_;
  assign new_n14146_ = ~new_n13842_ & ~new_n13845_;
  assign new_n14147_ = ~new_n14145_ & ~new_n14146_;
  assign new_n14148_ = \quotient[20]  & ~new_n14147_;
  assign new_n14149_ = ~new_n13544_ & ~new_n13962_;
  assign new_n14150_ = ~new_n13961_ & new_n14149_;
  assign new_n14151_ = ~new_n14148_ & ~new_n14150_;
  assign new_n14152_ = ~\b[23]  & ~new_n14151_;
  assign new_n14153_ = ~new_n13563_ & new_n13840_;
  assign new_n14154_ = ~new_n13836_ & new_n14153_;
  assign new_n14155_ = ~new_n13837_ & ~new_n13840_;
  assign new_n14156_ = ~new_n14154_ & ~new_n14155_;
  assign new_n14157_ = \quotient[20]  & ~new_n14156_;
  assign new_n14158_ = ~new_n13553_ & ~new_n13962_;
  assign new_n14159_ = ~new_n13961_ & new_n14158_;
  assign new_n14160_ = ~new_n14157_ & ~new_n14159_;
  assign new_n14161_ = ~\b[22]  & ~new_n14160_;
  assign new_n14162_ = ~new_n13572_ & new_n13835_;
  assign new_n14163_ = ~new_n13831_ & new_n14162_;
  assign new_n14164_ = ~new_n13832_ & ~new_n13835_;
  assign new_n14165_ = ~new_n14163_ & ~new_n14164_;
  assign new_n14166_ = \quotient[20]  & ~new_n14165_;
  assign new_n14167_ = ~new_n13562_ & ~new_n13962_;
  assign new_n14168_ = ~new_n13961_ & new_n14167_;
  assign new_n14169_ = ~new_n14166_ & ~new_n14168_;
  assign new_n14170_ = ~\b[21]  & ~new_n14169_;
  assign new_n14171_ = ~new_n13581_ & new_n13830_;
  assign new_n14172_ = ~new_n13826_ & new_n14171_;
  assign new_n14173_ = ~new_n13827_ & ~new_n13830_;
  assign new_n14174_ = ~new_n14172_ & ~new_n14173_;
  assign new_n14175_ = \quotient[20]  & ~new_n14174_;
  assign new_n14176_ = ~new_n13571_ & ~new_n13962_;
  assign new_n14177_ = ~new_n13961_ & new_n14176_;
  assign new_n14178_ = ~new_n14175_ & ~new_n14177_;
  assign new_n14179_ = ~\b[20]  & ~new_n14178_;
  assign new_n14180_ = ~new_n13590_ & new_n13825_;
  assign new_n14181_ = ~new_n13821_ & new_n14180_;
  assign new_n14182_ = ~new_n13822_ & ~new_n13825_;
  assign new_n14183_ = ~new_n14181_ & ~new_n14182_;
  assign new_n14184_ = \quotient[20]  & ~new_n14183_;
  assign new_n14185_ = ~new_n13580_ & ~new_n13962_;
  assign new_n14186_ = ~new_n13961_ & new_n14185_;
  assign new_n14187_ = ~new_n14184_ & ~new_n14186_;
  assign new_n14188_ = ~\b[19]  & ~new_n14187_;
  assign new_n14189_ = ~new_n13599_ & new_n13820_;
  assign new_n14190_ = ~new_n13816_ & new_n14189_;
  assign new_n14191_ = ~new_n13817_ & ~new_n13820_;
  assign new_n14192_ = ~new_n14190_ & ~new_n14191_;
  assign new_n14193_ = \quotient[20]  & ~new_n14192_;
  assign new_n14194_ = ~new_n13589_ & ~new_n13962_;
  assign new_n14195_ = ~new_n13961_ & new_n14194_;
  assign new_n14196_ = ~new_n14193_ & ~new_n14195_;
  assign new_n14197_ = ~\b[18]  & ~new_n14196_;
  assign new_n14198_ = ~new_n13608_ & new_n13815_;
  assign new_n14199_ = ~new_n13811_ & new_n14198_;
  assign new_n14200_ = ~new_n13812_ & ~new_n13815_;
  assign new_n14201_ = ~new_n14199_ & ~new_n14200_;
  assign new_n14202_ = \quotient[20]  & ~new_n14201_;
  assign new_n14203_ = ~new_n13598_ & ~new_n13962_;
  assign new_n14204_ = ~new_n13961_ & new_n14203_;
  assign new_n14205_ = ~new_n14202_ & ~new_n14204_;
  assign new_n14206_ = ~\b[17]  & ~new_n14205_;
  assign new_n14207_ = ~new_n13617_ & new_n13810_;
  assign new_n14208_ = ~new_n13806_ & new_n14207_;
  assign new_n14209_ = ~new_n13807_ & ~new_n13810_;
  assign new_n14210_ = ~new_n14208_ & ~new_n14209_;
  assign new_n14211_ = \quotient[20]  & ~new_n14210_;
  assign new_n14212_ = ~new_n13607_ & ~new_n13962_;
  assign new_n14213_ = ~new_n13961_ & new_n14212_;
  assign new_n14214_ = ~new_n14211_ & ~new_n14213_;
  assign new_n14215_ = ~\b[16]  & ~new_n14214_;
  assign new_n14216_ = ~new_n13626_ & new_n13805_;
  assign new_n14217_ = ~new_n13801_ & new_n14216_;
  assign new_n14218_ = ~new_n13802_ & ~new_n13805_;
  assign new_n14219_ = ~new_n14217_ & ~new_n14218_;
  assign new_n14220_ = \quotient[20]  & ~new_n14219_;
  assign new_n14221_ = ~new_n13616_ & ~new_n13962_;
  assign new_n14222_ = ~new_n13961_ & new_n14221_;
  assign new_n14223_ = ~new_n14220_ & ~new_n14222_;
  assign new_n14224_ = ~\b[15]  & ~new_n14223_;
  assign new_n14225_ = ~new_n13635_ & new_n13800_;
  assign new_n14226_ = ~new_n13796_ & new_n14225_;
  assign new_n14227_ = ~new_n13797_ & ~new_n13800_;
  assign new_n14228_ = ~new_n14226_ & ~new_n14227_;
  assign new_n14229_ = \quotient[20]  & ~new_n14228_;
  assign new_n14230_ = ~new_n13625_ & ~new_n13962_;
  assign new_n14231_ = ~new_n13961_ & new_n14230_;
  assign new_n14232_ = ~new_n14229_ & ~new_n14231_;
  assign new_n14233_ = ~\b[14]  & ~new_n14232_;
  assign new_n14234_ = ~new_n13644_ & new_n13795_;
  assign new_n14235_ = ~new_n13791_ & new_n14234_;
  assign new_n14236_ = ~new_n13792_ & ~new_n13795_;
  assign new_n14237_ = ~new_n14235_ & ~new_n14236_;
  assign new_n14238_ = \quotient[20]  & ~new_n14237_;
  assign new_n14239_ = ~new_n13634_ & ~new_n13962_;
  assign new_n14240_ = ~new_n13961_ & new_n14239_;
  assign new_n14241_ = ~new_n14238_ & ~new_n14240_;
  assign new_n14242_ = ~\b[13]  & ~new_n14241_;
  assign new_n14243_ = ~new_n13653_ & new_n13790_;
  assign new_n14244_ = ~new_n13786_ & new_n14243_;
  assign new_n14245_ = ~new_n13787_ & ~new_n13790_;
  assign new_n14246_ = ~new_n14244_ & ~new_n14245_;
  assign new_n14247_ = \quotient[20]  & ~new_n14246_;
  assign new_n14248_ = ~new_n13643_ & ~new_n13962_;
  assign new_n14249_ = ~new_n13961_ & new_n14248_;
  assign new_n14250_ = ~new_n14247_ & ~new_n14249_;
  assign new_n14251_ = ~\b[12]  & ~new_n14250_;
  assign new_n14252_ = ~new_n13662_ & new_n13785_;
  assign new_n14253_ = ~new_n13781_ & new_n14252_;
  assign new_n14254_ = ~new_n13782_ & ~new_n13785_;
  assign new_n14255_ = ~new_n14253_ & ~new_n14254_;
  assign new_n14256_ = \quotient[20]  & ~new_n14255_;
  assign new_n14257_ = ~new_n13652_ & ~new_n13962_;
  assign new_n14258_ = ~new_n13961_ & new_n14257_;
  assign new_n14259_ = ~new_n14256_ & ~new_n14258_;
  assign new_n14260_ = ~\b[11]  & ~new_n14259_;
  assign new_n14261_ = ~new_n13671_ & new_n13780_;
  assign new_n14262_ = ~new_n13776_ & new_n14261_;
  assign new_n14263_ = ~new_n13777_ & ~new_n13780_;
  assign new_n14264_ = ~new_n14262_ & ~new_n14263_;
  assign new_n14265_ = \quotient[20]  & ~new_n14264_;
  assign new_n14266_ = ~new_n13661_ & ~new_n13962_;
  assign new_n14267_ = ~new_n13961_ & new_n14266_;
  assign new_n14268_ = ~new_n14265_ & ~new_n14267_;
  assign new_n14269_ = ~\b[10]  & ~new_n14268_;
  assign new_n14270_ = ~new_n13680_ & new_n13775_;
  assign new_n14271_ = ~new_n13771_ & new_n14270_;
  assign new_n14272_ = ~new_n13772_ & ~new_n13775_;
  assign new_n14273_ = ~new_n14271_ & ~new_n14272_;
  assign new_n14274_ = \quotient[20]  & ~new_n14273_;
  assign new_n14275_ = ~new_n13670_ & ~new_n13962_;
  assign new_n14276_ = ~new_n13961_ & new_n14275_;
  assign new_n14277_ = ~new_n14274_ & ~new_n14276_;
  assign new_n14278_ = ~\b[9]  & ~new_n14277_;
  assign new_n14279_ = ~new_n13689_ & new_n13770_;
  assign new_n14280_ = ~new_n13766_ & new_n14279_;
  assign new_n14281_ = ~new_n13767_ & ~new_n13770_;
  assign new_n14282_ = ~new_n14280_ & ~new_n14281_;
  assign new_n14283_ = \quotient[20]  & ~new_n14282_;
  assign new_n14284_ = ~new_n13679_ & ~new_n13962_;
  assign new_n14285_ = ~new_n13961_ & new_n14284_;
  assign new_n14286_ = ~new_n14283_ & ~new_n14285_;
  assign new_n14287_ = ~\b[8]  & ~new_n14286_;
  assign new_n14288_ = ~new_n13698_ & new_n13765_;
  assign new_n14289_ = ~new_n13761_ & new_n14288_;
  assign new_n14290_ = ~new_n13762_ & ~new_n13765_;
  assign new_n14291_ = ~new_n14289_ & ~new_n14290_;
  assign new_n14292_ = \quotient[20]  & ~new_n14291_;
  assign new_n14293_ = ~new_n13688_ & ~new_n13962_;
  assign new_n14294_ = ~new_n13961_ & new_n14293_;
  assign new_n14295_ = ~new_n14292_ & ~new_n14294_;
  assign new_n14296_ = ~\b[7]  & ~new_n14295_;
  assign new_n14297_ = ~new_n13707_ & new_n13760_;
  assign new_n14298_ = ~new_n13756_ & new_n14297_;
  assign new_n14299_ = ~new_n13757_ & ~new_n13760_;
  assign new_n14300_ = ~new_n14298_ & ~new_n14299_;
  assign new_n14301_ = \quotient[20]  & ~new_n14300_;
  assign new_n14302_ = ~new_n13697_ & ~new_n13962_;
  assign new_n14303_ = ~new_n13961_ & new_n14302_;
  assign new_n14304_ = ~new_n14301_ & ~new_n14303_;
  assign new_n14305_ = ~\b[6]  & ~new_n14304_;
  assign new_n14306_ = ~new_n13716_ & new_n13755_;
  assign new_n14307_ = ~new_n13751_ & new_n14306_;
  assign new_n14308_ = ~new_n13752_ & ~new_n13755_;
  assign new_n14309_ = ~new_n14307_ & ~new_n14308_;
  assign new_n14310_ = \quotient[20]  & ~new_n14309_;
  assign new_n14311_ = ~new_n13706_ & ~new_n13962_;
  assign new_n14312_ = ~new_n13961_ & new_n14311_;
  assign new_n14313_ = ~new_n14310_ & ~new_n14312_;
  assign new_n14314_ = ~\b[5]  & ~new_n14313_;
  assign new_n14315_ = ~new_n13724_ & new_n13750_;
  assign new_n14316_ = ~new_n13746_ & new_n14315_;
  assign new_n14317_ = ~new_n13747_ & ~new_n13750_;
  assign new_n14318_ = ~new_n14316_ & ~new_n14317_;
  assign new_n14319_ = \quotient[20]  & ~new_n14318_;
  assign new_n14320_ = ~new_n13715_ & ~new_n13962_;
  assign new_n14321_ = ~new_n13961_ & new_n14320_;
  assign new_n14322_ = ~new_n14319_ & ~new_n14321_;
  assign new_n14323_ = ~\b[4]  & ~new_n14322_;
  assign new_n14324_ = ~new_n13741_ & new_n13745_;
  assign new_n14325_ = ~new_n13740_ & new_n14324_;
  assign new_n14326_ = ~new_n13742_ & ~new_n13745_;
  assign new_n14327_ = ~new_n14325_ & ~new_n14326_;
  assign new_n14328_ = \quotient[20]  & ~new_n14327_;
  assign new_n14329_ = ~new_n13723_ & ~new_n13962_;
  assign new_n14330_ = ~new_n13961_ & new_n14329_;
  assign new_n14331_ = ~new_n14328_ & ~new_n14330_;
  assign new_n14332_ = ~\b[3]  & ~new_n14331_;
  assign new_n14333_ = ~new_n13737_ & new_n13739_;
  assign new_n14334_ = ~new_n13735_ & new_n14333_;
  assign new_n14335_ = ~new_n13740_ & ~new_n14334_;
  assign new_n14336_ = \quotient[20]  & new_n14335_;
  assign new_n14337_ = ~new_n13734_ & ~new_n13962_;
  assign new_n14338_ = ~new_n13961_ & new_n14337_;
  assign new_n14339_ = ~new_n14336_ & ~new_n14338_;
  assign new_n14340_ = ~\b[2]  & ~new_n14339_;
  assign new_n14341_ = \b[0]  & \quotient[20] ;
  assign new_n14342_ = \a[20]  & ~new_n14341_;
  assign new_n14343_ = new_n13739_ & \quotient[20] ;
  assign new_n14344_ = ~new_n14342_ & ~new_n14343_;
  assign new_n14345_ = \b[1]  & ~new_n14344_;
  assign new_n14346_ = ~\b[1]  & ~new_n14343_;
  assign new_n14347_ = ~new_n14342_ & new_n14346_;
  assign new_n14348_ = ~new_n14345_ & ~new_n14347_;
  assign new_n14349_ = ~\a[19]  & \b[0] ;
  assign new_n14350_ = ~new_n14348_ & ~new_n14349_;
  assign new_n14351_ = ~\b[1]  & ~new_n14344_;
  assign new_n14352_ = ~new_n14350_ & ~new_n14351_;
  assign new_n14353_ = \b[2]  & ~new_n14338_;
  assign new_n14354_ = ~new_n14336_ & new_n14353_;
  assign new_n14355_ = ~new_n14340_ & ~new_n14354_;
  assign new_n14356_ = ~new_n14352_ & new_n14355_;
  assign new_n14357_ = ~new_n14340_ & ~new_n14356_;
  assign new_n14358_ = \b[3]  & ~new_n14330_;
  assign new_n14359_ = ~new_n14328_ & new_n14358_;
  assign new_n14360_ = ~new_n14332_ & ~new_n14359_;
  assign new_n14361_ = ~new_n14357_ & new_n14360_;
  assign new_n14362_ = ~new_n14332_ & ~new_n14361_;
  assign new_n14363_ = \b[4]  & ~new_n14321_;
  assign new_n14364_ = ~new_n14319_ & new_n14363_;
  assign new_n14365_ = ~new_n14323_ & ~new_n14364_;
  assign new_n14366_ = ~new_n14362_ & new_n14365_;
  assign new_n14367_ = ~new_n14323_ & ~new_n14366_;
  assign new_n14368_ = \b[5]  & ~new_n14312_;
  assign new_n14369_ = ~new_n14310_ & new_n14368_;
  assign new_n14370_ = ~new_n14314_ & ~new_n14369_;
  assign new_n14371_ = ~new_n14367_ & new_n14370_;
  assign new_n14372_ = ~new_n14314_ & ~new_n14371_;
  assign new_n14373_ = \b[6]  & ~new_n14303_;
  assign new_n14374_ = ~new_n14301_ & new_n14373_;
  assign new_n14375_ = ~new_n14305_ & ~new_n14374_;
  assign new_n14376_ = ~new_n14372_ & new_n14375_;
  assign new_n14377_ = ~new_n14305_ & ~new_n14376_;
  assign new_n14378_ = \b[7]  & ~new_n14294_;
  assign new_n14379_ = ~new_n14292_ & new_n14378_;
  assign new_n14380_ = ~new_n14296_ & ~new_n14379_;
  assign new_n14381_ = ~new_n14377_ & new_n14380_;
  assign new_n14382_ = ~new_n14296_ & ~new_n14381_;
  assign new_n14383_ = \b[8]  & ~new_n14285_;
  assign new_n14384_ = ~new_n14283_ & new_n14383_;
  assign new_n14385_ = ~new_n14287_ & ~new_n14384_;
  assign new_n14386_ = ~new_n14382_ & new_n14385_;
  assign new_n14387_ = ~new_n14287_ & ~new_n14386_;
  assign new_n14388_ = \b[9]  & ~new_n14276_;
  assign new_n14389_ = ~new_n14274_ & new_n14388_;
  assign new_n14390_ = ~new_n14278_ & ~new_n14389_;
  assign new_n14391_ = ~new_n14387_ & new_n14390_;
  assign new_n14392_ = ~new_n14278_ & ~new_n14391_;
  assign new_n14393_ = \b[10]  & ~new_n14267_;
  assign new_n14394_ = ~new_n14265_ & new_n14393_;
  assign new_n14395_ = ~new_n14269_ & ~new_n14394_;
  assign new_n14396_ = ~new_n14392_ & new_n14395_;
  assign new_n14397_ = ~new_n14269_ & ~new_n14396_;
  assign new_n14398_ = \b[11]  & ~new_n14258_;
  assign new_n14399_ = ~new_n14256_ & new_n14398_;
  assign new_n14400_ = ~new_n14260_ & ~new_n14399_;
  assign new_n14401_ = ~new_n14397_ & new_n14400_;
  assign new_n14402_ = ~new_n14260_ & ~new_n14401_;
  assign new_n14403_ = \b[12]  & ~new_n14249_;
  assign new_n14404_ = ~new_n14247_ & new_n14403_;
  assign new_n14405_ = ~new_n14251_ & ~new_n14404_;
  assign new_n14406_ = ~new_n14402_ & new_n14405_;
  assign new_n14407_ = ~new_n14251_ & ~new_n14406_;
  assign new_n14408_ = \b[13]  & ~new_n14240_;
  assign new_n14409_ = ~new_n14238_ & new_n14408_;
  assign new_n14410_ = ~new_n14242_ & ~new_n14409_;
  assign new_n14411_ = ~new_n14407_ & new_n14410_;
  assign new_n14412_ = ~new_n14242_ & ~new_n14411_;
  assign new_n14413_ = \b[14]  & ~new_n14231_;
  assign new_n14414_ = ~new_n14229_ & new_n14413_;
  assign new_n14415_ = ~new_n14233_ & ~new_n14414_;
  assign new_n14416_ = ~new_n14412_ & new_n14415_;
  assign new_n14417_ = ~new_n14233_ & ~new_n14416_;
  assign new_n14418_ = \b[15]  & ~new_n14222_;
  assign new_n14419_ = ~new_n14220_ & new_n14418_;
  assign new_n14420_ = ~new_n14224_ & ~new_n14419_;
  assign new_n14421_ = ~new_n14417_ & new_n14420_;
  assign new_n14422_ = ~new_n14224_ & ~new_n14421_;
  assign new_n14423_ = \b[16]  & ~new_n14213_;
  assign new_n14424_ = ~new_n14211_ & new_n14423_;
  assign new_n14425_ = ~new_n14215_ & ~new_n14424_;
  assign new_n14426_ = ~new_n14422_ & new_n14425_;
  assign new_n14427_ = ~new_n14215_ & ~new_n14426_;
  assign new_n14428_ = \b[17]  & ~new_n14204_;
  assign new_n14429_ = ~new_n14202_ & new_n14428_;
  assign new_n14430_ = ~new_n14206_ & ~new_n14429_;
  assign new_n14431_ = ~new_n14427_ & new_n14430_;
  assign new_n14432_ = ~new_n14206_ & ~new_n14431_;
  assign new_n14433_ = \b[18]  & ~new_n14195_;
  assign new_n14434_ = ~new_n14193_ & new_n14433_;
  assign new_n14435_ = ~new_n14197_ & ~new_n14434_;
  assign new_n14436_ = ~new_n14432_ & new_n14435_;
  assign new_n14437_ = ~new_n14197_ & ~new_n14436_;
  assign new_n14438_ = \b[19]  & ~new_n14186_;
  assign new_n14439_ = ~new_n14184_ & new_n14438_;
  assign new_n14440_ = ~new_n14188_ & ~new_n14439_;
  assign new_n14441_ = ~new_n14437_ & new_n14440_;
  assign new_n14442_ = ~new_n14188_ & ~new_n14441_;
  assign new_n14443_ = \b[20]  & ~new_n14177_;
  assign new_n14444_ = ~new_n14175_ & new_n14443_;
  assign new_n14445_ = ~new_n14179_ & ~new_n14444_;
  assign new_n14446_ = ~new_n14442_ & new_n14445_;
  assign new_n14447_ = ~new_n14179_ & ~new_n14446_;
  assign new_n14448_ = \b[21]  & ~new_n14168_;
  assign new_n14449_ = ~new_n14166_ & new_n14448_;
  assign new_n14450_ = ~new_n14170_ & ~new_n14449_;
  assign new_n14451_ = ~new_n14447_ & new_n14450_;
  assign new_n14452_ = ~new_n14170_ & ~new_n14451_;
  assign new_n14453_ = \b[22]  & ~new_n14159_;
  assign new_n14454_ = ~new_n14157_ & new_n14453_;
  assign new_n14455_ = ~new_n14161_ & ~new_n14454_;
  assign new_n14456_ = ~new_n14452_ & new_n14455_;
  assign new_n14457_ = ~new_n14161_ & ~new_n14456_;
  assign new_n14458_ = \b[23]  & ~new_n14150_;
  assign new_n14459_ = ~new_n14148_ & new_n14458_;
  assign new_n14460_ = ~new_n14152_ & ~new_n14459_;
  assign new_n14461_ = ~new_n14457_ & new_n14460_;
  assign new_n14462_ = ~new_n14152_ & ~new_n14461_;
  assign new_n14463_ = \b[24]  & ~new_n14141_;
  assign new_n14464_ = ~new_n14139_ & new_n14463_;
  assign new_n14465_ = ~new_n14143_ & ~new_n14464_;
  assign new_n14466_ = ~new_n14462_ & new_n14465_;
  assign new_n14467_ = ~new_n14143_ & ~new_n14466_;
  assign new_n14468_ = \b[25]  & ~new_n14132_;
  assign new_n14469_ = ~new_n14130_ & new_n14468_;
  assign new_n14470_ = ~new_n14134_ & ~new_n14469_;
  assign new_n14471_ = ~new_n14467_ & new_n14470_;
  assign new_n14472_ = ~new_n14134_ & ~new_n14471_;
  assign new_n14473_ = \b[26]  & ~new_n14123_;
  assign new_n14474_ = ~new_n14121_ & new_n14473_;
  assign new_n14475_ = ~new_n14125_ & ~new_n14474_;
  assign new_n14476_ = ~new_n14472_ & new_n14475_;
  assign new_n14477_ = ~new_n14125_ & ~new_n14476_;
  assign new_n14478_ = \b[27]  & ~new_n14114_;
  assign new_n14479_ = ~new_n14112_ & new_n14478_;
  assign new_n14480_ = ~new_n14116_ & ~new_n14479_;
  assign new_n14481_ = ~new_n14477_ & new_n14480_;
  assign new_n14482_ = ~new_n14116_ & ~new_n14481_;
  assign new_n14483_ = \b[28]  & ~new_n14105_;
  assign new_n14484_ = ~new_n14103_ & new_n14483_;
  assign new_n14485_ = ~new_n14107_ & ~new_n14484_;
  assign new_n14486_ = ~new_n14482_ & new_n14485_;
  assign new_n14487_ = ~new_n14107_ & ~new_n14486_;
  assign new_n14488_ = \b[29]  & ~new_n14096_;
  assign new_n14489_ = ~new_n14094_ & new_n14488_;
  assign new_n14490_ = ~new_n14098_ & ~new_n14489_;
  assign new_n14491_ = ~new_n14487_ & new_n14490_;
  assign new_n14492_ = ~new_n14098_ & ~new_n14491_;
  assign new_n14493_ = \b[30]  & ~new_n14087_;
  assign new_n14494_ = ~new_n14085_ & new_n14493_;
  assign new_n14495_ = ~new_n14089_ & ~new_n14494_;
  assign new_n14496_ = ~new_n14492_ & new_n14495_;
  assign new_n14497_ = ~new_n14089_ & ~new_n14496_;
  assign new_n14498_ = \b[31]  & ~new_n14078_;
  assign new_n14499_ = ~new_n14076_ & new_n14498_;
  assign new_n14500_ = ~new_n14080_ & ~new_n14499_;
  assign new_n14501_ = ~new_n14497_ & new_n14500_;
  assign new_n14502_ = ~new_n14080_ & ~new_n14501_;
  assign new_n14503_ = \b[32]  & ~new_n14069_;
  assign new_n14504_ = ~new_n14067_ & new_n14503_;
  assign new_n14505_ = ~new_n14071_ & ~new_n14504_;
  assign new_n14506_ = ~new_n14502_ & new_n14505_;
  assign new_n14507_ = ~new_n14071_ & ~new_n14506_;
  assign new_n14508_ = \b[33]  & ~new_n14060_;
  assign new_n14509_ = ~new_n14058_ & new_n14508_;
  assign new_n14510_ = ~new_n14062_ & ~new_n14509_;
  assign new_n14511_ = ~new_n14507_ & new_n14510_;
  assign new_n14512_ = ~new_n14062_ & ~new_n14511_;
  assign new_n14513_ = \b[34]  & ~new_n14051_;
  assign new_n14514_ = ~new_n14049_ & new_n14513_;
  assign new_n14515_ = ~new_n14053_ & ~new_n14514_;
  assign new_n14516_ = ~new_n14512_ & new_n14515_;
  assign new_n14517_ = ~new_n14053_ & ~new_n14516_;
  assign new_n14518_ = \b[35]  & ~new_n14042_;
  assign new_n14519_ = ~new_n14040_ & new_n14518_;
  assign new_n14520_ = ~new_n14044_ & ~new_n14519_;
  assign new_n14521_ = ~new_n14517_ & new_n14520_;
  assign new_n14522_ = ~new_n14044_ & ~new_n14521_;
  assign new_n14523_ = \b[36]  & ~new_n14033_;
  assign new_n14524_ = ~new_n14031_ & new_n14523_;
  assign new_n14525_ = ~new_n14035_ & ~new_n14524_;
  assign new_n14526_ = ~new_n14522_ & new_n14525_;
  assign new_n14527_ = ~new_n14035_ & ~new_n14526_;
  assign new_n14528_ = \b[37]  & ~new_n14024_;
  assign new_n14529_ = ~new_n14022_ & new_n14528_;
  assign new_n14530_ = ~new_n14026_ & ~new_n14529_;
  assign new_n14531_ = ~new_n14527_ & new_n14530_;
  assign new_n14532_ = ~new_n14026_ & ~new_n14531_;
  assign new_n14533_ = \b[38]  & ~new_n14015_;
  assign new_n14534_ = ~new_n14013_ & new_n14533_;
  assign new_n14535_ = ~new_n14017_ & ~new_n14534_;
  assign new_n14536_ = ~new_n14532_ & new_n14535_;
  assign new_n14537_ = ~new_n14017_ & ~new_n14536_;
  assign new_n14538_ = \b[39]  & ~new_n14006_;
  assign new_n14539_ = ~new_n14004_ & new_n14538_;
  assign new_n14540_ = ~new_n14008_ & ~new_n14539_;
  assign new_n14541_ = ~new_n14537_ & new_n14540_;
  assign new_n14542_ = ~new_n14008_ & ~new_n14541_;
  assign new_n14543_ = \b[40]  & ~new_n13997_;
  assign new_n14544_ = ~new_n13995_ & new_n14543_;
  assign new_n14545_ = ~new_n13999_ & ~new_n14544_;
  assign new_n14546_ = ~new_n14542_ & new_n14545_;
  assign new_n14547_ = ~new_n13999_ & ~new_n14546_;
  assign new_n14548_ = \b[41]  & ~new_n13988_;
  assign new_n14549_ = ~new_n13986_ & new_n14548_;
  assign new_n14550_ = ~new_n13990_ & ~new_n14549_;
  assign new_n14551_ = ~new_n14547_ & new_n14550_;
  assign new_n14552_ = ~new_n13990_ & ~new_n14551_;
  assign new_n14553_ = \b[42]  & ~new_n13979_;
  assign new_n14554_ = ~new_n13977_ & new_n14553_;
  assign new_n14555_ = ~new_n13981_ & ~new_n14554_;
  assign new_n14556_ = ~new_n14552_ & new_n14555_;
  assign new_n14557_ = ~new_n13981_ & ~new_n14556_;
  assign new_n14558_ = \b[43]  & ~new_n13970_;
  assign new_n14559_ = ~new_n13968_ & new_n14558_;
  assign new_n14560_ = ~new_n13972_ & ~new_n14559_;
  assign new_n14561_ = ~new_n14557_ & new_n14560_;
  assign new_n14562_ = ~new_n13972_ & ~new_n14561_;
  assign new_n14563_ = ~new_n13365_ & ~new_n13957_;
  assign new_n14564_ = ~new_n13955_ & new_n14563_;
  assign new_n14565_ = ~new_n13946_ & new_n14564_;
  assign new_n14566_ = ~new_n13955_ & ~new_n13957_;
  assign new_n14567_ = ~new_n13947_ & ~new_n14566_;
  assign new_n14568_ = ~new_n14565_ & ~new_n14567_;
  assign new_n14569_ = \quotient[20]  & ~new_n14568_;
  assign new_n14570_ = ~new_n13954_ & ~new_n13962_;
  assign new_n14571_ = ~new_n13961_ & new_n14570_;
  assign new_n14572_ = ~new_n14569_ & ~new_n14571_;
  assign new_n14573_ = ~\b[44]  & ~new_n14572_;
  assign new_n14574_ = \b[44]  & ~new_n14571_;
  assign new_n14575_ = ~new_n14569_ & new_n14574_;
  assign new_n14576_ = new_n595_ & new_n597_;
  assign new_n14577_ = ~new_n14575_ & new_n14576_;
  assign new_n14578_ = ~new_n14573_ & new_n14577_;
  assign new_n14579_ = ~new_n14562_ & new_n14578_;
  assign new_n14580_ = new_n13958_ & ~new_n14572_;
  assign \quotient[19]  = new_n14579_ | new_n14580_;
  assign new_n14582_ = ~new_n13981_ & new_n14560_;
  assign new_n14583_ = ~new_n14556_ & new_n14582_;
  assign new_n14584_ = ~new_n14557_ & ~new_n14560_;
  assign new_n14585_ = ~new_n14583_ & ~new_n14584_;
  assign new_n14586_ = \quotient[19]  & ~new_n14585_;
  assign new_n14587_ = ~new_n13971_ & ~new_n14580_;
  assign new_n14588_ = ~new_n14579_ & new_n14587_;
  assign new_n14589_ = ~new_n14586_ & ~new_n14588_;
  assign new_n14590_ = ~new_n13972_ & ~new_n14575_;
  assign new_n14591_ = ~new_n14573_ & new_n14590_;
  assign new_n14592_ = ~new_n14561_ & new_n14591_;
  assign new_n14593_ = ~new_n14573_ & ~new_n14575_;
  assign new_n14594_ = ~new_n14562_ & ~new_n14593_;
  assign new_n14595_ = ~new_n14592_ & ~new_n14594_;
  assign new_n14596_ = \quotient[19]  & ~new_n14595_;
  assign new_n14597_ = ~new_n14572_ & ~new_n14580_;
  assign new_n14598_ = ~new_n14579_ & new_n14597_;
  assign new_n14599_ = ~new_n14596_ & ~new_n14598_;
  assign new_n14600_ = ~\b[45]  & ~new_n14599_;
  assign new_n14601_ = ~\b[44]  & ~new_n14589_;
  assign new_n14602_ = ~new_n13990_ & new_n14555_;
  assign new_n14603_ = ~new_n14551_ & new_n14602_;
  assign new_n14604_ = ~new_n14552_ & ~new_n14555_;
  assign new_n14605_ = ~new_n14603_ & ~new_n14604_;
  assign new_n14606_ = \quotient[19]  & ~new_n14605_;
  assign new_n14607_ = ~new_n13980_ & ~new_n14580_;
  assign new_n14608_ = ~new_n14579_ & new_n14607_;
  assign new_n14609_ = ~new_n14606_ & ~new_n14608_;
  assign new_n14610_ = ~\b[43]  & ~new_n14609_;
  assign new_n14611_ = ~new_n13999_ & new_n14550_;
  assign new_n14612_ = ~new_n14546_ & new_n14611_;
  assign new_n14613_ = ~new_n14547_ & ~new_n14550_;
  assign new_n14614_ = ~new_n14612_ & ~new_n14613_;
  assign new_n14615_ = \quotient[19]  & ~new_n14614_;
  assign new_n14616_ = ~new_n13989_ & ~new_n14580_;
  assign new_n14617_ = ~new_n14579_ & new_n14616_;
  assign new_n14618_ = ~new_n14615_ & ~new_n14617_;
  assign new_n14619_ = ~\b[42]  & ~new_n14618_;
  assign new_n14620_ = ~new_n14008_ & new_n14545_;
  assign new_n14621_ = ~new_n14541_ & new_n14620_;
  assign new_n14622_ = ~new_n14542_ & ~new_n14545_;
  assign new_n14623_ = ~new_n14621_ & ~new_n14622_;
  assign new_n14624_ = \quotient[19]  & ~new_n14623_;
  assign new_n14625_ = ~new_n13998_ & ~new_n14580_;
  assign new_n14626_ = ~new_n14579_ & new_n14625_;
  assign new_n14627_ = ~new_n14624_ & ~new_n14626_;
  assign new_n14628_ = ~\b[41]  & ~new_n14627_;
  assign new_n14629_ = ~new_n14017_ & new_n14540_;
  assign new_n14630_ = ~new_n14536_ & new_n14629_;
  assign new_n14631_ = ~new_n14537_ & ~new_n14540_;
  assign new_n14632_ = ~new_n14630_ & ~new_n14631_;
  assign new_n14633_ = \quotient[19]  & ~new_n14632_;
  assign new_n14634_ = ~new_n14007_ & ~new_n14580_;
  assign new_n14635_ = ~new_n14579_ & new_n14634_;
  assign new_n14636_ = ~new_n14633_ & ~new_n14635_;
  assign new_n14637_ = ~\b[40]  & ~new_n14636_;
  assign new_n14638_ = ~new_n14026_ & new_n14535_;
  assign new_n14639_ = ~new_n14531_ & new_n14638_;
  assign new_n14640_ = ~new_n14532_ & ~new_n14535_;
  assign new_n14641_ = ~new_n14639_ & ~new_n14640_;
  assign new_n14642_ = \quotient[19]  & ~new_n14641_;
  assign new_n14643_ = ~new_n14016_ & ~new_n14580_;
  assign new_n14644_ = ~new_n14579_ & new_n14643_;
  assign new_n14645_ = ~new_n14642_ & ~new_n14644_;
  assign new_n14646_ = ~\b[39]  & ~new_n14645_;
  assign new_n14647_ = ~new_n14035_ & new_n14530_;
  assign new_n14648_ = ~new_n14526_ & new_n14647_;
  assign new_n14649_ = ~new_n14527_ & ~new_n14530_;
  assign new_n14650_ = ~new_n14648_ & ~new_n14649_;
  assign new_n14651_ = \quotient[19]  & ~new_n14650_;
  assign new_n14652_ = ~new_n14025_ & ~new_n14580_;
  assign new_n14653_ = ~new_n14579_ & new_n14652_;
  assign new_n14654_ = ~new_n14651_ & ~new_n14653_;
  assign new_n14655_ = ~\b[38]  & ~new_n14654_;
  assign new_n14656_ = ~new_n14044_ & new_n14525_;
  assign new_n14657_ = ~new_n14521_ & new_n14656_;
  assign new_n14658_ = ~new_n14522_ & ~new_n14525_;
  assign new_n14659_ = ~new_n14657_ & ~new_n14658_;
  assign new_n14660_ = \quotient[19]  & ~new_n14659_;
  assign new_n14661_ = ~new_n14034_ & ~new_n14580_;
  assign new_n14662_ = ~new_n14579_ & new_n14661_;
  assign new_n14663_ = ~new_n14660_ & ~new_n14662_;
  assign new_n14664_ = ~\b[37]  & ~new_n14663_;
  assign new_n14665_ = ~new_n14053_ & new_n14520_;
  assign new_n14666_ = ~new_n14516_ & new_n14665_;
  assign new_n14667_ = ~new_n14517_ & ~new_n14520_;
  assign new_n14668_ = ~new_n14666_ & ~new_n14667_;
  assign new_n14669_ = \quotient[19]  & ~new_n14668_;
  assign new_n14670_ = ~new_n14043_ & ~new_n14580_;
  assign new_n14671_ = ~new_n14579_ & new_n14670_;
  assign new_n14672_ = ~new_n14669_ & ~new_n14671_;
  assign new_n14673_ = ~\b[36]  & ~new_n14672_;
  assign new_n14674_ = ~new_n14062_ & new_n14515_;
  assign new_n14675_ = ~new_n14511_ & new_n14674_;
  assign new_n14676_ = ~new_n14512_ & ~new_n14515_;
  assign new_n14677_ = ~new_n14675_ & ~new_n14676_;
  assign new_n14678_ = \quotient[19]  & ~new_n14677_;
  assign new_n14679_ = ~new_n14052_ & ~new_n14580_;
  assign new_n14680_ = ~new_n14579_ & new_n14679_;
  assign new_n14681_ = ~new_n14678_ & ~new_n14680_;
  assign new_n14682_ = ~\b[35]  & ~new_n14681_;
  assign new_n14683_ = ~new_n14071_ & new_n14510_;
  assign new_n14684_ = ~new_n14506_ & new_n14683_;
  assign new_n14685_ = ~new_n14507_ & ~new_n14510_;
  assign new_n14686_ = ~new_n14684_ & ~new_n14685_;
  assign new_n14687_ = \quotient[19]  & ~new_n14686_;
  assign new_n14688_ = ~new_n14061_ & ~new_n14580_;
  assign new_n14689_ = ~new_n14579_ & new_n14688_;
  assign new_n14690_ = ~new_n14687_ & ~new_n14689_;
  assign new_n14691_ = ~\b[34]  & ~new_n14690_;
  assign new_n14692_ = ~new_n14080_ & new_n14505_;
  assign new_n14693_ = ~new_n14501_ & new_n14692_;
  assign new_n14694_ = ~new_n14502_ & ~new_n14505_;
  assign new_n14695_ = ~new_n14693_ & ~new_n14694_;
  assign new_n14696_ = \quotient[19]  & ~new_n14695_;
  assign new_n14697_ = ~new_n14070_ & ~new_n14580_;
  assign new_n14698_ = ~new_n14579_ & new_n14697_;
  assign new_n14699_ = ~new_n14696_ & ~new_n14698_;
  assign new_n14700_ = ~\b[33]  & ~new_n14699_;
  assign new_n14701_ = ~new_n14089_ & new_n14500_;
  assign new_n14702_ = ~new_n14496_ & new_n14701_;
  assign new_n14703_ = ~new_n14497_ & ~new_n14500_;
  assign new_n14704_ = ~new_n14702_ & ~new_n14703_;
  assign new_n14705_ = \quotient[19]  & ~new_n14704_;
  assign new_n14706_ = ~new_n14079_ & ~new_n14580_;
  assign new_n14707_ = ~new_n14579_ & new_n14706_;
  assign new_n14708_ = ~new_n14705_ & ~new_n14707_;
  assign new_n14709_ = ~\b[32]  & ~new_n14708_;
  assign new_n14710_ = ~new_n14098_ & new_n14495_;
  assign new_n14711_ = ~new_n14491_ & new_n14710_;
  assign new_n14712_ = ~new_n14492_ & ~new_n14495_;
  assign new_n14713_ = ~new_n14711_ & ~new_n14712_;
  assign new_n14714_ = \quotient[19]  & ~new_n14713_;
  assign new_n14715_ = ~new_n14088_ & ~new_n14580_;
  assign new_n14716_ = ~new_n14579_ & new_n14715_;
  assign new_n14717_ = ~new_n14714_ & ~new_n14716_;
  assign new_n14718_ = ~\b[31]  & ~new_n14717_;
  assign new_n14719_ = ~new_n14107_ & new_n14490_;
  assign new_n14720_ = ~new_n14486_ & new_n14719_;
  assign new_n14721_ = ~new_n14487_ & ~new_n14490_;
  assign new_n14722_ = ~new_n14720_ & ~new_n14721_;
  assign new_n14723_ = \quotient[19]  & ~new_n14722_;
  assign new_n14724_ = ~new_n14097_ & ~new_n14580_;
  assign new_n14725_ = ~new_n14579_ & new_n14724_;
  assign new_n14726_ = ~new_n14723_ & ~new_n14725_;
  assign new_n14727_ = ~\b[30]  & ~new_n14726_;
  assign new_n14728_ = ~new_n14116_ & new_n14485_;
  assign new_n14729_ = ~new_n14481_ & new_n14728_;
  assign new_n14730_ = ~new_n14482_ & ~new_n14485_;
  assign new_n14731_ = ~new_n14729_ & ~new_n14730_;
  assign new_n14732_ = \quotient[19]  & ~new_n14731_;
  assign new_n14733_ = ~new_n14106_ & ~new_n14580_;
  assign new_n14734_ = ~new_n14579_ & new_n14733_;
  assign new_n14735_ = ~new_n14732_ & ~new_n14734_;
  assign new_n14736_ = ~\b[29]  & ~new_n14735_;
  assign new_n14737_ = ~new_n14125_ & new_n14480_;
  assign new_n14738_ = ~new_n14476_ & new_n14737_;
  assign new_n14739_ = ~new_n14477_ & ~new_n14480_;
  assign new_n14740_ = ~new_n14738_ & ~new_n14739_;
  assign new_n14741_ = \quotient[19]  & ~new_n14740_;
  assign new_n14742_ = ~new_n14115_ & ~new_n14580_;
  assign new_n14743_ = ~new_n14579_ & new_n14742_;
  assign new_n14744_ = ~new_n14741_ & ~new_n14743_;
  assign new_n14745_ = ~\b[28]  & ~new_n14744_;
  assign new_n14746_ = ~new_n14134_ & new_n14475_;
  assign new_n14747_ = ~new_n14471_ & new_n14746_;
  assign new_n14748_ = ~new_n14472_ & ~new_n14475_;
  assign new_n14749_ = ~new_n14747_ & ~new_n14748_;
  assign new_n14750_ = \quotient[19]  & ~new_n14749_;
  assign new_n14751_ = ~new_n14124_ & ~new_n14580_;
  assign new_n14752_ = ~new_n14579_ & new_n14751_;
  assign new_n14753_ = ~new_n14750_ & ~new_n14752_;
  assign new_n14754_ = ~\b[27]  & ~new_n14753_;
  assign new_n14755_ = ~new_n14143_ & new_n14470_;
  assign new_n14756_ = ~new_n14466_ & new_n14755_;
  assign new_n14757_ = ~new_n14467_ & ~new_n14470_;
  assign new_n14758_ = ~new_n14756_ & ~new_n14757_;
  assign new_n14759_ = \quotient[19]  & ~new_n14758_;
  assign new_n14760_ = ~new_n14133_ & ~new_n14580_;
  assign new_n14761_ = ~new_n14579_ & new_n14760_;
  assign new_n14762_ = ~new_n14759_ & ~new_n14761_;
  assign new_n14763_ = ~\b[26]  & ~new_n14762_;
  assign new_n14764_ = ~new_n14152_ & new_n14465_;
  assign new_n14765_ = ~new_n14461_ & new_n14764_;
  assign new_n14766_ = ~new_n14462_ & ~new_n14465_;
  assign new_n14767_ = ~new_n14765_ & ~new_n14766_;
  assign new_n14768_ = \quotient[19]  & ~new_n14767_;
  assign new_n14769_ = ~new_n14142_ & ~new_n14580_;
  assign new_n14770_ = ~new_n14579_ & new_n14769_;
  assign new_n14771_ = ~new_n14768_ & ~new_n14770_;
  assign new_n14772_ = ~\b[25]  & ~new_n14771_;
  assign new_n14773_ = ~new_n14161_ & new_n14460_;
  assign new_n14774_ = ~new_n14456_ & new_n14773_;
  assign new_n14775_ = ~new_n14457_ & ~new_n14460_;
  assign new_n14776_ = ~new_n14774_ & ~new_n14775_;
  assign new_n14777_ = \quotient[19]  & ~new_n14776_;
  assign new_n14778_ = ~new_n14151_ & ~new_n14580_;
  assign new_n14779_ = ~new_n14579_ & new_n14778_;
  assign new_n14780_ = ~new_n14777_ & ~new_n14779_;
  assign new_n14781_ = ~\b[24]  & ~new_n14780_;
  assign new_n14782_ = ~new_n14170_ & new_n14455_;
  assign new_n14783_ = ~new_n14451_ & new_n14782_;
  assign new_n14784_ = ~new_n14452_ & ~new_n14455_;
  assign new_n14785_ = ~new_n14783_ & ~new_n14784_;
  assign new_n14786_ = \quotient[19]  & ~new_n14785_;
  assign new_n14787_ = ~new_n14160_ & ~new_n14580_;
  assign new_n14788_ = ~new_n14579_ & new_n14787_;
  assign new_n14789_ = ~new_n14786_ & ~new_n14788_;
  assign new_n14790_ = ~\b[23]  & ~new_n14789_;
  assign new_n14791_ = ~new_n14179_ & new_n14450_;
  assign new_n14792_ = ~new_n14446_ & new_n14791_;
  assign new_n14793_ = ~new_n14447_ & ~new_n14450_;
  assign new_n14794_ = ~new_n14792_ & ~new_n14793_;
  assign new_n14795_ = \quotient[19]  & ~new_n14794_;
  assign new_n14796_ = ~new_n14169_ & ~new_n14580_;
  assign new_n14797_ = ~new_n14579_ & new_n14796_;
  assign new_n14798_ = ~new_n14795_ & ~new_n14797_;
  assign new_n14799_ = ~\b[22]  & ~new_n14798_;
  assign new_n14800_ = ~new_n14188_ & new_n14445_;
  assign new_n14801_ = ~new_n14441_ & new_n14800_;
  assign new_n14802_ = ~new_n14442_ & ~new_n14445_;
  assign new_n14803_ = ~new_n14801_ & ~new_n14802_;
  assign new_n14804_ = \quotient[19]  & ~new_n14803_;
  assign new_n14805_ = ~new_n14178_ & ~new_n14580_;
  assign new_n14806_ = ~new_n14579_ & new_n14805_;
  assign new_n14807_ = ~new_n14804_ & ~new_n14806_;
  assign new_n14808_ = ~\b[21]  & ~new_n14807_;
  assign new_n14809_ = ~new_n14197_ & new_n14440_;
  assign new_n14810_ = ~new_n14436_ & new_n14809_;
  assign new_n14811_ = ~new_n14437_ & ~new_n14440_;
  assign new_n14812_ = ~new_n14810_ & ~new_n14811_;
  assign new_n14813_ = \quotient[19]  & ~new_n14812_;
  assign new_n14814_ = ~new_n14187_ & ~new_n14580_;
  assign new_n14815_ = ~new_n14579_ & new_n14814_;
  assign new_n14816_ = ~new_n14813_ & ~new_n14815_;
  assign new_n14817_ = ~\b[20]  & ~new_n14816_;
  assign new_n14818_ = ~new_n14206_ & new_n14435_;
  assign new_n14819_ = ~new_n14431_ & new_n14818_;
  assign new_n14820_ = ~new_n14432_ & ~new_n14435_;
  assign new_n14821_ = ~new_n14819_ & ~new_n14820_;
  assign new_n14822_ = \quotient[19]  & ~new_n14821_;
  assign new_n14823_ = ~new_n14196_ & ~new_n14580_;
  assign new_n14824_ = ~new_n14579_ & new_n14823_;
  assign new_n14825_ = ~new_n14822_ & ~new_n14824_;
  assign new_n14826_ = ~\b[19]  & ~new_n14825_;
  assign new_n14827_ = ~new_n14215_ & new_n14430_;
  assign new_n14828_ = ~new_n14426_ & new_n14827_;
  assign new_n14829_ = ~new_n14427_ & ~new_n14430_;
  assign new_n14830_ = ~new_n14828_ & ~new_n14829_;
  assign new_n14831_ = \quotient[19]  & ~new_n14830_;
  assign new_n14832_ = ~new_n14205_ & ~new_n14580_;
  assign new_n14833_ = ~new_n14579_ & new_n14832_;
  assign new_n14834_ = ~new_n14831_ & ~new_n14833_;
  assign new_n14835_ = ~\b[18]  & ~new_n14834_;
  assign new_n14836_ = ~new_n14224_ & new_n14425_;
  assign new_n14837_ = ~new_n14421_ & new_n14836_;
  assign new_n14838_ = ~new_n14422_ & ~new_n14425_;
  assign new_n14839_ = ~new_n14837_ & ~new_n14838_;
  assign new_n14840_ = \quotient[19]  & ~new_n14839_;
  assign new_n14841_ = ~new_n14214_ & ~new_n14580_;
  assign new_n14842_ = ~new_n14579_ & new_n14841_;
  assign new_n14843_ = ~new_n14840_ & ~new_n14842_;
  assign new_n14844_ = ~\b[17]  & ~new_n14843_;
  assign new_n14845_ = ~new_n14233_ & new_n14420_;
  assign new_n14846_ = ~new_n14416_ & new_n14845_;
  assign new_n14847_ = ~new_n14417_ & ~new_n14420_;
  assign new_n14848_ = ~new_n14846_ & ~new_n14847_;
  assign new_n14849_ = \quotient[19]  & ~new_n14848_;
  assign new_n14850_ = ~new_n14223_ & ~new_n14580_;
  assign new_n14851_ = ~new_n14579_ & new_n14850_;
  assign new_n14852_ = ~new_n14849_ & ~new_n14851_;
  assign new_n14853_ = ~\b[16]  & ~new_n14852_;
  assign new_n14854_ = ~new_n14242_ & new_n14415_;
  assign new_n14855_ = ~new_n14411_ & new_n14854_;
  assign new_n14856_ = ~new_n14412_ & ~new_n14415_;
  assign new_n14857_ = ~new_n14855_ & ~new_n14856_;
  assign new_n14858_ = \quotient[19]  & ~new_n14857_;
  assign new_n14859_ = ~new_n14232_ & ~new_n14580_;
  assign new_n14860_ = ~new_n14579_ & new_n14859_;
  assign new_n14861_ = ~new_n14858_ & ~new_n14860_;
  assign new_n14862_ = ~\b[15]  & ~new_n14861_;
  assign new_n14863_ = ~new_n14251_ & new_n14410_;
  assign new_n14864_ = ~new_n14406_ & new_n14863_;
  assign new_n14865_ = ~new_n14407_ & ~new_n14410_;
  assign new_n14866_ = ~new_n14864_ & ~new_n14865_;
  assign new_n14867_ = \quotient[19]  & ~new_n14866_;
  assign new_n14868_ = ~new_n14241_ & ~new_n14580_;
  assign new_n14869_ = ~new_n14579_ & new_n14868_;
  assign new_n14870_ = ~new_n14867_ & ~new_n14869_;
  assign new_n14871_ = ~\b[14]  & ~new_n14870_;
  assign new_n14872_ = ~new_n14260_ & new_n14405_;
  assign new_n14873_ = ~new_n14401_ & new_n14872_;
  assign new_n14874_ = ~new_n14402_ & ~new_n14405_;
  assign new_n14875_ = ~new_n14873_ & ~new_n14874_;
  assign new_n14876_ = \quotient[19]  & ~new_n14875_;
  assign new_n14877_ = ~new_n14250_ & ~new_n14580_;
  assign new_n14878_ = ~new_n14579_ & new_n14877_;
  assign new_n14879_ = ~new_n14876_ & ~new_n14878_;
  assign new_n14880_ = ~\b[13]  & ~new_n14879_;
  assign new_n14881_ = ~new_n14269_ & new_n14400_;
  assign new_n14882_ = ~new_n14396_ & new_n14881_;
  assign new_n14883_ = ~new_n14397_ & ~new_n14400_;
  assign new_n14884_ = ~new_n14882_ & ~new_n14883_;
  assign new_n14885_ = \quotient[19]  & ~new_n14884_;
  assign new_n14886_ = ~new_n14259_ & ~new_n14580_;
  assign new_n14887_ = ~new_n14579_ & new_n14886_;
  assign new_n14888_ = ~new_n14885_ & ~new_n14887_;
  assign new_n14889_ = ~\b[12]  & ~new_n14888_;
  assign new_n14890_ = ~new_n14278_ & new_n14395_;
  assign new_n14891_ = ~new_n14391_ & new_n14890_;
  assign new_n14892_ = ~new_n14392_ & ~new_n14395_;
  assign new_n14893_ = ~new_n14891_ & ~new_n14892_;
  assign new_n14894_ = \quotient[19]  & ~new_n14893_;
  assign new_n14895_ = ~new_n14268_ & ~new_n14580_;
  assign new_n14896_ = ~new_n14579_ & new_n14895_;
  assign new_n14897_ = ~new_n14894_ & ~new_n14896_;
  assign new_n14898_ = ~\b[11]  & ~new_n14897_;
  assign new_n14899_ = ~new_n14287_ & new_n14390_;
  assign new_n14900_ = ~new_n14386_ & new_n14899_;
  assign new_n14901_ = ~new_n14387_ & ~new_n14390_;
  assign new_n14902_ = ~new_n14900_ & ~new_n14901_;
  assign new_n14903_ = \quotient[19]  & ~new_n14902_;
  assign new_n14904_ = ~new_n14277_ & ~new_n14580_;
  assign new_n14905_ = ~new_n14579_ & new_n14904_;
  assign new_n14906_ = ~new_n14903_ & ~new_n14905_;
  assign new_n14907_ = ~\b[10]  & ~new_n14906_;
  assign new_n14908_ = ~new_n14296_ & new_n14385_;
  assign new_n14909_ = ~new_n14381_ & new_n14908_;
  assign new_n14910_ = ~new_n14382_ & ~new_n14385_;
  assign new_n14911_ = ~new_n14909_ & ~new_n14910_;
  assign new_n14912_ = \quotient[19]  & ~new_n14911_;
  assign new_n14913_ = ~new_n14286_ & ~new_n14580_;
  assign new_n14914_ = ~new_n14579_ & new_n14913_;
  assign new_n14915_ = ~new_n14912_ & ~new_n14914_;
  assign new_n14916_ = ~\b[9]  & ~new_n14915_;
  assign new_n14917_ = ~new_n14305_ & new_n14380_;
  assign new_n14918_ = ~new_n14376_ & new_n14917_;
  assign new_n14919_ = ~new_n14377_ & ~new_n14380_;
  assign new_n14920_ = ~new_n14918_ & ~new_n14919_;
  assign new_n14921_ = \quotient[19]  & ~new_n14920_;
  assign new_n14922_ = ~new_n14295_ & ~new_n14580_;
  assign new_n14923_ = ~new_n14579_ & new_n14922_;
  assign new_n14924_ = ~new_n14921_ & ~new_n14923_;
  assign new_n14925_ = ~\b[8]  & ~new_n14924_;
  assign new_n14926_ = ~new_n14314_ & new_n14375_;
  assign new_n14927_ = ~new_n14371_ & new_n14926_;
  assign new_n14928_ = ~new_n14372_ & ~new_n14375_;
  assign new_n14929_ = ~new_n14927_ & ~new_n14928_;
  assign new_n14930_ = \quotient[19]  & ~new_n14929_;
  assign new_n14931_ = ~new_n14304_ & ~new_n14580_;
  assign new_n14932_ = ~new_n14579_ & new_n14931_;
  assign new_n14933_ = ~new_n14930_ & ~new_n14932_;
  assign new_n14934_ = ~\b[7]  & ~new_n14933_;
  assign new_n14935_ = ~new_n14323_ & new_n14370_;
  assign new_n14936_ = ~new_n14366_ & new_n14935_;
  assign new_n14937_ = ~new_n14367_ & ~new_n14370_;
  assign new_n14938_ = ~new_n14936_ & ~new_n14937_;
  assign new_n14939_ = \quotient[19]  & ~new_n14938_;
  assign new_n14940_ = ~new_n14313_ & ~new_n14580_;
  assign new_n14941_ = ~new_n14579_ & new_n14940_;
  assign new_n14942_ = ~new_n14939_ & ~new_n14941_;
  assign new_n14943_ = ~\b[6]  & ~new_n14942_;
  assign new_n14944_ = ~new_n14332_ & new_n14365_;
  assign new_n14945_ = ~new_n14361_ & new_n14944_;
  assign new_n14946_ = ~new_n14362_ & ~new_n14365_;
  assign new_n14947_ = ~new_n14945_ & ~new_n14946_;
  assign new_n14948_ = \quotient[19]  & ~new_n14947_;
  assign new_n14949_ = ~new_n14322_ & ~new_n14580_;
  assign new_n14950_ = ~new_n14579_ & new_n14949_;
  assign new_n14951_ = ~new_n14948_ & ~new_n14950_;
  assign new_n14952_ = ~\b[5]  & ~new_n14951_;
  assign new_n14953_ = ~new_n14340_ & new_n14360_;
  assign new_n14954_ = ~new_n14356_ & new_n14953_;
  assign new_n14955_ = ~new_n14357_ & ~new_n14360_;
  assign new_n14956_ = ~new_n14954_ & ~new_n14955_;
  assign new_n14957_ = \quotient[19]  & ~new_n14956_;
  assign new_n14958_ = ~new_n14331_ & ~new_n14580_;
  assign new_n14959_ = ~new_n14579_ & new_n14958_;
  assign new_n14960_ = ~new_n14957_ & ~new_n14959_;
  assign new_n14961_ = ~\b[4]  & ~new_n14960_;
  assign new_n14962_ = ~new_n14351_ & new_n14355_;
  assign new_n14963_ = ~new_n14350_ & new_n14962_;
  assign new_n14964_ = ~new_n14352_ & ~new_n14355_;
  assign new_n14965_ = ~new_n14963_ & ~new_n14964_;
  assign new_n14966_ = \quotient[19]  & ~new_n14965_;
  assign new_n14967_ = ~new_n14339_ & ~new_n14580_;
  assign new_n14968_ = ~new_n14579_ & new_n14967_;
  assign new_n14969_ = ~new_n14966_ & ~new_n14968_;
  assign new_n14970_ = ~\b[3]  & ~new_n14969_;
  assign new_n14971_ = ~new_n14347_ & new_n14349_;
  assign new_n14972_ = ~new_n14345_ & new_n14971_;
  assign new_n14973_ = ~new_n14350_ & ~new_n14972_;
  assign new_n14974_ = \quotient[19]  & new_n14973_;
  assign new_n14975_ = ~new_n14344_ & ~new_n14580_;
  assign new_n14976_ = ~new_n14579_ & new_n14975_;
  assign new_n14977_ = ~new_n14974_ & ~new_n14976_;
  assign new_n14978_ = ~\b[2]  & ~new_n14977_;
  assign new_n14979_ = \b[0]  & \quotient[19] ;
  assign new_n14980_ = \a[19]  & ~new_n14979_;
  assign new_n14981_ = new_n14349_ & \quotient[19] ;
  assign new_n14982_ = ~new_n14980_ & ~new_n14981_;
  assign new_n14983_ = \b[1]  & ~new_n14982_;
  assign new_n14984_ = ~\b[1]  & ~new_n14981_;
  assign new_n14985_ = ~new_n14980_ & new_n14984_;
  assign new_n14986_ = ~new_n14983_ & ~new_n14985_;
  assign new_n14987_ = ~\a[18]  & \b[0] ;
  assign new_n14988_ = ~new_n14986_ & ~new_n14987_;
  assign new_n14989_ = ~\b[1]  & ~new_n14982_;
  assign new_n14990_ = ~new_n14988_ & ~new_n14989_;
  assign new_n14991_ = \b[2]  & ~new_n14976_;
  assign new_n14992_ = ~new_n14974_ & new_n14991_;
  assign new_n14993_ = ~new_n14978_ & ~new_n14992_;
  assign new_n14994_ = ~new_n14990_ & new_n14993_;
  assign new_n14995_ = ~new_n14978_ & ~new_n14994_;
  assign new_n14996_ = \b[3]  & ~new_n14968_;
  assign new_n14997_ = ~new_n14966_ & new_n14996_;
  assign new_n14998_ = ~new_n14970_ & ~new_n14997_;
  assign new_n14999_ = ~new_n14995_ & new_n14998_;
  assign new_n15000_ = ~new_n14970_ & ~new_n14999_;
  assign new_n15001_ = \b[4]  & ~new_n14959_;
  assign new_n15002_ = ~new_n14957_ & new_n15001_;
  assign new_n15003_ = ~new_n14961_ & ~new_n15002_;
  assign new_n15004_ = ~new_n15000_ & new_n15003_;
  assign new_n15005_ = ~new_n14961_ & ~new_n15004_;
  assign new_n15006_ = \b[5]  & ~new_n14950_;
  assign new_n15007_ = ~new_n14948_ & new_n15006_;
  assign new_n15008_ = ~new_n14952_ & ~new_n15007_;
  assign new_n15009_ = ~new_n15005_ & new_n15008_;
  assign new_n15010_ = ~new_n14952_ & ~new_n15009_;
  assign new_n15011_ = \b[6]  & ~new_n14941_;
  assign new_n15012_ = ~new_n14939_ & new_n15011_;
  assign new_n15013_ = ~new_n14943_ & ~new_n15012_;
  assign new_n15014_ = ~new_n15010_ & new_n15013_;
  assign new_n15015_ = ~new_n14943_ & ~new_n15014_;
  assign new_n15016_ = \b[7]  & ~new_n14932_;
  assign new_n15017_ = ~new_n14930_ & new_n15016_;
  assign new_n15018_ = ~new_n14934_ & ~new_n15017_;
  assign new_n15019_ = ~new_n15015_ & new_n15018_;
  assign new_n15020_ = ~new_n14934_ & ~new_n15019_;
  assign new_n15021_ = \b[8]  & ~new_n14923_;
  assign new_n15022_ = ~new_n14921_ & new_n15021_;
  assign new_n15023_ = ~new_n14925_ & ~new_n15022_;
  assign new_n15024_ = ~new_n15020_ & new_n15023_;
  assign new_n15025_ = ~new_n14925_ & ~new_n15024_;
  assign new_n15026_ = \b[9]  & ~new_n14914_;
  assign new_n15027_ = ~new_n14912_ & new_n15026_;
  assign new_n15028_ = ~new_n14916_ & ~new_n15027_;
  assign new_n15029_ = ~new_n15025_ & new_n15028_;
  assign new_n15030_ = ~new_n14916_ & ~new_n15029_;
  assign new_n15031_ = \b[10]  & ~new_n14905_;
  assign new_n15032_ = ~new_n14903_ & new_n15031_;
  assign new_n15033_ = ~new_n14907_ & ~new_n15032_;
  assign new_n15034_ = ~new_n15030_ & new_n15033_;
  assign new_n15035_ = ~new_n14907_ & ~new_n15034_;
  assign new_n15036_ = \b[11]  & ~new_n14896_;
  assign new_n15037_ = ~new_n14894_ & new_n15036_;
  assign new_n15038_ = ~new_n14898_ & ~new_n15037_;
  assign new_n15039_ = ~new_n15035_ & new_n15038_;
  assign new_n15040_ = ~new_n14898_ & ~new_n15039_;
  assign new_n15041_ = \b[12]  & ~new_n14887_;
  assign new_n15042_ = ~new_n14885_ & new_n15041_;
  assign new_n15043_ = ~new_n14889_ & ~new_n15042_;
  assign new_n15044_ = ~new_n15040_ & new_n15043_;
  assign new_n15045_ = ~new_n14889_ & ~new_n15044_;
  assign new_n15046_ = \b[13]  & ~new_n14878_;
  assign new_n15047_ = ~new_n14876_ & new_n15046_;
  assign new_n15048_ = ~new_n14880_ & ~new_n15047_;
  assign new_n15049_ = ~new_n15045_ & new_n15048_;
  assign new_n15050_ = ~new_n14880_ & ~new_n15049_;
  assign new_n15051_ = \b[14]  & ~new_n14869_;
  assign new_n15052_ = ~new_n14867_ & new_n15051_;
  assign new_n15053_ = ~new_n14871_ & ~new_n15052_;
  assign new_n15054_ = ~new_n15050_ & new_n15053_;
  assign new_n15055_ = ~new_n14871_ & ~new_n15054_;
  assign new_n15056_ = \b[15]  & ~new_n14860_;
  assign new_n15057_ = ~new_n14858_ & new_n15056_;
  assign new_n15058_ = ~new_n14862_ & ~new_n15057_;
  assign new_n15059_ = ~new_n15055_ & new_n15058_;
  assign new_n15060_ = ~new_n14862_ & ~new_n15059_;
  assign new_n15061_ = \b[16]  & ~new_n14851_;
  assign new_n15062_ = ~new_n14849_ & new_n15061_;
  assign new_n15063_ = ~new_n14853_ & ~new_n15062_;
  assign new_n15064_ = ~new_n15060_ & new_n15063_;
  assign new_n15065_ = ~new_n14853_ & ~new_n15064_;
  assign new_n15066_ = \b[17]  & ~new_n14842_;
  assign new_n15067_ = ~new_n14840_ & new_n15066_;
  assign new_n15068_ = ~new_n14844_ & ~new_n15067_;
  assign new_n15069_ = ~new_n15065_ & new_n15068_;
  assign new_n15070_ = ~new_n14844_ & ~new_n15069_;
  assign new_n15071_ = \b[18]  & ~new_n14833_;
  assign new_n15072_ = ~new_n14831_ & new_n15071_;
  assign new_n15073_ = ~new_n14835_ & ~new_n15072_;
  assign new_n15074_ = ~new_n15070_ & new_n15073_;
  assign new_n15075_ = ~new_n14835_ & ~new_n15074_;
  assign new_n15076_ = \b[19]  & ~new_n14824_;
  assign new_n15077_ = ~new_n14822_ & new_n15076_;
  assign new_n15078_ = ~new_n14826_ & ~new_n15077_;
  assign new_n15079_ = ~new_n15075_ & new_n15078_;
  assign new_n15080_ = ~new_n14826_ & ~new_n15079_;
  assign new_n15081_ = \b[20]  & ~new_n14815_;
  assign new_n15082_ = ~new_n14813_ & new_n15081_;
  assign new_n15083_ = ~new_n14817_ & ~new_n15082_;
  assign new_n15084_ = ~new_n15080_ & new_n15083_;
  assign new_n15085_ = ~new_n14817_ & ~new_n15084_;
  assign new_n15086_ = \b[21]  & ~new_n14806_;
  assign new_n15087_ = ~new_n14804_ & new_n15086_;
  assign new_n15088_ = ~new_n14808_ & ~new_n15087_;
  assign new_n15089_ = ~new_n15085_ & new_n15088_;
  assign new_n15090_ = ~new_n14808_ & ~new_n15089_;
  assign new_n15091_ = \b[22]  & ~new_n14797_;
  assign new_n15092_ = ~new_n14795_ & new_n15091_;
  assign new_n15093_ = ~new_n14799_ & ~new_n15092_;
  assign new_n15094_ = ~new_n15090_ & new_n15093_;
  assign new_n15095_ = ~new_n14799_ & ~new_n15094_;
  assign new_n15096_ = \b[23]  & ~new_n14788_;
  assign new_n15097_ = ~new_n14786_ & new_n15096_;
  assign new_n15098_ = ~new_n14790_ & ~new_n15097_;
  assign new_n15099_ = ~new_n15095_ & new_n15098_;
  assign new_n15100_ = ~new_n14790_ & ~new_n15099_;
  assign new_n15101_ = \b[24]  & ~new_n14779_;
  assign new_n15102_ = ~new_n14777_ & new_n15101_;
  assign new_n15103_ = ~new_n14781_ & ~new_n15102_;
  assign new_n15104_ = ~new_n15100_ & new_n15103_;
  assign new_n15105_ = ~new_n14781_ & ~new_n15104_;
  assign new_n15106_ = \b[25]  & ~new_n14770_;
  assign new_n15107_ = ~new_n14768_ & new_n15106_;
  assign new_n15108_ = ~new_n14772_ & ~new_n15107_;
  assign new_n15109_ = ~new_n15105_ & new_n15108_;
  assign new_n15110_ = ~new_n14772_ & ~new_n15109_;
  assign new_n15111_ = \b[26]  & ~new_n14761_;
  assign new_n15112_ = ~new_n14759_ & new_n15111_;
  assign new_n15113_ = ~new_n14763_ & ~new_n15112_;
  assign new_n15114_ = ~new_n15110_ & new_n15113_;
  assign new_n15115_ = ~new_n14763_ & ~new_n15114_;
  assign new_n15116_ = \b[27]  & ~new_n14752_;
  assign new_n15117_ = ~new_n14750_ & new_n15116_;
  assign new_n15118_ = ~new_n14754_ & ~new_n15117_;
  assign new_n15119_ = ~new_n15115_ & new_n15118_;
  assign new_n15120_ = ~new_n14754_ & ~new_n15119_;
  assign new_n15121_ = \b[28]  & ~new_n14743_;
  assign new_n15122_ = ~new_n14741_ & new_n15121_;
  assign new_n15123_ = ~new_n14745_ & ~new_n15122_;
  assign new_n15124_ = ~new_n15120_ & new_n15123_;
  assign new_n15125_ = ~new_n14745_ & ~new_n15124_;
  assign new_n15126_ = \b[29]  & ~new_n14734_;
  assign new_n15127_ = ~new_n14732_ & new_n15126_;
  assign new_n15128_ = ~new_n14736_ & ~new_n15127_;
  assign new_n15129_ = ~new_n15125_ & new_n15128_;
  assign new_n15130_ = ~new_n14736_ & ~new_n15129_;
  assign new_n15131_ = \b[30]  & ~new_n14725_;
  assign new_n15132_ = ~new_n14723_ & new_n15131_;
  assign new_n15133_ = ~new_n14727_ & ~new_n15132_;
  assign new_n15134_ = ~new_n15130_ & new_n15133_;
  assign new_n15135_ = ~new_n14727_ & ~new_n15134_;
  assign new_n15136_ = \b[31]  & ~new_n14716_;
  assign new_n15137_ = ~new_n14714_ & new_n15136_;
  assign new_n15138_ = ~new_n14718_ & ~new_n15137_;
  assign new_n15139_ = ~new_n15135_ & new_n15138_;
  assign new_n15140_ = ~new_n14718_ & ~new_n15139_;
  assign new_n15141_ = \b[32]  & ~new_n14707_;
  assign new_n15142_ = ~new_n14705_ & new_n15141_;
  assign new_n15143_ = ~new_n14709_ & ~new_n15142_;
  assign new_n15144_ = ~new_n15140_ & new_n15143_;
  assign new_n15145_ = ~new_n14709_ & ~new_n15144_;
  assign new_n15146_ = \b[33]  & ~new_n14698_;
  assign new_n15147_ = ~new_n14696_ & new_n15146_;
  assign new_n15148_ = ~new_n14700_ & ~new_n15147_;
  assign new_n15149_ = ~new_n15145_ & new_n15148_;
  assign new_n15150_ = ~new_n14700_ & ~new_n15149_;
  assign new_n15151_ = \b[34]  & ~new_n14689_;
  assign new_n15152_ = ~new_n14687_ & new_n15151_;
  assign new_n15153_ = ~new_n14691_ & ~new_n15152_;
  assign new_n15154_ = ~new_n15150_ & new_n15153_;
  assign new_n15155_ = ~new_n14691_ & ~new_n15154_;
  assign new_n15156_ = \b[35]  & ~new_n14680_;
  assign new_n15157_ = ~new_n14678_ & new_n15156_;
  assign new_n15158_ = ~new_n14682_ & ~new_n15157_;
  assign new_n15159_ = ~new_n15155_ & new_n15158_;
  assign new_n15160_ = ~new_n14682_ & ~new_n15159_;
  assign new_n15161_ = \b[36]  & ~new_n14671_;
  assign new_n15162_ = ~new_n14669_ & new_n15161_;
  assign new_n15163_ = ~new_n14673_ & ~new_n15162_;
  assign new_n15164_ = ~new_n15160_ & new_n15163_;
  assign new_n15165_ = ~new_n14673_ & ~new_n15164_;
  assign new_n15166_ = \b[37]  & ~new_n14662_;
  assign new_n15167_ = ~new_n14660_ & new_n15166_;
  assign new_n15168_ = ~new_n14664_ & ~new_n15167_;
  assign new_n15169_ = ~new_n15165_ & new_n15168_;
  assign new_n15170_ = ~new_n14664_ & ~new_n15169_;
  assign new_n15171_ = \b[38]  & ~new_n14653_;
  assign new_n15172_ = ~new_n14651_ & new_n15171_;
  assign new_n15173_ = ~new_n14655_ & ~new_n15172_;
  assign new_n15174_ = ~new_n15170_ & new_n15173_;
  assign new_n15175_ = ~new_n14655_ & ~new_n15174_;
  assign new_n15176_ = \b[39]  & ~new_n14644_;
  assign new_n15177_ = ~new_n14642_ & new_n15176_;
  assign new_n15178_ = ~new_n14646_ & ~new_n15177_;
  assign new_n15179_ = ~new_n15175_ & new_n15178_;
  assign new_n15180_ = ~new_n14646_ & ~new_n15179_;
  assign new_n15181_ = \b[40]  & ~new_n14635_;
  assign new_n15182_ = ~new_n14633_ & new_n15181_;
  assign new_n15183_ = ~new_n14637_ & ~new_n15182_;
  assign new_n15184_ = ~new_n15180_ & new_n15183_;
  assign new_n15185_ = ~new_n14637_ & ~new_n15184_;
  assign new_n15186_ = \b[41]  & ~new_n14626_;
  assign new_n15187_ = ~new_n14624_ & new_n15186_;
  assign new_n15188_ = ~new_n14628_ & ~new_n15187_;
  assign new_n15189_ = ~new_n15185_ & new_n15188_;
  assign new_n15190_ = ~new_n14628_ & ~new_n15189_;
  assign new_n15191_ = \b[42]  & ~new_n14617_;
  assign new_n15192_ = ~new_n14615_ & new_n15191_;
  assign new_n15193_ = ~new_n14619_ & ~new_n15192_;
  assign new_n15194_ = ~new_n15190_ & new_n15193_;
  assign new_n15195_ = ~new_n14619_ & ~new_n15194_;
  assign new_n15196_ = \b[43]  & ~new_n14608_;
  assign new_n15197_ = ~new_n14606_ & new_n15196_;
  assign new_n15198_ = ~new_n14610_ & ~new_n15197_;
  assign new_n15199_ = ~new_n15195_ & new_n15198_;
  assign new_n15200_ = ~new_n14610_ & ~new_n15199_;
  assign new_n15201_ = \b[44]  & ~new_n14588_;
  assign new_n15202_ = ~new_n14586_ & new_n15201_;
  assign new_n15203_ = ~new_n14601_ & ~new_n15202_;
  assign new_n15204_ = ~new_n15200_ & new_n15203_;
  assign new_n15205_ = ~new_n14601_ & ~new_n15204_;
  assign new_n15206_ = \b[45]  & ~new_n14598_;
  assign new_n15207_ = ~new_n14596_ & new_n15206_;
  assign new_n15208_ = ~new_n14600_ & ~new_n15207_;
  assign new_n15209_ = ~new_n15205_ & new_n15208_;
  assign new_n15210_ = ~new_n14600_ & ~new_n15209_;
  assign new_n15211_ = new_n298_ & new_n300_;
  assign new_n15212_ = new_n288_ & new_n15211_;
  assign \quotient[18]  = ~new_n15210_ & new_n15212_;
  assign new_n15214_ = ~new_n14589_ & ~\quotient[18] ;
  assign new_n15215_ = ~new_n14610_ & new_n15203_;
  assign new_n15216_ = ~new_n15199_ & new_n15215_;
  assign new_n15217_ = ~new_n15200_ & ~new_n15203_;
  assign new_n15218_ = ~new_n15216_ & ~new_n15217_;
  assign new_n15219_ = new_n15212_ & ~new_n15218_;
  assign new_n15220_ = ~new_n15210_ & new_n15219_;
  assign new_n15221_ = ~new_n15214_ & ~new_n15220_;
  assign new_n15222_ = ~\b[45]  & ~new_n15221_;
  assign new_n15223_ = ~new_n14609_ & ~\quotient[18] ;
  assign new_n15224_ = ~new_n14619_ & new_n15198_;
  assign new_n15225_ = ~new_n15194_ & new_n15224_;
  assign new_n15226_ = ~new_n15195_ & ~new_n15198_;
  assign new_n15227_ = ~new_n15225_ & ~new_n15226_;
  assign new_n15228_ = new_n15212_ & ~new_n15227_;
  assign new_n15229_ = ~new_n15210_ & new_n15228_;
  assign new_n15230_ = ~new_n15223_ & ~new_n15229_;
  assign new_n15231_ = ~\b[44]  & ~new_n15230_;
  assign new_n15232_ = ~new_n14618_ & ~\quotient[18] ;
  assign new_n15233_ = ~new_n14628_ & new_n15193_;
  assign new_n15234_ = ~new_n15189_ & new_n15233_;
  assign new_n15235_ = ~new_n15190_ & ~new_n15193_;
  assign new_n15236_ = ~new_n15234_ & ~new_n15235_;
  assign new_n15237_ = new_n15212_ & ~new_n15236_;
  assign new_n15238_ = ~new_n15210_ & new_n15237_;
  assign new_n15239_ = ~new_n15232_ & ~new_n15238_;
  assign new_n15240_ = ~\b[43]  & ~new_n15239_;
  assign new_n15241_ = ~new_n14627_ & ~\quotient[18] ;
  assign new_n15242_ = ~new_n14637_ & new_n15188_;
  assign new_n15243_ = ~new_n15184_ & new_n15242_;
  assign new_n15244_ = ~new_n15185_ & ~new_n15188_;
  assign new_n15245_ = ~new_n15243_ & ~new_n15244_;
  assign new_n15246_ = new_n15212_ & ~new_n15245_;
  assign new_n15247_ = ~new_n15210_ & new_n15246_;
  assign new_n15248_ = ~new_n15241_ & ~new_n15247_;
  assign new_n15249_ = ~\b[42]  & ~new_n15248_;
  assign new_n15250_ = ~new_n14636_ & ~\quotient[18] ;
  assign new_n15251_ = ~new_n14646_ & new_n15183_;
  assign new_n15252_ = ~new_n15179_ & new_n15251_;
  assign new_n15253_ = ~new_n15180_ & ~new_n15183_;
  assign new_n15254_ = ~new_n15252_ & ~new_n15253_;
  assign new_n15255_ = new_n15212_ & ~new_n15254_;
  assign new_n15256_ = ~new_n15210_ & new_n15255_;
  assign new_n15257_ = ~new_n15250_ & ~new_n15256_;
  assign new_n15258_ = ~\b[41]  & ~new_n15257_;
  assign new_n15259_ = ~new_n14645_ & ~\quotient[18] ;
  assign new_n15260_ = ~new_n14655_ & new_n15178_;
  assign new_n15261_ = ~new_n15174_ & new_n15260_;
  assign new_n15262_ = ~new_n15175_ & ~new_n15178_;
  assign new_n15263_ = ~new_n15261_ & ~new_n15262_;
  assign new_n15264_ = new_n15212_ & ~new_n15263_;
  assign new_n15265_ = ~new_n15210_ & new_n15264_;
  assign new_n15266_ = ~new_n15259_ & ~new_n15265_;
  assign new_n15267_ = ~\b[40]  & ~new_n15266_;
  assign new_n15268_ = ~new_n14654_ & ~\quotient[18] ;
  assign new_n15269_ = ~new_n14664_ & new_n15173_;
  assign new_n15270_ = ~new_n15169_ & new_n15269_;
  assign new_n15271_ = ~new_n15170_ & ~new_n15173_;
  assign new_n15272_ = ~new_n15270_ & ~new_n15271_;
  assign new_n15273_ = new_n15212_ & ~new_n15272_;
  assign new_n15274_ = ~new_n15210_ & new_n15273_;
  assign new_n15275_ = ~new_n15268_ & ~new_n15274_;
  assign new_n15276_ = ~\b[39]  & ~new_n15275_;
  assign new_n15277_ = ~new_n14663_ & ~\quotient[18] ;
  assign new_n15278_ = ~new_n14673_ & new_n15168_;
  assign new_n15279_ = ~new_n15164_ & new_n15278_;
  assign new_n15280_ = ~new_n15165_ & ~new_n15168_;
  assign new_n15281_ = ~new_n15279_ & ~new_n15280_;
  assign new_n15282_ = new_n15212_ & ~new_n15281_;
  assign new_n15283_ = ~new_n15210_ & new_n15282_;
  assign new_n15284_ = ~new_n15277_ & ~new_n15283_;
  assign new_n15285_ = ~\b[38]  & ~new_n15284_;
  assign new_n15286_ = ~new_n14672_ & ~\quotient[18] ;
  assign new_n15287_ = ~new_n14682_ & new_n15163_;
  assign new_n15288_ = ~new_n15159_ & new_n15287_;
  assign new_n15289_ = ~new_n15160_ & ~new_n15163_;
  assign new_n15290_ = ~new_n15288_ & ~new_n15289_;
  assign new_n15291_ = new_n15212_ & ~new_n15290_;
  assign new_n15292_ = ~new_n15210_ & new_n15291_;
  assign new_n15293_ = ~new_n15286_ & ~new_n15292_;
  assign new_n15294_ = ~\b[37]  & ~new_n15293_;
  assign new_n15295_ = ~new_n14681_ & ~\quotient[18] ;
  assign new_n15296_ = ~new_n14691_ & new_n15158_;
  assign new_n15297_ = ~new_n15154_ & new_n15296_;
  assign new_n15298_ = ~new_n15155_ & ~new_n15158_;
  assign new_n15299_ = ~new_n15297_ & ~new_n15298_;
  assign new_n15300_ = new_n15212_ & ~new_n15299_;
  assign new_n15301_ = ~new_n15210_ & new_n15300_;
  assign new_n15302_ = ~new_n15295_ & ~new_n15301_;
  assign new_n15303_ = ~\b[36]  & ~new_n15302_;
  assign new_n15304_ = ~new_n14690_ & ~\quotient[18] ;
  assign new_n15305_ = ~new_n14700_ & new_n15153_;
  assign new_n15306_ = ~new_n15149_ & new_n15305_;
  assign new_n15307_ = ~new_n15150_ & ~new_n15153_;
  assign new_n15308_ = ~new_n15306_ & ~new_n15307_;
  assign new_n15309_ = new_n15212_ & ~new_n15308_;
  assign new_n15310_ = ~new_n15210_ & new_n15309_;
  assign new_n15311_ = ~new_n15304_ & ~new_n15310_;
  assign new_n15312_ = ~\b[35]  & ~new_n15311_;
  assign new_n15313_ = ~new_n14699_ & ~\quotient[18] ;
  assign new_n15314_ = ~new_n14709_ & new_n15148_;
  assign new_n15315_ = ~new_n15144_ & new_n15314_;
  assign new_n15316_ = ~new_n15145_ & ~new_n15148_;
  assign new_n15317_ = ~new_n15315_ & ~new_n15316_;
  assign new_n15318_ = new_n15212_ & ~new_n15317_;
  assign new_n15319_ = ~new_n15210_ & new_n15318_;
  assign new_n15320_ = ~new_n15313_ & ~new_n15319_;
  assign new_n15321_ = ~\b[34]  & ~new_n15320_;
  assign new_n15322_ = ~new_n14708_ & ~\quotient[18] ;
  assign new_n15323_ = ~new_n14718_ & new_n15143_;
  assign new_n15324_ = ~new_n15139_ & new_n15323_;
  assign new_n15325_ = ~new_n15140_ & ~new_n15143_;
  assign new_n15326_ = ~new_n15324_ & ~new_n15325_;
  assign new_n15327_ = new_n15212_ & ~new_n15326_;
  assign new_n15328_ = ~new_n15210_ & new_n15327_;
  assign new_n15329_ = ~new_n15322_ & ~new_n15328_;
  assign new_n15330_ = ~\b[33]  & ~new_n15329_;
  assign new_n15331_ = ~new_n14717_ & ~\quotient[18] ;
  assign new_n15332_ = ~new_n14727_ & new_n15138_;
  assign new_n15333_ = ~new_n15134_ & new_n15332_;
  assign new_n15334_ = ~new_n15135_ & ~new_n15138_;
  assign new_n15335_ = ~new_n15333_ & ~new_n15334_;
  assign new_n15336_ = new_n15212_ & ~new_n15335_;
  assign new_n15337_ = ~new_n15210_ & new_n15336_;
  assign new_n15338_ = ~new_n15331_ & ~new_n15337_;
  assign new_n15339_ = ~\b[32]  & ~new_n15338_;
  assign new_n15340_ = ~new_n14726_ & ~\quotient[18] ;
  assign new_n15341_ = ~new_n14736_ & new_n15133_;
  assign new_n15342_ = ~new_n15129_ & new_n15341_;
  assign new_n15343_ = ~new_n15130_ & ~new_n15133_;
  assign new_n15344_ = ~new_n15342_ & ~new_n15343_;
  assign new_n15345_ = new_n15212_ & ~new_n15344_;
  assign new_n15346_ = ~new_n15210_ & new_n15345_;
  assign new_n15347_ = ~new_n15340_ & ~new_n15346_;
  assign new_n15348_ = ~\b[31]  & ~new_n15347_;
  assign new_n15349_ = ~new_n14735_ & ~\quotient[18] ;
  assign new_n15350_ = ~new_n14745_ & new_n15128_;
  assign new_n15351_ = ~new_n15124_ & new_n15350_;
  assign new_n15352_ = ~new_n15125_ & ~new_n15128_;
  assign new_n15353_ = ~new_n15351_ & ~new_n15352_;
  assign new_n15354_ = new_n15212_ & ~new_n15353_;
  assign new_n15355_ = ~new_n15210_ & new_n15354_;
  assign new_n15356_ = ~new_n15349_ & ~new_n15355_;
  assign new_n15357_ = ~\b[30]  & ~new_n15356_;
  assign new_n15358_ = ~new_n14744_ & ~\quotient[18] ;
  assign new_n15359_ = ~new_n14754_ & new_n15123_;
  assign new_n15360_ = ~new_n15119_ & new_n15359_;
  assign new_n15361_ = ~new_n15120_ & ~new_n15123_;
  assign new_n15362_ = ~new_n15360_ & ~new_n15361_;
  assign new_n15363_ = new_n15212_ & ~new_n15362_;
  assign new_n15364_ = ~new_n15210_ & new_n15363_;
  assign new_n15365_ = ~new_n15358_ & ~new_n15364_;
  assign new_n15366_ = ~\b[29]  & ~new_n15365_;
  assign new_n15367_ = ~new_n14753_ & ~\quotient[18] ;
  assign new_n15368_ = ~new_n14763_ & new_n15118_;
  assign new_n15369_ = ~new_n15114_ & new_n15368_;
  assign new_n15370_ = ~new_n15115_ & ~new_n15118_;
  assign new_n15371_ = ~new_n15369_ & ~new_n15370_;
  assign new_n15372_ = new_n15212_ & ~new_n15371_;
  assign new_n15373_ = ~new_n15210_ & new_n15372_;
  assign new_n15374_ = ~new_n15367_ & ~new_n15373_;
  assign new_n15375_ = ~\b[28]  & ~new_n15374_;
  assign new_n15376_ = ~new_n14762_ & ~\quotient[18] ;
  assign new_n15377_ = ~new_n14772_ & new_n15113_;
  assign new_n15378_ = ~new_n15109_ & new_n15377_;
  assign new_n15379_ = ~new_n15110_ & ~new_n15113_;
  assign new_n15380_ = ~new_n15378_ & ~new_n15379_;
  assign new_n15381_ = new_n15212_ & ~new_n15380_;
  assign new_n15382_ = ~new_n15210_ & new_n15381_;
  assign new_n15383_ = ~new_n15376_ & ~new_n15382_;
  assign new_n15384_ = ~\b[27]  & ~new_n15383_;
  assign new_n15385_ = ~new_n14771_ & ~\quotient[18] ;
  assign new_n15386_ = ~new_n14781_ & new_n15108_;
  assign new_n15387_ = ~new_n15104_ & new_n15386_;
  assign new_n15388_ = ~new_n15105_ & ~new_n15108_;
  assign new_n15389_ = ~new_n15387_ & ~new_n15388_;
  assign new_n15390_ = new_n15212_ & ~new_n15389_;
  assign new_n15391_ = ~new_n15210_ & new_n15390_;
  assign new_n15392_ = ~new_n15385_ & ~new_n15391_;
  assign new_n15393_ = ~\b[26]  & ~new_n15392_;
  assign new_n15394_ = ~new_n14780_ & ~\quotient[18] ;
  assign new_n15395_ = ~new_n14790_ & new_n15103_;
  assign new_n15396_ = ~new_n15099_ & new_n15395_;
  assign new_n15397_ = ~new_n15100_ & ~new_n15103_;
  assign new_n15398_ = ~new_n15396_ & ~new_n15397_;
  assign new_n15399_ = new_n15212_ & ~new_n15398_;
  assign new_n15400_ = ~new_n15210_ & new_n15399_;
  assign new_n15401_ = ~new_n15394_ & ~new_n15400_;
  assign new_n15402_ = ~\b[25]  & ~new_n15401_;
  assign new_n15403_ = ~new_n14789_ & ~\quotient[18] ;
  assign new_n15404_ = ~new_n14799_ & new_n15098_;
  assign new_n15405_ = ~new_n15094_ & new_n15404_;
  assign new_n15406_ = ~new_n15095_ & ~new_n15098_;
  assign new_n15407_ = ~new_n15405_ & ~new_n15406_;
  assign new_n15408_ = new_n15212_ & ~new_n15407_;
  assign new_n15409_ = ~new_n15210_ & new_n15408_;
  assign new_n15410_ = ~new_n15403_ & ~new_n15409_;
  assign new_n15411_ = ~\b[24]  & ~new_n15410_;
  assign new_n15412_ = ~new_n14798_ & ~\quotient[18] ;
  assign new_n15413_ = ~new_n14808_ & new_n15093_;
  assign new_n15414_ = ~new_n15089_ & new_n15413_;
  assign new_n15415_ = ~new_n15090_ & ~new_n15093_;
  assign new_n15416_ = ~new_n15414_ & ~new_n15415_;
  assign new_n15417_ = new_n15212_ & ~new_n15416_;
  assign new_n15418_ = ~new_n15210_ & new_n15417_;
  assign new_n15419_ = ~new_n15412_ & ~new_n15418_;
  assign new_n15420_ = ~\b[23]  & ~new_n15419_;
  assign new_n15421_ = ~new_n14807_ & ~\quotient[18] ;
  assign new_n15422_ = ~new_n14817_ & new_n15088_;
  assign new_n15423_ = ~new_n15084_ & new_n15422_;
  assign new_n15424_ = ~new_n15085_ & ~new_n15088_;
  assign new_n15425_ = ~new_n15423_ & ~new_n15424_;
  assign new_n15426_ = new_n15212_ & ~new_n15425_;
  assign new_n15427_ = ~new_n15210_ & new_n15426_;
  assign new_n15428_ = ~new_n15421_ & ~new_n15427_;
  assign new_n15429_ = ~\b[22]  & ~new_n15428_;
  assign new_n15430_ = ~new_n14816_ & ~\quotient[18] ;
  assign new_n15431_ = ~new_n14826_ & new_n15083_;
  assign new_n15432_ = ~new_n15079_ & new_n15431_;
  assign new_n15433_ = ~new_n15080_ & ~new_n15083_;
  assign new_n15434_ = ~new_n15432_ & ~new_n15433_;
  assign new_n15435_ = new_n15212_ & ~new_n15434_;
  assign new_n15436_ = ~new_n15210_ & new_n15435_;
  assign new_n15437_ = ~new_n15430_ & ~new_n15436_;
  assign new_n15438_ = ~\b[21]  & ~new_n15437_;
  assign new_n15439_ = ~new_n14825_ & ~\quotient[18] ;
  assign new_n15440_ = ~new_n14835_ & new_n15078_;
  assign new_n15441_ = ~new_n15074_ & new_n15440_;
  assign new_n15442_ = ~new_n15075_ & ~new_n15078_;
  assign new_n15443_ = ~new_n15441_ & ~new_n15442_;
  assign new_n15444_ = new_n15212_ & ~new_n15443_;
  assign new_n15445_ = ~new_n15210_ & new_n15444_;
  assign new_n15446_ = ~new_n15439_ & ~new_n15445_;
  assign new_n15447_ = ~\b[20]  & ~new_n15446_;
  assign new_n15448_ = ~new_n14834_ & ~\quotient[18] ;
  assign new_n15449_ = ~new_n14844_ & new_n15073_;
  assign new_n15450_ = ~new_n15069_ & new_n15449_;
  assign new_n15451_ = ~new_n15070_ & ~new_n15073_;
  assign new_n15452_ = ~new_n15450_ & ~new_n15451_;
  assign new_n15453_ = new_n15212_ & ~new_n15452_;
  assign new_n15454_ = ~new_n15210_ & new_n15453_;
  assign new_n15455_ = ~new_n15448_ & ~new_n15454_;
  assign new_n15456_ = ~\b[19]  & ~new_n15455_;
  assign new_n15457_ = ~new_n14843_ & ~\quotient[18] ;
  assign new_n15458_ = ~new_n14853_ & new_n15068_;
  assign new_n15459_ = ~new_n15064_ & new_n15458_;
  assign new_n15460_ = ~new_n15065_ & ~new_n15068_;
  assign new_n15461_ = ~new_n15459_ & ~new_n15460_;
  assign new_n15462_ = new_n15212_ & ~new_n15461_;
  assign new_n15463_ = ~new_n15210_ & new_n15462_;
  assign new_n15464_ = ~new_n15457_ & ~new_n15463_;
  assign new_n15465_ = ~\b[18]  & ~new_n15464_;
  assign new_n15466_ = ~new_n14852_ & ~\quotient[18] ;
  assign new_n15467_ = ~new_n14862_ & new_n15063_;
  assign new_n15468_ = ~new_n15059_ & new_n15467_;
  assign new_n15469_ = ~new_n15060_ & ~new_n15063_;
  assign new_n15470_ = ~new_n15468_ & ~new_n15469_;
  assign new_n15471_ = new_n15212_ & ~new_n15470_;
  assign new_n15472_ = ~new_n15210_ & new_n15471_;
  assign new_n15473_ = ~new_n15466_ & ~new_n15472_;
  assign new_n15474_ = ~\b[17]  & ~new_n15473_;
  assign new_n15475_ = ~new_n14861_ & ~\quotient[18] ;
  assign new_n15476_ = ~new_n14871_ & new_n15058_;
  assign new_n15477_ = ~new_n15054_ & new_n15476_;
  assign new_n15478_ = ~new_n15055_ & ~new_n15058_;
  assign new_n15479_ = ~new_n15477_ & ~new_n15478_;
  assign new_n15480_ = new_n15212_ & ~new_n15479_;
  assign new_n15481_ = ~new_n15210_ & new_n15480_;
  assign new_n15482_ = ~new_n15475_ & ~new_n15481_;
  assign new_n15483_ = ~\b[16]  & ~new_n15482_;
  assign new_n15484_ = ~new_n14870_ & ~\quotient[18] ;
  assign new_n15485_ = ~new_n14880_ & new_n15053_;
  assign new_n15486_ = ~new_n15049_ & new_n15485_;
  assign new_n15487_ = ~new_n15050_ & ~new_n15053_;
  assign new_n15488_ = ~new_n15486_ & ~new_n15487_;
  assign new_n15489_ = new_n15212_ & ~new_n15488_;
  assign new_n15490_ = ~new_n15210_ & new_n15489_;
  assign new_n15491_ = ~new_n15484_ & ~new_n15490_;
  assign new_n15492_ = ~\b[15]  & ~new_n15491_;
  assign new_n15493_ = ~new_n14879_ & ~\quotient[18] ;
  assign new_n15494_ = ~new_n14889_ & new_n15048_;
  assign new_n15495_ = ~new_n15044_ & new_n15494_;
  assign new_n15496_ = ~new_n15045_ & ~new_n15048_;
  assign new_n15497_ = ~new_n15495_ & ~new_n15496_;
  assign new_n15498_ = new_n15212_ & ~new_n15497_;
  assign new_n15499_ = ~new_n15210_ & new_n15498_;
  assign new_n15500_ = ~new_n15493_ & ~new_n15499_;
  assign new_n15501_ = ~\b[14]  & ~new_n15500_;
  assign new_n15502_ = ~new_n14888_ & ~\quotient[18] ;
  assign new_n15503_ = ~new_n14898_ & new_n15043_;
  assign new_n15504_ = ~new_n15039_ & new_n15503_;
  assign new_n15505_ = ~new_n15040_ & ~new_n15043_;
  assign new_n15506_ = ~new_n15504_ & ~new_n15505_;
  assign new_n15507_ = new_n15212_ & ~new_n15506_;
  assign new_n15508_ = ~new_n15210_ & new_n15507_;
  assign new_n15509_ = ~new_n15502_ & ~new_n15508_;
  assign new_n15510_ = ~\b[13]  & ~new_n15509_;
  assign new_n15511_ = ~new_n14897_ & ~\quotient[18] ;
  assign new_n15512_ = ~new_n14907_ & new_n15038_;
  assign new_n15513_ = ~new_n15034_ & new_n15512_;
  assign new_n15514_ = ~new_n15035_ & ~new_n15038_;
  assign new_n15515_ = ~new_n15513_ & ~new_n15514_;
  assign new_n15516_ = new_n15212_ & ~new_n15515_;
  assign new_n15517_ = ~new_n15210_ & new_n15516_;
  assign new_n15518_ = ~new_n15511_ & ~new_n15517_;
  assign new_n15519_ = ~\b[12]  & ~new_n15518_;
  assign new_n15520_ = ~new_n14906_ & ~\quotient[18] ;
  assign new_n15521_ = ~new_n14916_ & new_n15033_;
  assign new_n15522_ = ~new_n15029_ & new_n15521_;
  assign new_n15523_ = ~new_n15030_ & ~new_n15033_;
  assign new_n15524_ = ~new_n15522_ & ~new_n15523_;
  assign new_n15525_ = new_n15212_ & ~new_n15524_;
  assign new_n15526_ = ~new_n15210_ & new_n15525_;
  assign new_n15527_ = ~new_n15520_ & ~new_n15526_;
  assign new_n15528_ = ~\b[11]  & ~new_n15527_;
  assign new_n15529_ = ~new_n14915_ & ~\quotient[18] ;
  assign new_n15530_ = ~new_n14925_ & new_n15028_;
  assign new_n15531_ = ~new_n15024_ & new_n15530_;
  assign new_n15532_ = ~new_n15025_ & ~new_n15028_;
  assign new_n15533_ = ~new_n15531_ & ~new_n15532_;
  assign new_n15534_ = new_n15212_ & ~new_n15533_;
  assign new_n15535_ = ~new_n15210_ & new_n15534_;
  assign new_n15536_ = ~new_n15529_ & ~new_n15535_;
  assign new_n15537_ = ~\b[10]  & ~new_n15536_;
  assign new_n15538_ = ~new_n14924_ & ~\quotient[18] ;
  assign new_n15539_ = ~new_n14934_ & new_n15023_;
  assign new_n15540_ = ~new_n15019_ & new_n15539_;
  assign new_n15541_ = ~new_n15020_ & ~new_n15023_;
  assign new_n15542_ = ~new_n15540_ & ~new_n15541_;
  assign new_n15543_ = new_n15212_ & ~new_n15542_;
  assign new_n15544_ = ~new_n15210_ & new_n15543_;
  assign new_n15545_ = ~new_n15538_ & ~new_n15544_;
  assign new_n15546_ = ~\b[9]  & ~new_n15545_;
  assign new_n15547_ = ~new_n14933_ & ~\quotient[18] ;
  assign new_n15548_ = ~new_n14943_ & new_n15018_;
  assign new_n15549_ = ~new_n15014_ & new_n15548_;
  assign new_n15550_ = ~new_n15015_ & ~new_n15018_;
  assign new_n15551_ = ~new_n15549_ & ~new_n15550_;
  assign new_n15552_ = new_n15212_ & ~new_n15551_;
  assign new_n15553_ = ~new_n15210_ & new_n15552_;
  assign new_n15554_ = ~new_n15547_ & ~new_n15553_;
  assign new_n15555_ = ~\b[8]  & ~new_n15554_;
  assign new_n15556_ = ~new_n14942_ & ~\quotient[18] ;
  assign new_n15557_ = ~new_n14952_ & new_n15013_;
  assign new_n15558_ = ~new_n15009_ & new_n15557_;
  assign new_n15559_ = ~new_n15010_ & ~new_n15013_;
  assign new_n15560_ = ~new_n15558_ & ~new_n15559_;
  assign new_n15561_ = new_n15212_ & ~new_n15560_;
  assign new_n15562_ = ~new_n15210_ & new_n15561_;
  assign new_n15563_ = ~new_n15556_ & ~new_n15562_;
  assign new_n15564_ = ~\b[7]  & ~new_n15563_;
  assign new_n15565_ = ~new_n14951_ & ~\quotient[18] ;
  assign new_n15566_ = ~new_n14961_ & new_n15008_;
  assign new_n15567_ = ~new_n15004_ & new_n15566_;
  assign new_n15568_ = ~new_n15005_ & ~new_n15008_;
  assign new_n15569_ = ~new_n15567_ & ~new_n15568_;
  assign new_n15570_ = new_n15212_ & ~new_n15569_;
  assign new_n15571_ = ~new_n15210_ & new_n15570_;
  assign new_n15572_ = ~new_n15565_ & ~new_n15571_;
  assign new_n15573_ = ~\b[6]  & ~new_n15572_;
  assign new_n15574_ = ~new_n14960_ & ~\quotient[18] ;
  assign new_n15575_ = ~new_n14970_ & new_n15003_;
  assign new_n15576_ = ~new_n14999_ & new_n15575_;
  assign new_n15577_ = ~new_n15000_ & ~new_n15003_;
  assign new_n15578_ = ~new_n15576_ & ~new_n15577_;
  assign new_n15579_ = new_n15212_ & ~new_n15578_;
  assign new_n15580_ = ~new_n15210_ & new_n15579_;
  assign new_n15581_ = ~new_n15574_ & ~new_n15580_;
  assign new_n15582_ = ~\b[5]  & ~new_n15581_;
  assign new_n15583_ = ~new_n14969_ & ~\quotient[18] ;
  assign new_n15584_ = ~new_n14978_ & new_n14998_;
  assign new_n15585_ = ~new_n14994_ & new_n15584_;
  assign new_n15586_ = ~new_n14995_ & ~new_n14998_;
  assign new_n15587_ = ~new_n15585_ & ~new_n15586_;
  assign new_n15588_ = new_n15212_ & ~new_n15587_;
  assign new_n15589_ = ~new_n15210_ & new_n15588_;
  assign new_n15590_ = ~new_n15583_ & ~new_n15589_;
  assign new_n15591_ = ~\b[4]  & ~new_n15590_;
  assign new_n15592_ = ~new_n14977_ & ~\quotient[18] ;
  assign new_n15593_ = ~new_n14989_ & new_n14993_;
  assign new_n15594_ = ~new_n14988_ & new_n15593_;
  assign new_n15595_ = ~new_n14990_ & ~new_n14993_;
  assign new_n15596_ = ~new_n15594_ & ~new_n15595_;
  assign new_n15597_ = new_n15212_ & ~new_n15596_;
  assign new_n15598_ = ~new_n15210_ & new_n15597_;
  assign new_n15599_ = ~new_n15592_ & ~new_n15598_;
  assign new_n15600_ = ~\b[3]  & ~new_n15599_;
  assign new_n15601_ = ~new_n14982_ & ~\quotient[18] ;
  assign new_n15602_ = ~new_n14985_ & new_n14987_;
  assign new_n15603_ = ~new_n14983_ & new_n15602_;
  assign new_n15604_ = new_n15212_ & ~new_n15603_;
  assign new_n15605_ = ~new_n14988_ & new_n15604_;
  assign new_n15606_ = ~new_n15210_ & new_n15605_;
  assign new_n15607_ = ~new_n15601_ & ~new_n15606_;
  assign new_n15608_ = ~\b[2]  & ~new_n15607_;
  assign new_n15609_ = \b[0]  & ~\b[46] ;
  assign new_n15610_ = new_n417_ & new_n15609_;
  assign new_n15611_ = new_n400_ & new_n15610_;
  assign new_n15612_ = new_n595_ & new_n15611_;
  assign new_n15613_ = ~new_n15210_ & new_n15612_;
  assign new_n15614_ = \a[18]  & ~new_n15613_;
  assign new_n15615_ = new_n300_ & new_n14987_;
  assign new_n15616_ = new_n298_ & new_n15615_;
  assign new_n15617_ = new_n288_ & new_n15616_;
  assign new_n15618_ = ~new_n15210_ & new_n15617_;
  assign new_n15619_ = ~new_n15614_ & ~new_n15618_;
  assign new_n15620_ = \b[1]  & ~new_n15619_;
  assign new_n15621_ = ~\b[1]  & ~new_n15618_;
  assign new_n15622_ = ~new_n15614_ & new_n15621_;
  assign new_n15623_ = ~new_n15620_ & ~new_n15622_;
  assign new_n15624_ = ~\a[17]  & \b[0] ;
  assign new_n15625_ = ~new_n15623_ & ~new_n15624_;
  assign new_n15626_ = ~\b[1]  & ~new_n15619_;
  assign new_n15627_ = ~new_n15625_ & ~new_n15626_;
  assign new_n15628_ = \b[2]  & ~new_n15606_;
  assign new_n15629_ = ~new_n15601_ & new_n15628_;
  assign new_n15630_ = ~new_n15608_ & ~new_n15629_;
  assign new_n15631_ = ~new_n15627_ & new_n15630_;
  assign new_n15632_ = ~new_n15608_ & ~new_n15631_;
  assign new_n15633_ = \b[3]  & ~new_n15598_;
  assign new_n15634_ = ~new_n15592_ & new_n15633_;
  assign new_n15635_ = ~new_n15600_ & ~new_n15634_;
  assign new_n15636_ = ~new_n15632_ & new_n15635_;
  assign new_n15637_ = ~new_n15600_ & ~new_n15636_;
  assign new_n15638_ = \b[4]  & ~new_n15589_;
  assign new_n15639_ = ~new_n15583_ & new_n15638_;
  assign new_n15640_ = ~new_n15591_ & ~new_n15639_;
  assign new_n15641_ = ~new_n15637_ & new_n15640_;
  assign new_n15642_ = ~new_n15591_ & ~new_n15641_;
  assign new_n15643_ = \b[5]  & ~new_n15580_;
  assign new_n15644_ = ~new_n15574_ & new_n15643_;
  assign new_n15645_ = ~new_n15582_ & ~new_n15644_;
  assign new_n15646_ = ~new_n15642_ & new_n15645_;
  assign new_n15647_ = ~new_n15582_ & ~new_n15646_;
  assign new_n15648_ = \b[6]  & ~new_n15571_;
  assign new_n15649_ = ~new_n15565_ & new_n15648_;
  assign new_n15650_ = ~new_n15573_ & ~new_n15649_;
  assign new_n15651_ = ~new_n15647_ & new_n15650_;
  assign new_n15652_ = ~new_n15573_ & ~new_n15651_;
  assign new_n15653_ = \b[7]  & ~new_n15562_;
  assign new_n15654_ = ~new_n15556_ & new_n15653_;
  assign new_n15655_ = ~new_n15564_ & ~new_n15654_;
  assign new_n15656_ = ~new_n15652_ & new_n15655_;
  assign new_n15657_ = ~new_n15564_ & ~new_n15656_;
  assign new_n15658_ = \b[8]  & ~new_n15553_;
  assign new_n15659_ = ~new_n15547_ & new_n15658_;
  assign new_n15660_ = ~new_n15555_ & ~new_n15659_;
  assign new_n15661_ = ~new_n15657_ & new_n15660_;
  assign new_n15662_ = ~new_n15555_ & ~new_n15661_;
  assign new_n15663_ = \b[9]  & ~new_n15544_;
  assign new_n15664_ = ~new_n15538_ & new_n15663_;
  assign new_n15665_ = ~new_n15546_ & ~new_n15664_;
  assign new_n15666_ = ~new_n15662_ & new_n15665_;
  assign new_n15667_ = ~new_n15546_ & ~new_n15666_;
  assign new_n15668_ = \b[10]  & ~new_n15535_;
  assign new_n15669_ = ~new_n15529_ & new_n15668_;
  assign new_n15670_ = ~new_n15537_ & ~new_n15669_;
  assign new_n15671_ = ~new_n15667_ & new_n15670_;
  assign new_n15672_ = ~new_n15537_ & ~new_n15671_;
  assign new_n15673_ = \b[11]  & ~new_n15526_;
  assign new_n15674_ = ~new_n15520_ & new_n15673_;
  assign new_n15675_ = ~new_n15528_ & ~new_n15674_;
  assign new_n15676_ = ~new_n15672_ & new_n15675_;
  assign new_n15677_ = ~new_n15528_ & ~new_n15676_;
  assign new_n15678_ = \b[12]  & ~new_n15517_;
  assign new_n15679_ = ~new_n15511_ & new_n15678_;
  assign new_n15680_ = ~new_n15519_ & ~new_n15679_;
  assign new_n15681_ = ~new_n15677_ & new_n15680_;
  assign new_n15682_ = ~new_n15519_ & ~new_n15681_;
  assign new_n15683_ = \b[13]  & ~new_n15508_;
  assign new_n15684_ = ~new_n15502_ & new_n15683_;
  assign new_n15685_ = ~new_n15510_ & ~new_n15684_;
  assign new_n15686_ = ~new_n15682_ & new_n15685_;
  assign new_n15687_ = ~new_n15510_ & ~new_n15686_;
  assign new_n15688_ = \b[14]  & ~new_n15499_;
  assign new_n15689_ = ~new_n15493_ & new_n15688_;
  assign new_n15690_ = ~new_n15501_ & ~new_n15689_;
  assign new_n15691_ = ~new_n15687_ & new_n15690_;
  assign new_n15692_ = ~new_n15501_ & ~new_n15691_;
  assign new_n15693_ = \b[15]  & ~new_n15490_;
  assign new_n15694_ = ~new_n15484_ & new_n15693_;
  assign new_n15695_ = ~new_n15492_ & ~new_n15694_;
  assign new_n15696_ = ~new_n15692_ & new_n15695_;
  assign new_n15697_ = ~new_n15492_ & ~new_n15696_;
  assign new_n15698_ = \b[16]  & ~new_n15481_;
  assign new_n15699_ = ~new_n15475_ & new_n15698_;
  assign new_n15700_ = ~new_n15483_ & ~new_n15699_;
  assign new_n15701_ = ~new_n15697_ & new_n15700_;
  assign new_n15702_ = ~new_n15483_ & ~new_n15701_;
  assign new_n15703_ = \b[17]  & ~new_n15472_;
  assign new_n15704_ = ~new_n15466_ & new_n15703_;
  assign new_n15705_ = ~new_n15474_ & ~new_n15704_;
  assign new_n15706_ = ~new_n15702_ & new_n15705_;
  assign new_n15707_ = ~new_n15474_ & ~new_n15706_;
  assign new_n15708_ = \b[18]  & ~new_n15463_;
  assign new_n15709_ = ~new_n15457_ & new_n15708_;
  assign new_n15710_ = ~new_n15465_ & ~new_n15709_;
  assign new_n15711_ = ~new_n15707_ & new_n15710_;
  assign new_n15712_ = ~new_n15465_ & ~new_n15711_;
  assign new_n15713_ = \b[19]  & ~new_n15454_;
  assign new_n15714_ = ~new_n15448_ & new_n15713_;
  assign new_n15715_ = ~new_n15456_ & ~new_n15714_;
  assign new_n15716_ = ~new_n15712_ & new_n15715_;
  assign new_n15717_ = ~new_n15456_ & ~new_n15716_;
  assign new_n15718_ = \b[20]  & ~new_n15445_;
  assign new_n15719_ = ~new_n15439_ & new_n15718_;
  assign new_n15720_ = ~new_n15447_ & ~new_n15719_;
  assign new_n15721_ = ~new_n15717_ & new_n15720_;
  assign new_n15722_ = ~new_n15447_ & ~new_n15721_;
  assign new_n15723_ = \b[21]  & ~new_n15436_;
  assign new_n15724_ = ~new_n15430_ & new_n15723_;
  assign new_n15725_ = ~new_n15438_ & ~new_n15724_;
  assign new_n15726_ = ~new_n15722_ & new_n15725_;
  assign new_n15727_ = ~new_n15438_ & ~new_n15726_;
  assign new_n15728_ = \b[22]  & ~new_n15427_;
  assign new_n15729_ = ~new_n15421_ & new_n15728_;
  assign new_n15730_ = ~new_n15429_ & ~new_n15729_;
  assign new_n15731_ = ~new_n15727_ & new_n15730_;
  assign new_n15732_ = ~new_n15429_ & ~new_n15731_;
  assign new_n15733_ = \b[23]  & ~new_n15418_;
  assign new_n15734_ = ~new_n15412_ & new_n15733_;
  assign new_n15735_ = ~new_n15420_ & ~new_n15734_;
  assign new_n15736_ = ~new_n15732_ & new_n15735_;
  assign new_n15737_ = ~new_n15420_ & ~new_n15736_;
  assign new_n15738_ = \b[24]  & ~new_n15409_;
  assign new_n15739_ = ~new_n15403_ & new_n15738_;
  assign new_n15740_ = ~new_n15411_ & ~new_n15739_;
  assign new_n15741_ = ~new_n15737_ & new_n15740_;
  assign new_n15742_ = ~new_n15411_ & ~new_n15741_;
  assign new_n15743_ = \b[25]  & ~new_n15400_;
  assign new_n15744_ = ~new_n15394_ & new_n15743_;
  assign new_n15745_ = ~new_n15402_ & ~new_n15744_;
  assign new_n15746_ = ~new_n15742_ & new_n15745_;
  assign new_n15747_ = ~new_n15402_ & ~new_n15746_;
  assign new_n15748_ = \b[26]  & ~new_n15391_;
  assign new_n15749_ = ~new_n15385_ & new_n15748_;
  assign new_n15750_ = ~new_n15393_ & ~new_n15749_;
  assign new_n15751_ = ~new_n15747_ & new_n15750_;
  assign new_n15752_ = ~new_n15393_ & ~new_n15751_;
  assign new_n15753_ = \b[27]  & ~new_n15382_;
  assign new_n15754_ = ~new_n15376_ & new_n15753_;
  assign new_n15755_ = ~new_n15384_ & ~new_n15754_;
  assign new_n15756_ = ~new_n15752_ & new_n15755_;
  assign new_n15757_ = ~new_n15384_ & ~new_n15756_;
  assign new_n15758_ = \b[28]  & ~new_n15373_;
  assign new_n15759_ = ~new_n15367_ & new_n15758_;
  assign new_n15760_ = ~new_n15375_ & ~new_n15759_;
  assign new_n15761_ = ~new_n15757_ & new_n15760_;
  assign new_n15762_ = ~new_n15375_ & ~new_n15761_;
  assign new_n15763_ = \b[29]  & ~new_n15364_;
  assign new_n15764_ = ~new_n15358_ & new_n15763_;
  assign new_n15765_ = ~new_n15366_ & ~new_n15764_;
  assign new_n15766_ = ~new_n15762_ & new_n15765_;
  assign new_n15767_ = ~new_n15366_ & ~new_n15766_;
  assign new_n15768_ = \b[30]  & ~new_n15355_;
  assign new_n15769_ = ~new_n15349_ & new_n15768_;
  assign new_n15770_ = ~new_n15357_ & ~new_n15769_;
  assign new_n15771_ = ~new_n15767_ & new_n15770_;
  assign new_n15772_ = ~new_n15357_ & ~new_n15771_;
  assign new_n15773_ = \b[31]  & ~new_n15346_;
  assign new_n15774_ = ~new_n15340_ & new_n15773_;
  assign new_n15775_ = ~new_n15348_ & ~new_n15774_;
  assign new_n15776_ = ~new_n15772_ & new_n15775_;
  assign new_n15777_ = ~new_n15348_ & ~new_n15776_;
  assign new_n15778_ = \b[32]  & ~new_n15337_;
  assign new_n15779_ = ~new_n15331_ & new_n15778_;
  assign new_n15780_ = ~new_n15339_ & ~new_n15779_;
  assign new_n15781_ = ~new_n15777_ & new_n15780_;
  assign new_n15782_ = ~new_n15339_ & ~new_n15781_;
  assign new_n15783_ = \b[33]  & ~new_n15328_;
  assign new_n15784_ = ~new_n15322_ & new_n15783_;
  assign new_n15785_ = ~new_n15330_ & ~new_n15784_;
  assign new_n15786_ = ~new_n15782_ & new_n15785_;
  assign new_n15787_ = ~new_n15330_ & ~new_n15786_;
  assign new_n15788_ = \b[34]  & ~new_n15319_;
  assign new_n15789_ = ~new_n15313_ & new_n15788_;
  assign new_n15790_ = ~new_n15321_ & ~new_n15789_;
  assign new_n15791_ = ~new_n15787_ & new_n15790_;
  assign new_n15792_ = ~new_n15321_ & ~new_n15791_;
  assign new_n15793_ = \b[35]  & ~new_n15310_;
  assign new_n15794_ = ~new_n15304_ & new_n15793_;
  assign new_n15795_ = ~new_n15312_ & ~new_n15794_;
  assign new_n15796_ = ~new_n15792_ & new_n15795_;
  assign new_n15797_ = ~new_n15312_ & ~new_n15796_;
  assign new_n15798_ = \b[36]  & ~new_n15301_;
  assign new_n15799_ = ~new_n15295_ & new_n15798_;
  assign new_n15800_ = ~new_n15303_ & ~new_n15799_;
  assign new_n15801_ = ~new_n15797_ & new_n15800_;
  assign new_n15802_ = ~new_n15303_ & ~new_n15801_;
  assign new_n15803_ = \b[37]  & ~new_n15292_;
  assign new_n15804_ = ~new_n15286_ & new_n15803_;
  assign new_n15805_ = ~new_n15294_ & ~new_n15804_;
  assign new_n15806_ = ~new_n15802_ & new_n15805_;
  assign new_n15807_ = ~new_n15294_ & ~new_n15806_;
  assign new_n15808_ = \b[38]  & ~new_n15283_;
  assign new_n15809_ = ~new_n15277_ & new_n15808_;
  assign new_n15810_ = ~new_n15285_ & ~new_n15809_;
  assign new_n15811_ = ~new_n15807_ & new_n15810_;
  assign new_n15812_ = ~new_n15285_ & ~new_n15811_;
  assign new_n15813_ = \b[39]  & ~new_n15274_;
  assign new_n15814_ = ~new_n15268_ & new_n15813_;
  assign new_n15815_ = ~new_n15276_ & ~new_n15814_;
  assign new_n15816_ = ~new_n15812_ & new_n15815_;
  assign new_n15817_ = ~new_n15276_ & ~new_n15816_;
  assign new_n15818_ = \b[40]  & ~new_n15265_;
  assign new_n15819_ = ~new_n15259_ & new_n15818_;
  assign new_n15820_ = ~new_n15267_ & ~new_n15819_;
  assign new_n15821_ = ~new_n15817_ & new_n15820_;
  assign new_n15822_ = ~new_n15267_ & ~new_n15821_;
  assign new_n15823_ = \b[41]  & ~new_n15256_;
  assign new_n15824_ = ~new_n15250_ & new_n15823_;
  assign new_n15825_ = ~new_n15258_ & ~new_n15824_;
  assign new_n15826_ = ~new_n15822_ & new_n15825_;
  assign new_n15827_ = ~new_n15258_ & ~new_n15826_;
  assign new_n15828_ = \b[42]  & ~new_n15247_;
  assign new_n15829_ = ~new_n15241_ & new_n15828_;
  assign new_n15830_ = ~new_n15249_ & ~new_n15829_;
  assign new_n15831_ = ~new_n15827_ & new_n15830_;
  assign new_n15832_ = ~new_n15249_ & ~new_n15831_;
  assign new_n15833_ = \b[43]  & ~new_n15238_;
  assign new_n15834_ = ~new_n15232_ & new_n15833_;
  assign new_n15835_ = ~new_n15240_ & ~new_n15834_;
  assign new_n15836_ = ~new_n15832_ & new_n15835_;
  assign new_n15837_ = ~new_n15240_ & ~new_n15836_;
  assign new_n15838_ = \b[44]  & ~new_n15229_;
  assign new_n15839_ = ~new_n15223_ & new_n15838_;
  assign new_n15840_ = ~new_n15231_ & ~new_n15839_;
  assign new_n15841_ = ~new_n15837_ & new_n15840_;
  assign new_n15842_ = ~new_n15231_ & ~new_n15841_;
  assign new_n15843_ = \b[45]  & ~new_n15220_;
  assign new_n15844_ = ~new_n15214_ & new_n15843_;
  assign new_n15845_ = ~new_n15222_ & ~new_n15844_;
  assign new_n15846_ = ~new_n15842_ & new_n15845_;
  assign new_n15847_ = ~new_n15222_ & ~new_n15846_;
  assign new_n15848_ = ~new_n14599_ & ~\quotient[18] ;
  assign new_n15849_ = ~new_n14601_ & new_n15208_;
  assign new_n15850_ = ~new_n15204_ & new_n15849_;
  assign new_n15851_ = ~new_n15205_ & ~new_n15208_;
  assign new_n15852_ = ~new_n15850_ & ~new_n15851_;
  assign new_n15853_ = \quotient[18]  & ~new_n15852_;
  assign new_n15854_ = ~new_n15848_ & ~new_n15853_;
  assign new_n15855_ = ~\b[46]  & ~new_n15854_;
  assign new_n15856_ = \b[46]  & ~new_n15848_;
  assign new_n15857_ = ~new_n15853_ & new_n15856_;
  assign new_n15858_ = new_n400_ & new_n417_;
  assign new_n15859_ = new_n595_ & new_n15858_;
  assign new_n15860_ = ~new_n15857_ & new_n15859_;
  assign new_n15861_ = ~new_n15855_ & new_n15860_;
  assign new_n15862_ = ~new_n15847_ & new_n15861_;
  assign new_n15863_ = new_n15212_ & ~new_n15854_;
  assign \quotient[17]  = new_n15862_ | new_n15863_;
  assign new_n15865_ = ~new_n15231_ & new_n15845_;
  assign new_n15866_ = ~new_n15841_ & new_n15865_;
  assign new_n15867_ = ~new_n15842_ & ~new_n15845_;
  assign new_n15868_ = ~new_n15866_ & ~new_n15867_;
  assign new_n15869_ = \quotient[17]  & ~new_n15868_;
  assign new_n15870_ = ~new_n15221_ & ~new_n15863_;
  assign new_n15871_ = ~new_n15862_ & new_n15870_;
  assign new_n15872_ = ~new_n15869_ & ~new_n15871_;
  assign new_n15873_ = ~\b[46]  & ~new_n15872_;
  assign new_n15874_ = ~new_n15240_ & new_n15840_;
  assign new_n15875_ = ~new_n15836_ & new_n15874_;
  assign new_n15876_ = ~new_n15837_ & ~new_n15840_;
  assign new_n15877_ = ~new_n15875_ & ~new_n15876_;
  assign new_n15878_ = \quotient[17]  & ~new_n15877_;
  assign new_n15879_ = ~new_n15230_ & ~new_n15863_;
  assign new_n15880_ = ~new_n15862_ & new_n15879_;
  assign new_n15881_ = ~new_n15878_ & ~new_n15880_;
  assign new_n15882_ = ~\b[45]  & ~new_n15881_;
  assign new_n15883_ = ~new_n15249_ & new_n15835_;
  assign new_n15884_ = ~new_n15831_ & new_n15883_;
  assign new_n15885_ = ~new_n15832_ & ~new_n15835_;
  assign new_n15886_ = ~new_n15884_ & ~new_n15885_;
  assign new_n15887_ = \quotient[17]  & ~new_n15886_;
  assign new_n15888_ = ~new_n15239_ & ~new_n15863_;
  assign new_n15889_ = ~new_n15862_ & new_n15888_;
  assign new_n15890_ = ~new_n15887_ & ~new_n15889_;
  assign new_n15891_ = ~\b[44]  & ~new_n15890_;
  assign new_n15892_ = ~new_n15258_ & new_n15830_;
  assign new_n15893_ = ~new_n15826_ & new_n15892_;
  assign new_n15894_ = ~new_n15827_ & ~new_n15830_;
  assign new_n15895_ = ~new_n15893_ & ~new_n15894_;
  assign new_n15896_ = \quotient[17]  & ~new_n15895_;
  assign new_n15897_ = ~new_n15248_ & ~new_n15863_;
  assign new_n15898_ = ~new_n15862_ & new_n15897_;
  assign new_n15899_ = ~new_n15896_ & ~new_n15898_;
  assign new_n15900_ = ~\b[43]  & ~new_n15899_;
  assign new_n15901_ = ~new_n15267_ & new_n15825_;
  assign new_n15902_ = ~new_n15821_ & new_n15901_;
  assign new_n15903_ = ~new_n15822_ & ~new_n15825_;
  assign new_n15904_ = ~new_n15902_ & ~new_n15903_;
  assign new_n15905_ = \quotient[17]  & ~new_n15904_;
  assign new_n15906_ = ~new_n15257_ & ~new_n15863_;
  assign new_n15907_ = ~new_n15862_ & new_n15906_;
  assign new_n15908_ = ~new_n15905_ & ~new_n15907_;
  assign new_n15909_ = ~\b[42]  & ~new_n15908_;
  assign new_n15910_ = ~new_n15276_ & new_n15820_;
  assign new_n15911_ = ~new_n15816_ & new_n15910_;
  assign new_n15912_ = ~new_n15817_ & ~new_n15820_;
  assign new_n15913_ = ~new_n15911_ & ~new_n15912_;
  assign new_n15914_ = \quotient[17]  & ~new_n15913_;
  assign new_n15915_ = ~new_n15266_ & ~new_n15863_;
  assign new_n15916_ = ~new_n15862_ & new_n15915_;
  assign new_n15917_ = ~new_n15914_ & ~new_n15916_;
  assign new_n15918_ = ~\b[41]  & ~new_n15917_;
  assign new_n15919_ = ~new_n15285_ & new_n15815_;
  assign new_n15920_ = ~new_n15811_ & new_n15919_;
  assign new_n15921_ = ~new_n15812_ & ~new_n15815_;
  assign new_n15922_ = ~new_n15920_ & ~new_n15921_;
  assign new_n15923_ = \quotient[17]  & ~new_n15922_;
  assign new_n15924_ = ~new_n15275_ & ~new_n15863_;
  assign new_n15925_ = ~new_n15862_ & new_n15924_;
  assign new_n15926_ = ~new_n15923_ & ~new_n15925_;
  assign new_n15927_ = ~\b[40]  & ~new_n15926_;
  assign new_n15928_ = ~new_n15294_ & new_n15810_;
  assign new_n15929_ = ~new_n15806_ & new_n15928_;
  assign new_n15930_ = ~new_n15807_ & ~new_n15810_;
  assign new_n15931_ = ~new_n15929_ & ~new_n15930_;
  assign new_n15932_ = \quotient[17]  & ~new_n15931_;
  assign new_n15933_ = ~new_n15284_ & ~new_n15863_;
  assign new_n15934_ = ~new_n15862_ & new_n15933_;
  assign new_n15935_ = ~new_n15932_ & ~new_n15934_;
  assign new_n15936_ = ~\b[39]  & ~new_n15935_;
  assign new_n15937_ = ~new_n15303_ & new_n15805_;
  assign new_n15938_ = ~new_n15801_ & new_n15937_;
  assign new_n15939_ = ~new_n15802_ & ~new_n15805_;
  assign new_n15940_ = ~new_n15938_ & ~new_n15939_;
  assign new_n15941_ = \quotient[17]  & ~new_n15940_;
  assign new_n15942_ = ~new_n15293_ & ~new_n15863_;
  assign new_n15943_ = ~new_n15862_ & new_n15942_;
  assign new_n15944_ = ~new_n15941_ & ~new_n15943_;
  assign new_n15945_ = ~\b[38]  & ~new_n15944_;
  assign new_n15946_ = ~new_n15312_ & new_n15800_;
  assign new_n15947_ = ~new_n15796_ & new_n15946_;
  assign new_n15948_ = ~new_n15797_ & ~new_n15800_;
  assign new_n15949_ = ~new_n15947_ & ~new_n15948_;
  assign new_n15950_ = \quotient[17]  & ~new_n15949_;
  assign new_n15951_ = ~new_n15302_ & ~new_n15863_;
  assign new_n15952_ = ~new_n15862_ & new_n15951_;
  assign new_n15953_ = ~new_n15950_ & ~new_n15952_;
  assign new_n15954_ = ~\b[37]  & ~new_n15953_;
  assign new_n15955_ = ~new_n15321_ & new_n15795_;
  assign new_n15956_ = ~new_n15791_ & new_n15955_;
  assign new_n15957_ = ~new_n15792_ & ~new_n15795_;
  assign new_n15958_ = ~new_n15956_ & ~new_n15957_;
  assign new_n15959_ = \quotient[17]  & ~new_n15958_;
  assign new_n15960_ = ~new_n15311_ & ~new_n15863_;
  assign new_n15961_ = ~new_n15862_ & new_n15960_;
  assign new_n15962_ = ~new_n15959_ & ~new_n15961_;
  assign new_n15963_ = ~\b[36]  & ~new_n15962_;
  assign new_n15964_ = ~new_n15330_ & new_n15790_;
  assign new_n15965_ = ~new_n15786_ & new_n15964_;
  assign new_n15966_ = ~new_n15787_ & ~new_n15790_;
  assign new_n15967_ = ~new_n15965_ & ~new_n15966_;
  assign new_n15968_ = \quotient[17]  & ~new_n15967_;
  assign new_n15969_ = ~new_n15320_ & ~new_n15863_;
  assign new_n15970_ = ~new_n15862_ & new_n15969_;
  assign new_n15971_ = ~new_n15968_ & ~new_n15970_;
  assign new_n15972_ = ~\b[35]  & ~new_n15971_;
  assign new_n15973_ = ~new_n15339_ & new_n15785_;
  assign new_n15974_ = ~new_n15781_ & new_n15973_;
  assign new_n15975_ = ~new_n15782_ & ~new_n15785_;
  assign new_n15976_ = ~new_n15974_ & ~new_n15975_;
  assign new_n15977_ = \quotient[17]  & ~new_n15976_;
  assign new_n15978_ = ~new_n15329_ & ~new_n15863_;
  assign new_n15979_ = ~new_n15862_ & new_n15978_;
  assign new_n15980_ = ~new_n15977_ & ~new_n15979_;
  assign new_n15981_ = ~\b[34]  & ~new_n15980_;
  assign new_n15982_ = ~new_n15348_ & new_n15780_;
  assign new_n15983_ = ~new_n15776_ & new_n15982_;
  assign new_n15984_ = ~new_n15777_ & ~new_n15780_;
  assign new_n15985_ = ~new_n15983_ & ~new_n15984_;
  assign new_n15986_ = \quotient[17]  & ~new_n15985_;
  assign new_n15987_ = ~new_n15338_ & ~new_n15863_;
  assign new_n15988_ = ~new_n15862_ & new_n15987_;
  assign new_n15989_ = ~new_n15986_ & ~new_n15988_;
  assign new_n15990_ = ~\b[33]  & ~new_n15989_;
  assign new_n15991_ = ~new_n15357_ & new_n15775_;
  assign new_n15992_ = ~new_n15771_ & new_n15991_;
  assign new_n15993_ = ~new_n15772_ & ~new_n15775_;
  assign new_n15994_ = ~new_n15992_ & ~new_n15993_;
  assign new_n15995_ = \quotient[17]  & ~new_n15994_;
  assign new_n15996_ = ~new_n15347_ & ~new_n15863_;
  assign new_n15997_ = ~new_n15862_ & new_n15996_;
  assign new_n15998_ = ~new_n15995_ & ~new_n15997_;
  assign new_n15999_ = ~\b[32]  & ~new_n15998_;
  assign new_n16000_ = ~new_n15366_ & new_n15770_;
  assign new_n16001_ = ~new_n15766_ & new_n16000_;
  assign new_n16002_ = ~new_n15767_ & ~new_n15770_;
  assign new_n16003_ = ~new_n16001_ & ~new_n16002_;
  assign new_n16004_ = \quotient[17]  & ~new_n16003_;
  assign new_n16005_ = ~new_n15356_ & ~new_n15863_;
  assign new_n16006_ = ~new_n15862_ & new_n16005_;
  assign new_n16007_ = ~new_n16004_ & ~new_n16006_;
  assign new_n16008_ = ~\b[31]  & ~new_n16007_;
  assign new_n16009_ = ~new_n15375_ & new_n15765_;
  assign new_n16010_ = ~new_n15761_ & new_n16009_;
  assign new_n16011_ = ~new_n15762_ & ~new_n15765_;
  assign new_n16012_ = ~new_n16010_ & ~new_n16011_;
  assign new_n16013_ = \quotient[17]  & ~new_n16012_;
  assign new_n16014_ = ~new_n15365_ & ~new_n15863_;
  assign new_n16015_ = ~new_n15862_ & new_n16014_;
  assign new_n16016_ = ~new_n16013_ & ~new_n16015_;
  assign new_n16017_ = ~\b[30]  & ~new_n16016_;
  assign new_n16018_ = ~new_n15384_ & new_n15760_;
  assign new_n16019_ = ~new_n15756_ & new_n16018_;
  assign new_n16020_ = ~new_n15757_ & ~new_n15760_;
  assign new_n16021_ = ~new_n16019_ & ~new_n16020_;
  assign new_n16022_ = \quotient[17]  & ~new_n16021_;
  assign new_n16023_ = ~new_n15374_ & ~new_n15863_;
  assign new_n16024_ = ~new_n15862_ & new_n16023_;
  assign new_n16025_ = ~new_n16022_ & ~new_n16024_;
  assign new_n16026_ = ~\b[29]  & ~new_n16025_;
  assign new_n16027_ = ~new_n15393_ & new_n15755_;
  assign new_n16028_ = ~new_n15751_ & new_n16027_;
  assign new_n16029_ = ~new_n15752_ & ~new_n15755_;
  assign new_n16030_ = ~new_n16028_ & ~new_n16029_;
  assign new_n16031_ = \quotient[17]  & ~new_n16030_;
  assign new_n16032_ = ~new_n15383_ & ~new_n15863_;
  assign new_n16033_ = ~new_n15862_ & new_n16032_;
  assign new_n16034_ = ~new_n16031_ & ~new_n16033_;
  assign new_n16035_ = ~\b[28]  & ~new_n16034_;
  assign new_n16036_ = ~new_n15402_ & new_n15750_;
  assign new_n16037_ = ~new_n15746_ & new_n16036_;
  assign new_n16038_ = ~new_n15747_ & ~new_n15750_;
  assign new_n16039_ = ~new_n16037_ & ~new_n16038_;
  assign new_n16040_ = \quotient[17]  & ~new_n16039_;
  assign new_n16041_ = ~new_n15392_ & ~new_n15863_;
  assign new_n16042_ = ~new_n15862_ & new_n16041_;
  assign new_n16043_ = ~new_n16040_ & ~new_n16042_;
  assign new_n16044_ = ~\b[27]  & ~new_n16043_;
  assign new_n16045_ = ~new_n15411_ & new_n15745_;
  assign new_n16046_ = ~new_n15741_ & new_n16045_;
  assign new_n16047_ = ~new_n15742_ & ~new_n15745_;
  assign new_n16048_ = ~new_n16046_ & ~new_n16047_;
  assign new_n16049_ = \quotient[17]  & ~new_n16048_;
  assign new_n16050_ = ~new_n15401_ & ~new_n15863_;
  assign new_n16051_ = ~new_n15862_ & new_n16050_;
  assign new_n16052_ = ~new_n16049_ & ~new_n16051_;
  assign new_n16053_ = ~\b[26]  & ~new_n16052_;
  assign new_n16054_ = ~new_n15420_ & new_n15740_;
  assign new_n16055_ = ~new_n15736_ & new_n16054_;
  assign new_n16056_ = ~new_n15737_ & ~new_n15740_;
  assign new_n16057_ = ~new_n16055_ & ~new_n16056_;
  assign new_n16058_ = \quotient[17]  & ~new_n16057_;
  assign new_n16059_ = ~new_n15410_ & ~new_n15863_;
  assign new_n16060_ = ~new_n15862_ & new_n16059_;
  assign new_n16061_ = ~new_n16058_ & ~new_n16060_;
  assign new_n16062_ = ~\b[25]  & ~new_n16061_;
  assign new_n16063_ = ~new_n15429_ & new_n15735_;
  assign new_n16064_ = ~new_n15731_ & new_n16063_;
  assign new_n16065_ = ~new_n15732_ & ~new_n15735_;
  assign new_n16066_ = ~new_n16064_ & ~new_n16065_;
  assign new_n16067_ = \quotient[17]  & ~new_n16066_;
  assign new_n16068_ = ~new_n15419_ & ~new_n15863_;
  assign new_n16069_ = ~new_n15862_ & new_n16068_;
  assign new_n16070_ = ~new_n16067_ & ~new_n16069_;
  assign new_n16071_ = ~\b[24]  & ~new_n16070_;
  assign new_n16072_ = ~new_n15438_ & new_n15730_;
  assign new_n16073_ = ~new_n15726_ & new_n16072_;
  assign new_n16074_ = ~new_n15727_ & ~new_n15730_;
  assign new_n16075_ = ~new_n16073_ & ~new_n16074_;
  assign new_n16076_ = \quotient[17]  & ~new_n16075_;
  assign new_n16077_ = ~new_n15428_ & ~new_n15863_;
  assign new_n16078_ = ~new_n15862_ & new_n16077_;
  assign new_n16079_ = ~new_n16076_ & ~new_n16078_;
  assign new_n16080_ = ~\b[23]  & ~new_n16079_;
  assign new_n16081_ = ~new_n15447_ & new_n15725_;
  assign new_n16082_ = ~new_n15721_ & new_n16081_;
  assign new_n16083_ = ~new_n15722_ & ~new_n15725_;
  assign new_n16084_ = ~new_n16082_ & ~new_n16083_;
  assign new_n16085_ = \quotient[17]  & ~new_n16084_;
  assign new_n16086_ = ~new_n15437_ & ~new_n15863_;
  assign new_n16087_ = ~new_n15862_ & new_n16086_;
  assign new_n16088_ = ~new_n16085_ & ~new_n16087_;
  assign new_n16089_ = ~\b[22]  & ~new_n16088_;
  assign new_n16090_ = ~new_n15456_ & new_n15720_;
  assign new_n16091_ = ~new_n15716_ & new_n16090_;
  assign new_n16092_ = ~new_n15717_ & ~new_n15720_;
  assign new_n16093_ = ~new_n16091_ & ~new_n16092_;
  assign new_n16094_ = \quotient[17]  & ~new_n16093_;
  assign new_n16095_ = ~new_n15446_ & ~new_n15863_;
  assign new_n16096_ = ~new_n15862_ & new_n16095_;
  assign new_n16097_ = ~new_n16094_ & ~new_n16096_;
  assign new_n16098_ = ~\b[21]  & ~new_n16097_;
  assign new_n16099_ = ~new_n15465_ & new_n15715_;
  assign new_n16100_ = ~new_n15711_ & new_n16099_;
  assign new_n16101_ = ~new_n15712_ & ~new_n15715_;
  assign new_n16102_ = ~new_n16100_ & ~new_n16101_;
  assign new_n16103_ = \quotient[17]  & ~new_n16102_;
  assign new_n16104_ = ~new_n15455_ & ~new_n15863_;
  assign new_n16105_ = ~new_n15862_ & new_n16104_;
  assign new_n16106_ = ~new_n16103_ & ~new_n16105_;
  assign new_n16107_ = ~\b[20]  & ~new_n16106_;
  assign new_n16108_ = ~new_n15474_ & new_n15710_;
  assign new_n16109_ = ~new_n15706_ & new_n16108_;
  assign new_n16110_ = ~new_n15707_ & ~new_n15710_;
  assign new_n16111_ = ~new_n16109_ & ~new_n16110_;
  assign new_n16112_ = \quotient[17]  & ~new_n16111_;
  assign new_n16113_ = ~new_n15464_ & ~new_n15863_;
  assign new_n16114_ = ~new_n15862_ & new_n16113_;
  assign new_n16115_ = ~new_n16112_ & ~new_n16114_;
  assign new_n16116_ = ~\b[19]  & ~new_n16115_;
  assign new_n16117_ = ~new_n15483_ & new_n15705_;
  assign new_n16118_ = ~new_n15701_ & new_n16117_;
  assign new_n16119_ = ~new_n15702_ & ~new_n15705_;
  assign new_n16120_ = ~new_n16118_ & ~new_n16119_;
  assign new_n16121_ = \quotient[17]  & ~new_n16120_;
  assign new_n16122_ = ~new_n15473_ & ~new_n15863_;
  assign new_n16123_ = ~new_n15862_ & new_n16122_;
  assign new_n16124_ = ~new_n16121_ & ~new_n16123_;
  assign new_n16125_ = ~\b[18]  & ~new_n16124_;
  assign new_n16126_ = ~new_n15492_ & new_n15700_;
  assign new_n16127_ = ~new_n15696_ & new_n16126_;
  assign new_n16128_ = ~new_n15697_ & ~new_n15700_;
  assign new_n16129_ = ~new_n16127_ & ~new_n16128_;
  assign new_n16130_ = \quotient[17]  & ~new_n16129_;
  assign new_n16131_ = ~new_n15482_ & ~new_n15863_;
  assign new_n16132_ = ~new_n15862_ & new_n16131_;
  assign new_n16133_ = ~new_n16130_ & ~new_n16132_;
  assign new_n16134_ = ~\b[17]  & ~new_n16133_;
  assign new_n16135_ = ~new_n15501_ & new_n15695_;
  assign new_n16136_ = ~new_n15691_ & new_n16135_;
  assign new_n16137_ = ~new_n15692_ & ~new_n15695_;
  assign new_n16138_ = ~new_n16136_ & ~new_n16137_;
  assign new_n16139_ = \quotient[17]  & ~new_n16138_;
  assign new_n16140_ = ~new_n15491_ & ~new_n15863_;
  assign new_n16141_ = ~new_n15862_ & new_n16140_;
  assign new_n16142_ = ~new_n16139_ & ~new_n16141_;
  assign new_n16143_ = ~\b[16]  & ~new_n16142_;
  assign new_n16144_ = ~new_n15510_ & new_n15690_;
  assign new_n16145_ = ~new_n15686_ & new_n16144_;
  assign new_n16146_ = ~new_n15687_ & ~new_n15690_;
  assign new_n16147_ = ~new_n16145_ & ~new_n16146_;
  assign new_n16148_ = \quotient[17]  & ~new_n16147_;
  assign new_n16149_ = ~new_n15500_ & ~new_n15863_;
  assign new_n16150_ = ~new_n15862_ & new_n16149_;
  assign new_n16151_ = ~new_n16148_ & ~new_n16150_;
  assign new_n16152_ = ~\b[15]  & ~new_n16151_;
  assign new_n16153_ = ~new_n15519_ & new_n15685_;
  assign new_n16154_ = ~new_n15681_ & new_n16153_;
  assign new_n16155_ = ~new_n15682_ & ~new_n15685_;
  assign new_n16156_ = ~new_n16154_ & ~new_n16155_;
  assign new_n16157_ = \quotient[17]  & ~new_n16156_;
  assign new_n16158_ = ~new_n15509_ & ~new_n15863_;
  assign new_n16159_ = ~new_n15862_ & new_n16158_;
  assign new_n16160_ = ~new_n16157_ & ~new_n16159_;
  assign new_n16161_ = ~\b[14]  & ~new_n16160_;
  assign new_n16162_ = ~new_n15528_ & new_n15680_;
  assign new_n16163_ = ~new_n15676_ & new_n16162_;
  assign new_n16164_ = ~new_n15677_ & ~new_n15680_;
  assign new_n16165_ = ~new_n16163_ & ~new_n16164_;
  assign new_n16166_ = \quotient[17]  & ~new_n16165_;
  assign new_n16167_ = ~new_n15518_ & ~new_n15863_;
  assign new_n16168_ = ~new_n15862_ & new_n16167_;
  assign new_n16169_ = ~new_n16166_ & ~new_n16168_;
  assign new_n16170_ = ~\b[13]  & ~new_n16169_;
  assign new_n16171_ = ~new_n15537_ & new_n15675_;
  assign new_n16172_ = ~new_n15671_ & new_n16171_;
  assign new_n16173_ = ~new_n15672_ & ~new_n15675_;
  assign new_n16174_ = ~new_n16172_ & ~new_n16173_;
  assign new_n16175_ = \quotient[17]  & ~new_n16174_;
  assign new_n16176_ = ~new_n15527_ & ~new_n15863_;
  assign new_n16177_ = ~new_n15862_ & new_n16176_;
  assign new_n16178_ = ~new_n16175_ & ~new_n16177_;
  assign new_n16179_ = ~\b[12]  & ~new_n16178_;
  assign new_n16180_ = ~new_n15546_ & new_n15670_;
  assign new_n16181_ = ~new_n15666_ & new_n16180_;
  assign new_n16182_ = ~new_n15667_ & ~new_n15670_;
  assign new_n16183_ = ~new_n16181_ & ~new_n16182_;
  assign new_n16184_ = \quotient[17]  & ~new_n16183_;
  assign new_n16185_ = ~new_n15536_ & ~new_n15863_;
  assign new_n16186_ = ~new_n15862_ & new_n16185_;
  assign new_n16187_ = ~new_n16184_ & ~new_n16186_;
  assign new_n16188_ = ~\b[11]  & ~new_n16187_;
  assign new_n16189_ = ~new_n15555_ & new_n15665_;
  assign new_n16190_ = ~new_n15661_ & new_n16189_;
  assign new_n16191_ = ~new_n15662_ & ~new_n15665_;
  assign new_n16192_ = ~new_n16190_ & ~new_n16191_;
  assign new_n16193_ = \quotient[17]  & ~new_n16192_;
  assign new_n16194_ = ~new_n15545_ & ~new_n15863_;
  assign new_n16195_ = ~new_n15862_ & new_n16194_;
  assign new_n16196_ = ~new_n16193_ & ~new_n16195_;
  assign new_n16197_ = ~\b[10]  & ~new_n16196_;
  assign new_n16198_ = ~new_n15564_ & new_n15660_;
  assign new_n16199_ = ~new_n15656_ & new_n16198_;
  assign new_n16200_ = ~new_n15657_ & ~new_n15660_;
  assign new_n16201_ = ~new_n16199_ & ~new_n16200_;
  assign new_n16202_ = \quotient[17]  & ~new_n16201_;
  assign new_n16203_ = ~new_n15554_ & ~new_n15863_;
  assign new_n16204_ = ~new_n15862_ & new_n16203_;
  assign new_n16205_ = ~new_n16202_ & ~new_n16204_;
  assign new_n16206_ = ~\b[9]  & ~new_n16205_;
  assign new_n16207_ = ~new_n15573_ & new_n15655_;
  assign new_n16208_ = ~new_n15651_ & new_n16207_;
  assign new_n16209_ = ~new_n15652_ & ~new_n15655_;
  assign new_n16210_ = ~new_n16208_ & ~new_n16209_;
  assign new_n16211_ = \quotient[17]  & ~new_n16210_;
  assign new_n16212_ = ~new_n15563_ & ~new_n15863_;
  assign new_n16213_ = ~new_n15862_ & new_n16212_;
  assign new_n16214_ = ~new_n16211_ & ~new_n16213_;
  assign new_n16215_ = ~\b[8]  & ~new_n16214_;
  assign new_n16216_ = ~new_n15582_ & new_n15650_;
  assign new_n16217_ = ~new_n15646_ & new_n16216_;
  assign new_n16218_ = ~new_n15647_ & ~new_n15650_;
  assign new_n16219_ = ~new_n16217_ & ~new_n16218_;
  assign new_n16220_ = \quotient[17]  & ~new_n16219_;
  assign new_n16221_ = ~new_n15572_ & ~new_n15863_;
  assign new_n16222_ = ~new_n15862_ & new_n16221_;
  assign new_n16223_ = ~new_n16220_ & ~new_n16222_;
  assign new_n16224_ = ~\b[7]  & ~new_n16223_;
  assign new_n16225_ = ~new_n15591_ & new_n15645_;
  assign new_n16226_ = ~new_n15641_ & new_n16225_;
  assign new_n16227_ = ~new_n15642_ & ~new_n15645_;
  assign new_n16228_ = ~new_n16226_ & ~new_n16227_;
  assign new_n16229_ = \quotient[17]  & ~new_n16228_;
  assign new_n16230_ = ~new_n15581_ & ~new_n15863_;
  assign new_n16231_ = ~new_n15862_ & new_n16230_;
  assign new_n16232_ = ~new_n16229_ & ~new_n16231_;
  assign new_n16233_ = ~\b[6]  & ~new_n16232_;
  assign new_n16234_ = ~new_n15600_ & new_n15640_;
  assign new_n16235_ = ~new_n15636_ & new_n16234_;
  assign new_n16236_ = ~new_n15637_ & ~new_n15640_;
  assign new_n16237_ = ~new_n16235_ & ~new_n16236_;
  assign new_n16238_ = \quotient[17]  & ~new_n16237_;
  assign new_n16239_ = ~new_n15590_ & ~new_n15863_;
  assign new_n16240_ = ~new_n15862_ & new_n16239_;
  assign new_n16241_ = ~new_n16238_ & ~new_n16240_;
  assign new_n16242_ = ~\b[5]  & ~new_n16241_;
  assign new_n16243_ = ~new_n15608_ & new_n15635_;
  assign new_n16244_ = ~new_n15631_ & new_n16243_;
  assign new_n16245_ = ~new_n15632_ & ~new_n15635_;
  assign new_n16246_ = ~new_n16244_ & ~new_n16245_;
  assign new_n16247_ = \quotient[17]  & ~new_n16246_;
  assign new_n16248_ = ~new_n15599_ & ~new_n15863_;
  assign new_n16249_ = ~new_n15862_ & new_n16248_;
  assign new_n16250_ = ~new_n16247_ & ~new_n16249_;
  assign new_n16251_ = ~\b[4]  & ~new_n16250_;
  assign new_n16252_ = ~new_n15626_ & new_n15630_;
  assign new_n16253_ = ~new_n15625_ & new_n16252_;
  assign new_n16254_ = ~new_n15627_ & ~new_n15630_;
  assign new_n16255_ = ~new_n16253_ & ~new_n16254_;
  assign new_n16256_ = \quotient[17]  & ~new_n16255_;
  assign new_n16257_ = ~new_n15607_ & ~new_n15863_;
  assign new_n16258_ = ~new_n15862_ & new_n16257_;
  assign new_n16259_ = ~new_n16256_ & ~new_n16258_;
  assign new_n16260_ = ~\b[3]  & ~new_n16259_;
  assign new_n16261_ = ~new_n15622_ & new_n15624_;
  assign new_n16262_ = ~new_n15620_ & new_n16261_;
  assign new_n16263_ = ~new_n15625_ & ~new_n16262_;
  assign new_n16264_ = \quotient[17]  & new_n16263_;
  assign new_n16265_ = ~new_n15619_ & ~new_n15863_;
  assign new_n16266_ = ~new_n15862_ & new_n16265_;
  assign new_n16267_ = ~new_n16264_ & ~new_n16266_;
  assign new_n16268_ = ~\b[2]  & ~new_n16267_;
  assign new_n16269_ = \b[0]  & \quotient[17] ;
  assign new_n16270_ = \a[17]  & ~new_n16269_;
  assign new_n16271_ = new_n15624_ & \quotient[17] ;
  assign new_n16272_ = ~new_n16270_ & ~new_n16271_;
  assign new_n16273_ = \b[1]  & ~new_n16272_;
  assign new_n16274_ = ~\b[1]  & ~new_n16271_;
  assign new_n16275_ = ~new_n16270_ & new_n16274_;
  assign new_n16276_ = ~new_n16273_ & ~new_n16275_;
  assign new_n16277_ = ~\a[16]  & \b[0] ;
  assign new_n16278_ = ~new_n16276_ & ~new_n16277_;
  assign new_n16279_ = ~\b[1]  & ~new_n16272_;
  assign new_n16280_ = ~new_n16278_ & ~new_n16279_;
  assign new_n16281_ = \b[2]  & ~new_n16266_;
  assign new_n16282_ = ~new_n16264_ & new_n16281_;
  assign new_n16283_ = ~new_n16268_ & ~new_n16282_;
  assign new_n16284_ = ~new_n16280_ & new_n16283_;
  assign new_n16285_ = ~new_n16268_ & ~new_n16284_;
  assign new_n16286_ = \b[3]  & ~new_n16258_;
  assign new_n16287_ = ~new_n16256_ & new_n16286_;
  assign new_n16288_ = ~new_n16260_ & ~new_n16287_;
  assign new_n16289_ = ~new_n16285_ & new_n16288_;
  assign new_n16290_ = ~new_n16260_ & ~new_n16289_;
  assign new_n16291_ = \b[4]  & ~new_n16249_;
  assign new_n16292_ = ~new_n16247_ & new_n16291_;
  assign new_n16293_ = ~new_n16251_ & ~new_n16292_;
  assign new_n16294_ = ~new_n16290_ & new_n16293_;
  assign new_n16295_ = ~new_n16251_ & ~new_n16294_;
  assign new_n16296_ = \b[5]  & ~new_n16240_;
  assign new_n16297_ = ~new_n16238_ & new_n16296_;
  assign new_n16298_ = ~new_n16242_ & ~new_n16297_;
  assign new_n16299_ = ~new_n16295_ & new_n16298_;
  assign new_n16300_ = ~new_n16242_ & ~new_n16299_;
  assign new_n16301_ = \b[6]  & ~new_n16231_;
  assign new_n16302_ = ~new_n16229_ & new_n16301_;
  assign new_n16303_ = ~new_n16233_ & ~new_n16302_;
  assign new_n16304_ = ~new_n16300_ & new_n16303_;
  assign new_n16305_ = ~new_n16233_ & ~new_n16304_;
  assign new_n16306_ = \b[7]  & ~new_n16222_;
  assign new_n16307_ = ~new_n16220_ & new_n16306_;
  assign new_n16308_ = ~new_n16224_ & ~new_n16307_;
  assign new_n16309_ = ~new_n16305_ & new_n16308_;
  assign new_n16310_ = ~new_n16224_ & ~new_n16309_;
  assign new_n16311_ = \b[8]  & ~new_n16213_;
  assign new_n16312_ = ~new_n16211_ & new_n16311_;
  assign new_n16313_ = ~new_n16215_ & ~new_n16312_;
  assign new_n16314_ = ~new_n16310_ & new_n16313_;
  assign new_n16315_ = ~new_n16215_ & ~new_n16314_;
  assign new_n16316_ = \b[9]  & ~new_n16204_;
  assign new_n16317_ = ~new_n16202_ & new_n16316_;
  assign new_n16318_ = ~new_n16206_ & ~new_n16317_;
  assign new_n16319_ = ~new_n16315_ & new_n16318_;
  assign new_n16320_ = ~new_n16206_ & ~new_n16319_;
  assign new_n16321_ = \b[10]  & ~new_n16195_;
  assign new_n16322_ = ~new_n16193_ & new_n16321_;
  assign new_n16323_ = ~new_n16197_ & ~new_n16322_;
  assign new_n16324_ = ~new_n16320_ & new_n16323_;
  assign new_n16325_ = ~new_n16197_ & ~new_n16324_;
  assign new_n16326_ = \b[11]  & ~new_n16186_;
  assign new_n16327_ = ~new_n16184_ & new_n16326_;
  assign new_n16328_ = ~new_n16188_ & ~new_n16327_;
  assign new_n16329_ = ~new_n16325_ & new_n16328_;
  assign new_n16330_ = ~new_n16188_ & ~new_n16329_;
  assign new_n16331_ = \b[12]  & ~new_n16177_;
  assign new_n16332_ = ~new_n16175_ & new_n16331_;
  assign new_n16333_ = ~new_n16179_ & ~new_n16332_;
  assign new_n16334_ = ~new_n16330_ & new_n16333_;
  assign new_n16335_ = ~new_n16179_ & ~new_n16334_;
  assign new_n16336_ = \b[13]  & ~new_n16168_;
  assign new_n16337_ = ~new_n16166_ & new_n16336_;
  assign new_n16338_ = ~new_n16170_ & ~new_n16337_;
  assign new_n16339_ = ~new_n16335_ & new_n16338_;
  assign new_n16340_ = ~new_n16170_ & ~new_n16339_;
  assign new_n16341_ = \b[14]  & ~new_n16159_;
  assign new_n16342_ = ~new_n16157_ & new_n16341_;
  assign new_n16343_ = ~new_n16161_ & ~new_n16342_;
  assign new_n16344_ = ~new_n16340_ & new_n16343_;
  assign new_n16345_ = ~new_n16161_ & ~new_n16344_;
  assign new_n16346_ = \b[15]  & ~new_n16150_;
  assign new_n16347_ = ~new_n16148_ & new_n16346_;
  assign new_n16348_ = ~new_n16152_ & ~new_n16347_;
  assign new_n16349_ = ~new_n16345_ & new_n16348_;
  assign new_n16350_ = ~new_n16152_ & ~new_n16349_;
  assign new_n16351_ = \b[16]  & ~new_n16141_;
  assign new_n16352_ = ~new_n16139_ & new_n16351_;
  assign new_n16353_ = ~new_n16143_ & ~new_n16352_;
  assign new_n16354_ = ~new_n16350_ & new_n16353_;
  assign new_n16355_ = ~new_n16143_ & ~new_n16354_;
  assign new_n16356_ = \b[17]  & ~new_n16132_;
  assign new_n16357_ = ~new_n16130_ & new_n16356_;
  assign new_n16358_ = ~new_n16134_ & ~new_n16357_;
  assign new_n16359_ = ~new_n16355_ & new_n16358_;
  assign new_n16360_ = ~new_n16134_ & ~new_n16359_;
  assign new_n16361_ = \b[18]  & ~new_n16123_;
  assign new_n16362_ = ~new_n16121_ & new_n16361_;
  assign new_n16363_ = ~new_n16125_ & ~new_n16362_;
  assign new_n16364_ = ~new_n16360_ & new_n16363_;
  assign new_n16365_ = ~new_n16125_ & ~new_n16364_;
  assign new_n16366_ = \b[19]  & ~new_n16114_;
  assign new_n16367_ = ~new_n16112_ & new_n16366_;
  assign new_n16368_ = ~new_n16116_ & ~new_n16367_;
  assign new_n16369_ = ~new_n16365_ & new_n16368_;
  assign new_n16370_ = ~new_n16116_ & ~new_n16369_;
  assign new_n16371_ = \b[20]  & ~new_n16105_;
  assign new_n16372_ = ~new_n16103_ & new_n16371_;
  assign new_n16373_ = ~new_n16107_ & ~new_n16372_;
  assign new_n16374_ = ~new_n16370_ & new_n16373_;
  assign new_n16375_ = ~new_n16107_ & ~new_n16374_;
  assign new_n16376_ = \b[21]  & ~new_n16096_;
  assign new_n16377_ = ~new_n16094_ & new_n16376_;
  assign new_n16378_ = ~new_n16098_ & ~new_n16377_;
  assign new_n16379_ = ~new_n16375_ & new_n16378_;
  assign new_n16380_ = ~new_n16098_ & ~new_n16379_;
  assign new_n16381_ = \b[22]  & ~new_n16087_;
  assign new_n16382_ = ~new_n16085_ & new_n16381_;
  assign new_n16383_ = ~new_n16089_ & ~new_n16382_;
  assign new_n16384_ = ~new_n16380_ & new_n16383_;
  assign new_n16385_ = ~new_n16089_ & ~new_n16384_;
  assign new_n16386_ = \b[23]  & ~new_n16078_;
  assign new_n16387_ = ~new_n16076_ & new_n16386_;
  assign new_n16388_ = ~new_n16080_ & ~new_n16387_;
  assign new_n16389_ = ~new_n16385_ & new_n16388_;
  assign new_n16390_ = ~new_n16080_ & ~new_n16389_;
  assign new_n16391_ = \b[24]  & ~new_n16069_;
  assign new_n16392_ = ~new_n16067_ & new_n16391_;
  assign new_n16393_ = ~new_n16071_ & ~new_n16392_;
  assign new_n16394_ = ~new_n16390_ & new_n16393_;
  assign new_n16395_ = ~new_n16071_ & ~new_n16394_;
  assign new_n16396_ = \b[25]  & ~new_n16060_;
  assign new_n16397_ = ~new_n16058_ & new_n16396_;
  assign new_n16398_ = ~new_n16062_ & ~new_n16397_;
  assign new_n16399_ = ~new_n16395_ & new_n16398_;
  assign new_n16400_ = ~new_n16062_ & ~new_n16399_;
  assign new_n16401_ = \b[26]  & ~new_n16051_;
  assign new_n16402_ = ~new_n16049_ & new_n16401_;
  assign new_n16403_ = ~new_n16053_ & ~new_n16402_;
  assign new_n16404_ = ~new_n16400_ & new_n16403_;
  assign new_n16405_ = ~new_n16053_ & ~new_n16404_;
  assign new_n16406_ = \b[27]  & ~new_n16042_;
  assign new_n16407_ = ~new_n16040_ & new_n16406_;
  assign new_n16408_ = ~new_n16044_ & ~new_n16407_;
  assign new_n16409_ = ~new_n16405_ & new_n16408_;
  assign new_n16410_ = ~new_n16044_ & ~new_n16409_;
  assign new_n16411_ = \b[28]  & ~new_n16033_;
  assign new_n16412_ = ~new_n16031_ & new_n16411_;
  assign new_n16413_ = ~new_n16035_ & ~new_n16412_;
  assign new_n16414_ = ~new_n16410_ & new_n16413_;
  assign new_n16415_ = ~new_n16035_ & ~new_n16414_;
  assign new_n16416_ = \b[29]  & ~new_n16024_;
  assign new_n16417_ = ~new_n16022_ & new_n16416_;
  assign new_n16418_ = ~new_n16026_ & ~new_n16417_;
  assign new_n16419_ = ~new_n16415_ & new_n16418_;
  assign new_n16420_ = ~new_n16026_ & ~new_n16419_;
  assign new_n16421_ = \b[30]  & ~new_n16015_;
  assign new_n16422_ = ~new_n16013_ & new_n16421_;
  assign new_n16423_ = ~new_n16017_ & ~new_n16422_;
  assign new_n16424_ = ~new_n16420_ & new_n16423_;
  assign new_n16425_ = ~new_n16017_ & ~new_n16424_;
  assign new_n16426_ = \b[31]  & ~new_n16006_;
  assign new_n16427_ = ~new_n16004_ & new_n16426_;
  assign new_n16428_ = ~new_n16008_ & ~new_n16427_;
  assign new_n16429_ = ~new_n16425_ & new_n16428_;
  assign new_n16430_ = ~new_n16008_ & ~new_n16429_;
  assign new_n16431_ = \b[32]  & ~new_n15997_;
  assign new_n16432_ = ~new_n15995_ & new_n16431_;
  assign new_n16433_ = ~new_n15999_ & ~new_n16432_;
  assign new_n16434_ = ~new_n16430_ & new_n16433_;
  assign new_n16435_ = ~new_n15999_ & ~new_n16434_;
  assign new_n16436_ = \b[33]  & ~new_n15988_;
  assign new_n16437_ = ~new_n15986_ & new_n16436_;
  assign new_n16438_ = ~new_n15990_ & ~new_n16437_;
  assign new_n16439_ = ~new_n16435_ & new_n16438_;
  assign new_n16440_ = ~new_n15990_ & ~new_n16439_;
  assign new_n16441_ = \b[34]  & ~new_n15979_;
  assign new_n16442_ = ~new_n15977_ & new_n16441_;
  assign new_n16443_ = ~new_n15981_ & ~new_n16442_;
  assign new_n16444_ = ~new_n16440_ & new_n16443_;
  assign new_n16445_ = ~new_n15981_ & ~new_n16444_;
  assign new_n16446_ = \b[35]  & ~new_n15970_;
  assign new_n16447_ = ~new_n15968_ & new_n16446_;
  assign new_n16448_ = ~new_n15972_ & ~new_n16447_;
  assign new_n16449_ = ~new_n16445_ & new_n16448_;
  assign new_n16450_ = ~new_n15972_ & ~new_n16449_;
  assign new_n16451_ = \b[36]  & ~new_n15961_;
  assign new_n16452_ = ~new_n15959_ & new_n16451_;
  assign new_n16453_ = ~new_n15963_ & ~new_n16452_;
  assign new_n16454_ = ~new_n16450_ & new_n16453_;
  assign new_n16455_ = ~new_n15963_ & ~new_n16454_;
  assign new_n16456_ = \b[37]  & ~new_n15952_;
  assign new_n16457_ = ~new_n15950_ & new_n16456_;
  assign new_n16458_ = ~new_n15954_ & ~new_n16457_;
  assign new_n16459_ = ~new_n16455_ & new_n16458_;
  assign new_n16460_ = ~new_n15954_ & ~new_n16459_;
  assign new_n16461_ = \b[38]  & ~new_n15943_;
  assign new_n16462_ = ~new_n15941_ & new_n16461_;
  assign new_n16463_ = ~new_n15945_ & ~new_n16462_;
  assign new_n16464_ = ~new_n16460_ & new_n16463_;
  assign new_n16465_ = ~new_n15945_ & ~new_n16464_;
  assign new_n16466_ = \b[39]  & ~new_n15934_;
  assign new_n16467_ = ~new_n15932_ & new_n16466_;
  assign new_n16468_ = ~new_n15936_ & ~new_n16467_;
  assign new_n16469_ = ~new_n16465_ & new_n16468_;
  assign new_n16470_ = ~new_n15936_ & ~new_n16469_;
  assign new_n16471_ = \b[40]  & ~new_n15925_;
  assign new_n16472_ = ~new_n15923_ & new_n16471_;
  assign new_n16473_ = ~new_n15927_ & ~new_n16472_;
  assign new_n16474_ = ~new_n16470_ & new_n16473_;
  assign new_n16475_ = ~new_n15927_ & ~new_n16474_;
  assign new_n16476_ = \b[41]  & ~new_n15916_;
  assign new_n16477_ = ~new_n15914_ & new_n16476_;
  assign new_n16478_ = ~new_n15918_ & ~new_n16477_;
  assign new_n16479_ = ~new_n16475_ & new_n16478_;
  assign new_n16480_ = ~new_n15918_ & ~new_n16479_;
  assign new_n16481_ = \b[42]  & ~new_n15907_;
  assign new_n16482_ = ~new_n15905_ & new_n16481_;
  assign new_n16483_ = ~new_n15909_ & ~new_n16482_;
  assign new_n16484_ = ~new_n16480_ & new_n16483_;
  assign new_n16485_ = ~new_n15909_ & ~new_n16484_;
  assign new_n16486_ = \b[43]  & ~new_n15898_;
  assign new_n16487_ = ~new_n15896_ & new_n16486_;
  assign new_n16488_ = ~new_n15900_ & ~new_n16487_;
  assign new_n16489_ = ~new_n16485_ & new_n16488_;
  assign new_n16490_ = ~new_n15900_ & ~new_n16489_;
  assign new_n16491_ = \b[44]  & ~new_n15889_;
  assign new_n16492_ = ~new_n15887_ & new_n16491_;
  assign new_n16493_ = ~new_n15891_ & ~new_n16492_;
  assign new_n16494_ = ~new_n16490_ & new_n16493_;
  assign new_n16495_ = ~new_n15891_ & ~new_n16494_;
  assign new_n16496_ = \b[45]  & ~new_n15880_;
  assign new_n16497_ = ~new_n15878_ & new_n16496_;
  assign new_n16498_ = ~new_n15882_ & ~new_n16497_;
  assign new_n16499_ = ~new_n16495_ & new_n16498_;
  assign new_n16500_ = ~new_n15882_ & ~new_n16499_;
  assign new_n16501_ = \b[46]  & ~new_n15871_;
  assign new_n16502_ = ~new_n15869_ & new_n16501_;
  assign new_n16503_ = ~new_n15873_ & ~new_n16502_;
  assign new_n16504_ = ~new_n16500_ & new_n16503_;
  assign new_n16505_ = ~new_n15873_ & ~new_n16504_;
  assign new_n16506_ = ~new_n15222_ & ~new_n15857_;
  assign new_n16507_ = ~new_n15855_ & new_n16506_;
  assign new_n16508_ = ~new_n15846_ & new_n16507_;
  assign new_n16509_ = ~new_n15855_ & ~new_n15857_;
  assign new_n16510_ = ~new_n15847_ & ~new_n16509_;
  assign new_n16511_ = ~new_n16508_ & ~new_n16510_;
  assign new_n16512_ = \quotient[17]  & ~new_n16511_;
  assign new_n16513_ = ~new_n15854_ & ~new_n15863_;
  assign new_n16514_ = ~new_n15862_ & new_n16513_;
  assign new_n16515_ = ~new_n16512_ & ~new_n16514_;
  assign new_n16516_ = ~\b[47]  & ~new_n16515_;
  assign new_n16517_ = \b[47]  & ~new_n16514_;
  assign new_n16518_ = ~new_n16512_ & new_n16517_;
  assign new_n16519_ = new_n338_ & ~new_n16518_;
  assign new_n16520_ = ~new_n16516_ & new_n16519_;
  assign new_n16521_ = ~new_n16505_ & new_n16520_;
  assign new_n16522_ = new_n15859_ & ~new_n16515_;
  assign \quotient[16]  = new_n16521_ | new_n16522_;
  assign new_n16524_ = ~new_n15882_ & new_n16503_;
  assign new_n16525_ = ~new_n16499_ & new_n16524_;
  assign new_n16526_ = ~new_n16500_ & ~new_n16503_;
  assign new_n16527_ = ~new_n16525_ & ~new_n16526_;
  assign new_n16528_ = \quotient[16]  & ~new_n16527_;
  assign new_n16529_ = ~new_n15872_ & ~new_n16522_;
  assign new_n16530_ = ~new_n16521_ & new_n16529_;
  assign new_n16531_ = ~new_n16528_ & ~new_n16530_;
  assign new_n16532_ = ~new_n15873_ & ~new_n16518_;
  assign new_n16533_ = ~new_n16516_ & new_n16532_;
  assign new_n16534_ = ~new_n16504_ & new_n16533_;
  assign new_n16535_ = ~new_n16516_ & ~new_n16518_;
  assign new_n16536_ = ~new_n16505_ & ~new_n16535_;
  assign new_n16537_ = ~new_n16534_ & ~new_n16536_;
  assign new_n16538_ = \quotient[16]  & ~new_n16537_;
  assign new_n16539_ = ~new_n16515_ & ~new_n16522_;
  assign new_n16540_ = ~new_n16521_ & new_n16539_;
  assign new_n16541_ = ~new_n16538_ & ~new_n16540_;
  assign new_n16542_ = ~\b[48]  & ~new_n16541_;
  assign new_n16543_ = ~\b[47]  & ~new_n16531_;
  assign new_n16544_ = ~new_n15891_ & new_n16498_;
  assign new_n16545_ = ~new_n16494_ & new_n16544_;
  assign new_n16546_ = ~new_n16495_ & ~new_n16498_;
  assign new_n16547_ = ~new_n16545_ & ~new_n16546_;
  assign new_n16548_ = \quotient[16]  & ~new_n16547_;
  assign new_n16549_ = ~new_n15881_ & ~new_n16522_;
  assign new_n16550_ = ~new_n16521_ & new_n16549_;
  assign new_n16551_ = ~new_n16548_ & ~new_n16550_;
  assign new_n16552_ = ~\b[46]  & ~new_n16551_;
  assign new_n16553_ = ~new_n15900_ & new_n16493_;
  assign new_n16554_ = ~new_n16489_ & new_n16553_;
  assign new_n16555_ = ~new_n16490_ & ~new_n16493_;
  assign new_n16556_ = ~new_n16554_ & ~new_n16555_;
  assign new_n16557_ = \quotient[16]  & ~new_n16556_;
  assign new_n16558_ = ~new_n15890_ & ~new_n16522_;
  assign new_n16559_ = ~new_n16521_ & new_n16558_;
  assign new_n16560_ = ~new_n16557_ & ~new_n16559_;
  assign new_n16561_ = ~\b[45]  & ~new_n16560_;
  assign new_n16562_ = ~new_n15909_ & new_n16488_;
  assign new_n16563_ = ~new_n16484_ & new_n16562_;
  assign new_n16564_ = ~new_n16485_ & ~new_n16488_;
  assign new_n16565_ = ~new_n16563_ & ~new_n16564_;
  assign new_n16566_ = \quotient[16]  & ~new_n16565_;
  assign new_n16567_ = ~new_n15899_ & ~new_n16522_;
  assign new_n16568_ = ~new_n16521_ & new_n16567_;
  assign new_n16569_ = ~new_n16566_ & ~new_n16568_;
  assign new_n16570_ = ~\b[44]  & ~new_n16569_;
  assign new_n16571_ = ~new_n15918_ & new_n16483_;
  assign new_n16572_ = ~new_n16479_ & new_n16571_;
  assign new_n16573_ = ~new_n16480_ & ~new_n16483_;
  assign new_n16574_ = ~new_n16572_ & ~new_n16573_;
  assign new_n16575_ = \quotient[16]  & ~new_n16574_;
  assign new_n16576_ = ~new_n15908_ & ~new_n16522_;
  assign new_n16577_ = ~new_n16521_ & new_n16576_;
  assign new_n16578_ = ~new_n16575_ & ~new_n16577_;
  assign new_n16579_ = ~\b[43]  & ~new_n16578_;
  assign new_n16580_ = ~new_n15927_ & new_n16478_;
  assign new_n16581_ = ~new_n16474_ & new_n16580_;
  assign new_n16582_ = ~new_n16475_ & ~new_n16478_;
  assign new_n16583_ = ~new_n16581_ & ~new_n16582_;
  assign new_n16584_ = \quotient[16]  & ~new_n16583_;
  assign new_n16585_ = ~new_n15917_ & ~new_n16522_;
  assign new_n16586_ = ~new_n16521_ & new_n16585_;
  assign new_n16587_ = ~new_n16584_ & ~new_n16586_;
  assign new_n16588_ = ~\b[42]  & ~new_n16587_;
  assign new_n16589_ = ~new_n15936_ & new_n16473_;
  assign new_n16590_ = ~new_n16469_ & new_n16589_;
  assign new_n16591_ = ~new_n16470_ & ~new_n16473_;
  assign new_n16592_ = ~new_n16590_ & ~new_n16591_;
  assign new_n16593_ = \quotient[16]  & ~new_n16592_;
  assign new_n16594_ = ~new_n15926_ & ~new_n16522_;
  assign new_n16595_ = ~new_n16521_ & new_n16594_;
  assign new_n16596_ = ~new_n16593_ & ~new_n16595_;
  assign new_n16597_ = ~\b[41]  & ~new_n16596_;
  assign new_n16598_ = ~new_n15945_ & new_n16468_;
  assign new_n16599_ = ~new_n16464_ & new_n16598_;
  assign new_n16600_ = ~new_n16465_ & ~new_n16468_;
  assign new_n16601_ = ~new_n16599_ & ~new_n16600_;
  assign new_n16602_ = \quotient[16]  & ~new_n16601_;
  assign new_n16603_ = ~new_n15935_ & ~new_n16522_;
  assign new_n16604_ = ~new_n16521_ & new_n16603_;
  assign new_n16605_ = ~new_n16602_ & ~new_n16604_;
  assign new_n16606_ = ~\b[40]  & ~new_n16605_;
  assign new_n16607_ = ~new_n15954_ & new_n16463_;
  assign new_n16608_ = ~new_n16459_ & new_n16607_;
  assign new_n16609_ = ~new_n16460_ & ~new_n16463_;
  assign new_n16610_ = ~new_n16608_ & ~new_n16609_;
  assign new_n16611_ = \quotient[16]  & ~new_n16610_;
  assign new_n16612_ = ~new_n15944_ & ~new_n16522_;
  assign new_n16613_ = ~new_n16521_ & new_n16612_;
  assign new_n16614_ = ~new_n16611_ & ~new_n16613_;
  assign new_n16615_ = ~\b[39]  & ~new_n16614_;
  assign new_n16616_ = ~new_n15963_ & new_n16458_;
  assign new_n16617_ = ~new_n16454_ & new_n16616_;
  assign new_n16618_ = ~new_n16455_ & ~new_n16458_;
  assign new_n16619_ = ~new_n16617_ & ~new_n16618_;
  assign new_n16620_ = \quotient[16]  & ~new_n16619_;
  assign new_n16621_ = ~new_n15953_ & ~new_n16522_;
  assign new_n16622_ = ~new_n16521_ & new_n16621_;
  assign new_n16623_ = ~new_n16620_ & ~new_n16622_;
  assign new_n16624_ = ~\b[38]  & ~new_n16623_;
  assign new_n16625_ = ~new_n15972_ & new_n16453_;
  assign new_n16626_ = ~new_n16449_ & new_n16625_;
  assign new_n16627_ = ~new_n16450_ & ~new_n16453_;
  assign new_n16628_ = ~new_n16626_ & ~new_n16627_;
  assign new_n16629_ = \quotient[16]  & ~new_n16628_;
  assign new_n16630_ = ~new_n15962_ & ~new_n16522_;
  assign new_n16631_ = ~new_n16521_ & new_n16630_;
  assign new_n16632_ = ~new_n16629_ & ~new_n16631_;
  assign new_n16633_ = ~\b[37]  & ~new_n16632_;
  assign new_n16634_ = ~new_n15981_ & new_n16448_;
  assign new_n16635_ = ~new_n16444_ & new_n16634_;
  assign new_n16636_ = ~new_n16445_ & ~new_n16448_;
  assign new_n16637_ = ~new_n16635_ & ~new_n16636_;
  assign new_n16638_ = \quotient[16]  & ~new_n16637_;
  assign new_n16639_ = ~new_n15971_ & ~new_n16522_;
  assign new_n16640_ = ~new_n16521_ & new_n16639_;
  assign new_n16641_ = ~new_n16638_ & ~new_n16640_;
  assign new_n16642_ = ~\b[36]  & ~new_n16641_;
  assign new_n16643_ = ~new_n15990_ & new_n16443_;
  assign new_n16644_ = ~new_n16439_ & new_n16643_;
  assign new_n16645_ = ~new_n16440_ & ~new_n16443_;
  assign new_n16646_ = ~new_n16644_ & ~new_n16645_;
  assign new_n16647_ = \quotient[16]  & ~new_n16646_;
  assign new_n16648_ = ~new_n15980_ & ~new_n16522_;
  assign new_n16649_ = ~new_n16521_ & new_n16648_;
  assign new_n16650_ = ~new_n16647_ & ~new_n16649_;
  assign new_n16651_ = ~\b[35]  & ~new_n16650_;
  assign new_n16652_ = ~new_n15999_ & new_n16438_;
  assign new_n16653_ = ~new_n16434_ & new_n16652_;
  assign new_n16654_ = ~new_n16435_ & ~new_n16438_;
  assign new_n16655_ = ~new_n16653_ & ~new_n16654_;
  assign new_n16656_ = \quotient[16]  & ~new_n16655_;
  assign new_n16657_ = ~new_n15989_ & ~new_n16522_;
  assign new_n16658_ = ~new_n16521_ & new_n16657_;
  assign new_n16659_ = ~new_n16656_ & ~new_n16658_;
  assign new_n16660_ = ~\b[34]  & ~new_n16659_;
  assign new_n16661_ = ~new_n16008_ & new_n16433_;
  assign new_n16662_ = ~new_n16429_ & new_n16661_;
  assign new_n16663_ = ~new_n16430_ & ~new_n16433_;
  assign new_n16664_ = ~new_n16662_ & ~new_n16663_;
  assign new_n16665_ = \quotient[16]  & ~new_n16664_;
  assign new_n16666_ = ~new_n15998_ & ~new_n16522_;
  assign new_n16667_ = ~new_n16521_ & new_n16666_;
  assign new_n16668_ = ~new_n16665_ & ~new_n16667_;
  assign new_n16669_ = ~\b[33]  & ~new_n16668_;
  assign new_n16670_ = ~new_n16017_ & new_n16428_;
  assign new_n16671_ = ~new_n16424_ & new_n16670_;
  assign new_n16672_ = ~new_n16425_ & ~new_n16428_;
  assign new_n16673_ = ~new_n16671_ & ~new_n16672_;
  assign new_n16674_ = \quotient[16]  & ~new_n16673_;
  assign new_n16675_ = ~new_n16007_ & ~new_n16522_;
  assign new_n16676_ = ~new_n16521_ & new_n16675_;
  assign new_n16677_ = ~new_n16674_ & ~new_n16676_;
  assign new_n16678_ = ~\b[32]  & ~new_n16677_;
  assign new_n16679_ = ~new_n16026_ & new_n16423_;
  assign new_n16680_ = ~new_n16419_ & new_n16679_;
  assign new_n16681_ = ~new_n16420_ & ~new_n16423_;
  assign new_n16682_ = ~new_n16680_ & ~new_n16681_;
  assign new_n16683_ = \quotient[16]  & ~new_n16682_;
  assign new_n16684_ = ~new_n16016_ & ~new_n16522_;
  assign new_n16685_ = ~new_n16521_ & new_n16684_;
  assign new_n16686_ = ~new_n16683_ & ~new_n16685_;
  assign new_n16687_ = ~\b[31]  & ~new_n16686_;
  assign new_n16688_ = ~new_n16035_ & new_n16418_;
  assign new_n16689_ = ~new_n16414_ & new_n16688_;
  assign new_n16690_ = ~new_n16415_ & ~new_n16418_;
  assign new_n16691_ = ~new_n16689_ & ~new_n16690_;
  assign new_n16692_ = \quotient[16]  & ~new_n16691_;
  assign new_n16693_ = ~new_n16025_ & ~new_n16522_;
  assign new_n16694_ = ~new_n16521_ & new_n16693_;
  assign new_n16695_ = ~new_n16692_ & ~new_n16694_;
  assign new_n16696_ = ~\b[30]  & ~new_n16695_;
  assign new_n16697_ = ~new_n16044_ & new_n16413_;
  assign new_n16698_ = ~new_n16409_ & new_n16697_;
  assign new_n16699_ = ~new_n16410_ & ~new_n16413_;
  assign new_n16700_ = ~new_n16698_ & ~new_n16699_;
  assign new_n16701_ = \quotient[16]  & ~new_n16700_;
  assign new_n16702_ = ~new_n16034_ & ~new_n16522_;
  assign new_n16703_ = ~new_n16521_ & new_n16702_;
  assign new_n16704_ = ~new_n16701_ & ~new_n16703_;
  assign new_n16705_ = ~\b[29]  & ~new_n16704_;
  assign new_n16706_ = ~new_n16053_ & new_n16408_;
  assign new_n16707_ = ~new_n16404_ & new_n16706_;
  assign new_n16708_ = ~new_n16405_ & ~new_n16408_;
  assign new_n16709_ = ~new_n16707_ & ~new_n16708_;
  assign new_n16710_ = \quotient[16]  & ~new_n16709_;
  assign new_n16711_ = ~new_n16043_ & ~new_n16522_;
  assign new_n16712_ = ~new_n16521_ & new_n16711_;
  assign new_n16713_ = ~new_n16710_ & ~new_n16712_;
  assign new_n16714_ = ~\b[28]  & ~new_n16713_;
  assign new_n16715_ = ~new_n16062_ & new_n16403_;
  assign new_n16716_ = ~new_n16399_ & new_n16715_;
  assign new_n16717_ = ~new_n16400_ & ~new_n16403_;
  assign new_n16718_ = ~new_n16716_ & ~new_n16717_;
  assign new_n16719_ = \quotient[16]  & ~new_n16718_;
  assign new_n16720_ = ~new_n16052_ & ~new_n16522_;
  assign new_n16721_ = ~new_n16521_ & new_n16720_;
  assign new_n16722_ = ~new_n16719_ & ~new_n16721_;
  assign new_n16723_ = ~\b[27]  & ~new_n16722_;
  assign new_n16724_ = ~new_n16071_ & new_n16398_;
  assign new_n16725_ = ~new_n16394_ & new_n16724_;
  assign new_n16726_ = ~new_n16395_ & ~new_n16398_;
  assign new_n16727_ = ~new_n16725_ & ~new_n16726_;
  assign new_n16728_ = \quotient[16]  & ~new_n16727_;
  assign new_n16729_ = ~new_n16061_ & ~new_n16522_;
  assign new_n16730_ = ~new_n16521_ & new_n16729_;
  assign new_n16731_ = ~new_n16728_ & ~new_n16730_;
  assign new_n16732_ = ~\b[26]  & ~new_n16731_;
  assign new_n16733_ = ~new_n16080_ & new_n16393_;
  assign new_n16734_ = ~new_n16389_ & new_n16733_;
  assign new_n16735_ = ~new_n16390_ & ~new_n16393_;
  assign new_n16736_ = ~new_n16734_ & ~new_n16735_;
  assign new_n16737_ = \quotient[16]  & ~new_n16736_;
  assign new_n16738_ = ~new_n16070_ & ~new_n16522_;
  assign new_n16739_ = ~new_n16521_ & new_n16738_;
  assign new_n16740_ = ~new_n16737_ & ~new_n16739_;
  assign new_n16741_ = ~\b[25]  & ~new_n16740_;
  assign new_n16742_ = ~new_n16089_ & new_n16388_;
  assign new_n16743_ = ~new_n16384_ & new_n16742_;
  assign new_n16744_ = ~new_n16385_ & ~new_n16388_;
  assign new_n16745_ = ~new_n16743_ & ~new_n16744_;
  assign new_n16746_ = \quotient[16]  & ~new_n16745_;
  assign new_n16747_ = ~new_n16079_ & ~new_n16522_;
  assign new_n16748_ = ~new_n16521_ & new_n16747_;
  assign new_n16749_ = ~new_n16746_ & ~new_n16748_;
  assign new_n16750_ = ~\b[24]  & ~new_n16749_;
  assign new_n16751_ = ~new_n16098_ & new_n16383_;
  assign new_n16752_ = ~new_n16379_ & new_n16751_;
  assign new_n16753_ = ~new_n16380_ & ~new_n16383_;
  assign new_n16754_ = ~new_n16752_ & ~new_n16753_;
  assign new_n16755_ = \quotient[16]  & ~new_n16754_;
  assign new_n16756_ = ~new_n16088_ & ~new_n16522_;
  assign new_n16757_ = ~new_n16521_ & new_n16756_;
  assign new_n16758_ = ~new_n16755_ & ~new_n16757_;
  assign new_n16759_ = ~\b[23]  & ~new_n16758_;
  assign new_n16760_ = ~new_n16107_ & new_n16378_;
  assign new_n16761_ = ~new_n16374_ & new_n16760_;
  assign new_n16762_ = ~new_n16375_ & ~new_n16378_;
  assign new_n16763_ = ~new_n16761_ & ~new_n16762_;
  assign new_n16764_ = \quotient[16]  & ~new_n16763_;
  assign new_n16765_ = ~new_n16097_ & ~new_n16522_;
  assign new_n16766_ = ~new_n16521_ & new_n16765_;
  assign new_n16767_ = ~new_n16764_ & ~new_n16766_;
  assign new_n16768_ = ~\b[22]  & ~new_n16767_;
  assign new_n16769_ = ~new_n16116_ & new_n16373_;
  assign new_n16770_ = ~new_n16369_ & new_n16769_;
  assign new_n16771_ = ~new_n16370_ & ~new_n16373_;
  assign new_n16772_ = ~new_n16770_ & ~new_n16771_;
  assign new_n16773_ = \quotient[16]  & ~new_n16772_;
  assign new_n16774_ = ~new_n16106_ & ~new_n16522_;
  assign new_n16775_ = ~new_n16521_ & new_n16774_;
  assign new_n16776_ = ~new_n16773_ & ~new_n16775_;
  assign new_n16777_ = ~\b[21]  & ~new_n16776_;
  assign new_n16778_ = ~new_n16125_ & new_n16368_;
  assign new_n16779_ = ~new_n16364_ & new_n16778_;
  assign new_n16780_ = ~new_n16365_ & ~new_n16368_;
  assign new_n16781_ = ~new_n16779_ & ~new_n16780_;
  assign new_n16782_ = \quotient[16]  & ~new_n16781_;
  assign new_n16783_ = ~new_n16115_ & ~new_n16522_;
  assign new_n16784_ = ~new_n16521_ & new_n16783_;
  assign new_n16785_ = ~new_n16782_ & ~new_n16784_;
  assign new_n16786_ = ~\b[20]  & ~new_n16785_;
  assign new_n16787_ = ~new_n16134_ & new_n16363_;
  assign new_n16788_ = ~new_n16359_ & new_n16787_;
  assign new_n16789_ = ~new_n16360_ & ~new_n16363_;
  assign new_n16790_ = ~new_n16788_ & ~new_n16789_;
  assign new_n16791_ = \quotient[16]  & ~new_n16790_;
  assign new_n16792_ = ~new_n16124_ & ~new_n16522_;
  assign new_n16793_ = ~new_n16521_ & new_n16792_;
  assign new_n16794_ = ~new_n16791_ & ~new_n16793_;
  assign new_n16795_ = ~\b[19]  & ~new_n16794_;
  assign new_n16796_ = ~new_n16143_ & new_n16358_;
  assign new_n16797_ = ~new_n16354_ & new_n16796_;
  assign new_n16798_ = ~new_n16355_ & ~new_n16358_;
  assign new_n16799_ = ~new_n16797_ & ~new_n16798_;
  assign new_n16800_ = \quotient[16]  & ~new_n16799_;
  assign new_n16801_ = ~new_n16133_ & ~new_n16522_;
  assign new_n16802_ = ~new_n16521_ & new_n16801_;
  assign new_n16803_ = ~new_n16800_ & ~new_n16802_;
  assign new_n16804_ = ~\b[18]  & ~new_n16803_;
  assign new_n16805_ = ~new_n16152_ & new_n16353_;
  assign new_n16806_ = ~new_n16349_ & new_n16805_;
  assign new_n16807_ = ~new_n16350_ & ~new_n16353_;
  assign new_n16808_ = ~new_n16806_ & ~new_n16807_;
  assign new_n16809_ = \quotient[16]  & ~new_n16808_;
  assign new_n16810_ = ~new_n16142_ & ~new_n16522_;
  assign new_n16811_ = ~new_n16521_ & new_n16810_;
  assign new_n16812_ = ~new_n16809_ & ~new_n16811_;
  assign new_n16813_ = ~\b[17]  & ~new_n16812_;
  assign new_n16814_ = ~new_n16161_ & new_n16348_;
  assign new_n16815_ = ~new_n16344_ & new_n16814_;
  assign new_n16816_ = ~new_n16345_ & ~new_n16348_;
  assign new_n16817_ = ~new_n16815_ & ~new_n16816_;
  assign new_n16818_ = \quotient[16]  & ~new_n16817_;
  assign new_n16819_ = ~new_n16151_ & ~new_n16522_;
  assign new_n16820_ = ~new_n16521_ & new_n16819_;
  assign new_n16821_ = ~new_n16818_ & ~new_n16820_;
  assign new_n16822_ = ~\b[16]  & ~new_n16821_;
  assign new_n16823_ = ~new_n16170_ & new_n16343_;
  assign new_n16824_ = ~new_n16339_ & new_n16823_;
  assign new_n16825_ = ~new_n16340_ & ~new_n16343_;
  assign new_n16826_ = ~new_n16824_ & ~new_n16825_;
  assign new_n16827_ = \quotient[16]  & ~new_n16826_;
  assign new_n16828_ = ~new_n16160_ & ~new_n16522_;
  assign new_n16829_ = ~new_n16521_ & new_n16828_;
  assign new_n16830_ = ~new_n16827_ & ~new_n16829_;
  assign new_n16831_ = ~\b[15]  & ~new_n16830_;
  assign new_n16832_ = ~new_n16179_ & new_n16338_;
  assign new_n16833_ = ~new_n16334_ & new_n16832_;
  assign new_n16834_ = ~new_n16335_ & ~new_n16338_;
  assign new_n16835_ = ~new_n16833_ & ~new_n16834_;
  assign new_n16836_ = \quotient[16]  & ~new_n16835_;
  assign new_n16837_ = ~new_n16169_ & ~new_n16522_;
  assign new_n16838_ = ~new_n16521_ & new_n16837_;
  assign new_n16839_ = ~new_n16836_ & ~new_n16838_;
  assign new_n16840_ = ~\b[14]  & ~new_n16839_;
  assign new_n16841_ = ~new_n16188_ & new_n16333_;
  assign new_n16842_ = ~new_n16329_ & new_n16841_;
  assign new_n16843_ = ~new_n16330_ & ~new_n16333_;
  assign new_n16844_ = ~new_n16842_ & ~new_n16843_;
  assign new_n16845_ = \quotient[16]  & ~new_n16844_;
  assign new_n16846_ = ~new_n16178_ & ~new_n16522_;
  assign new_n16847_ = ~new_n16521_ & new_n16846_;
  assign new_n16848_ = ~new_n16845_ & ~new_n16847_;
  assign new_n16849_ = ~\b[13]  & ~new_n16848_;
  assign new_n16850_ = ~new_n16197_ & new_n16328_;
  assign new_n16851_ = ~new_n16324_ & new_n16850_;
  assign new_n16852_ = ~new_n16325_ & ~new_n16328_;
  assign new_n16853_ = ~new_n16851_ & ~new_n16852_;
  assign new_n16854_ = \quotient[16]  & ~new_n16853_;
  assign new_n16855_ = ~new_n16187_ & ~new_n16522_;
  assign new_n16856_ = ~new_n16521_ & new_n16855_;
  assign new_n16857_ = ~new_n16854_ & ~new_n16856_;
  assign new_n16858_ = ~\b[12]  & ~new_n16857_;
  assign new_n16859_ = ~new_n16206_ & new_n16323_;
  assign new_n16860_ = ~new_n16319_ & new_n16859_;
  assign new_n16861_ = ~new_n16320_ & ~new_n16323_;
  assign new_n16862_ = ~new_n16860_ & ~new_n16861_;
  assign new_n16863_ = \quotient[16]  & ~new_n16862_;
  assign new_n16864_ = ~new_n16196_ & ~new_n16522_;
  assign new_n16865_ = ~new_n16521_ & new_n16864_;
  assign new_n16866_ = ~new_n16863_ & ~new_n16865_;
  assign new_n16867_ = ~\b[11]  & ~new_n16866_;
  assign new_n16868_ = ~new_n16215_ & new_n16318_;
  assign new_n16869_ = ~new_n16314_ & new_n16868_;
  assign new_n16870_ = ~new_n16315_ & ~new_n16318_;
  assign new_n16871_ = ~new_n16869_ & ~new_n16870_;
  assign new_n16872_ = \quotient[16]  & ~new_n16871_;
  assign new_n16873_ = ~new_n16205_ & ~new_n16522_;
  assign new_n16874_ = ~new_n16521_ & new_n16873_;
  assign new_n16875_ = ~new_n16872_ & ~new_n16874_;
  assign new_n16876_ = ~\b[10]  & ~new_n16875_;
  assign new_n16877_ = ~new_n16224_ & new_n16313_;
  assign new_n16878_ = ~new_n16309_ & new_n16877_;
  assign new_n16879_ = ~new_n16310_ & ~new_n16313_;
  assign new_n16880_ = ~new_n16878_ & ~new_n16879_;
  assign new_n16881_ = \quotient[16]  & ~new_n16880_;
  assign new_n16882_ = ~new_n16214_ & ~new_n16522_;
  assign new_n16883_ = ~new_n16521_ & new_n16882_;
  assign new_n16884_ = ~new_n16881_ & ~new_n16883_;
  assign new_n16885_ = ~\b[9]  & ~new_n16884_;
  assign new_n16886_ = ~new_n16233_ & new_n16308_;
  assign new_n16887_ = ~new_n16304_ & new_n16886_;
  assign new_n16888_ = ~new_n16305_ & ~new_n16308_;
  assign new_n16889_ = ~new_n16887_ & ~new_n16888_;
  assign new_n16890_ = \quotient[16]  & ~new_n16889_;
  assign new_n16891_ = ~new_n16223_ & ~new_n16522_;
  assign new_n16892_ = ~new_n16521_ & new_n16891_;
  assign new_n16893_ = ~new_n16890_ & ~new_n16892_;
  assign new_n16894_ = ~\b[8]  & ~new_n16893_;
  assign new_n16895_ = ~new_n16242_ & new_n16303_;
  assign new_n16896_ = ~new_n16299_ & new_n16895_;
  assign new_n16897_ = ~new_n16300_ & ~new_n16303_;
  assign new_n16898_ = ~new_n16896_ & ~new_n16897_;
  assign new_n16899_ = \quotient[16]  & ~new_n16898_;
  assign new_n16900_ = ~new_n16232_ & ~new_n16522_;
  assign new_n16901_ = ~new_n16521_ & new_n16900_;
  assign new_n16902_ = ~new_n16899_ & ~new_n16901_;
  assign new_n16903_ = ~\b[7]  & ~new_n16902_;
  assign new_n16904_ = ~new_n16251_ & new_n16298_;
  assign new_n16905_ = ~new_n16294_ & new_n16904_;
  assign new_n16906_ = ~new_n16295_ & ~new_n16298_;
  assign new_n16907_ = ~new_n16905_ & ~new_n16906_;
  assign new_n16908_ = \quotient[16]  & ~new_n16907_;
  assign new_n16909_ = ~new_n16241_ & ~new_n16522_;
  assign new_n16910_ = ~new_n16521_ & new_n16909_;
  assign new_n16911_ = ~new_n16908_ & ~new_n16910_;
  assign new_n16912_ = ~\b[6]  & ~new_n16911_;
  assign new_n16913_ = ~new_n16260_ & new_n16293_;
  assign new_n16914_ = ~new_n16289_ & new_n16913_;
  assign new_n16915_ = ~new_n16290_ & ~new_n16293_;
  assign new_n16916_ = ~new_n16914_ & ~new_n16915_;
  assign new_n16917_ = \quotient[16]  & ~new_n16916_;
  assign new_n16918_ = ~new_n16250_ & ~new_n16522_;
  assign new_n16919_ = ~new_n16521_ & new_n16918_;
  assign new_n16920_ = ~new_n16917_ & ~new_n16919_;
  assign new_n16921_ = ~\b[5]  & ~new_n16920_;
  assign new_n16922_ = ~new_n16268_ & new_n16288_;
  assign new_n16923_ = ~new_n16284_ & new_n16922_;
  assign new_n16924_ = ~new_n16285_ & ~new_n16288_;
  assign new_n16925_ = ~new_n16923_ & ~new_n16924_;
  assign new_n16926_ = \quotient[16]  & ~new_n16925_;
  assign new_n16927_ = ~new_n16259_ & ~new_n16522_;
  assign new_n16928_ = ~new_n16521_ & new_n16927_;
  assign new_n16929_ = ~new_n16926_ & ~new_n16928_;
  assign new_n16930_ = ~\b[4]  & ~new_n16929_;
  assign new_n16931_ = ~new_n16279_ & new_n16283_;
  assign new_n16932_ = ~new_n16278_ & new_n16931_;
  assign new_n16933_ = ~new_n16280_ & ~new_n16283_;
  assign new_n16934_ = ~new_n16932_ & ~new_n16933_;
  assign new_n16935_ = \quotient[16]  & ~new_n16934_;
  assign new_n16936_ = ~new_n16267_ & ~new_n16522_;
  assign new_n16937_ = ~new_n16521_ & new_n16936_;
  assign new_n16938_ = ~new_n16935_ & ~new_n16937_;
  assign new_n16939_ = ~\b[3]  & ~new_n16938_;
  assign new_n16940_ = ~new_n16275_ & new_n16277_;
  assign new_n16941_ = ~new_n16273_ & new_n16940_;
  assign new_n16942_ = ~new_n16278_ & ~new_n16941_;
  assign new_n16943_ = \quotient[16]  & new_n16942_;
  assign new_n16944_ = ~new_n16272_ & ~new_n16522_;
  assign new_n16945_ = ~new_n16521_ & new_n16944_;
  assign new_n16946_ = ~new_n16943_ & ~new_n16945_;
  assign new_n16947_ = ~\b[2]  & ~new_n16946_;
  assign new_n16948_ = \b[0]  & \quotient[16] ;
  assign new_n16949_ = \a[16]  & ~new_n16948_;
  assign new_n16950_ = new_n16277_ & \quotient[16] ;
  assign new_n16951_ = ~new_n16949_ & ~new_n16950_;
  assign new_n16952_ = \b[1]  & ~new_n16951_;
  assign new_n16953_ = ~\b[1]  & ~new_n16950_;
  assign new_n16954_ = ~new_n16949_ & new_n16953_;
  assign new_n16955_ = ~new_n16952_ & ~new_n16954_;
  assign new_n16956_ = ~\a[15]  & \b[0] ;
  assign new_n16957_ = ~new_n16955_ & ~new_n16956_;
  assign new_n16958_ = ~\b[1]  & ~new_n16951_;
  assign new_n16959_ = ~new_n16957_ & ~new_n16958_;
  assign new_n16960_ = \b[2]  & ~new_n16945_;
  assign new_n16961_ = ~new_n16943_ & new_n16960_;
  assign new_n16962_ = ~new_n16947_ & ~new_n16961_;
  assign new_n16963_ = ~new_n16959_ & new_n16962_;
  assign new_n16964_ = ~new_n16947_ & ~new_n16963_;
  assign new_n16965_ = \b[3]  & ~new_n16937_;
  assign new_n16966_ = ~new_n16935_ & new_n16965_;
  assign new_n16967_ = ~new_n16939_ & ~new_n16966_;
  assign new_n16968_ = ~new_n16964_ & new_n16967_;
  assign new_n16969_ = ~new_n16939_ & ~new_n16968_;
  assign new_n16970_ = \b[4]  & ~new_n16928_;
  assign new_n16971_ = ~new_n16926_ & new_n16970_;
  assign new_n16972_ = ~new_n16930_ & ~new_n16971_;
  assign new_n16973_ = ~new_n16969_ & new_n16972_;
  assign new_n16974_ = ~new_n16930_ & ~new_n16973_;
  assign new_n16975_ = \b[5]  & ~new_n16919_;
  assign new_n16976_ = ~new_n16917_ & new_n16975_;
  assign new_n16977_ = ~new_n16921_ & ~new_n16976_;
  assign new_n16978_ = ~new_n16974_ & new_n16977_;
  assign new_n16979_ = ~new_n16921_ & ~new_n16978_;
  assign new_n16980_ = \b[6]  & ~new_n16910_;
  assign new_n16981_ = ~new_n16908_ & new_n16980_;
  assign new_n16982_ = ~new_n16912_ & ~new_n16981_;
  assign new_n16983_ = ~new_n16979_ & new_n16982_;
  assign new_n16984_ = ~new_n16912_ & ~new_n16983_;
  assign new_n16985_ = \b[7]  & ~new_n16901_;
  assign new_n16986_ = ~new_n16899_ & new_n16985_;
  assign new_n16987_ = ~new_n16903_ & ~new_n16986_;
  assign new_n16988_ = ~new_n16984_ & new_n16987_;
  assign new_n16989_ = ~new_n16903_ & ~new_n16988_;
  assign new_n16990_ = \b[8]  & ~new_n16892_;
  assign new_n16991_ = ~new_n16890_ & new_n16990_;
  assign new_n16992_ = ~new_n16894_ & ~new_n16991_;
  assign new_n16993_ = ~new_n16989_ & new_n16992_;
  assign new_n16994_ = ~new_n16894_ & ~new_n16993_;
  assign new_n16995_ = \b[9]  & ~new_n16883_;
  assign new_n16996_ = ~new_n16881_ & new_n16995_;
  assign new_n16997_ = ~new_n16885_ & ~new_n16996_;
  assign new_n16998_ = ~new_n16994_ & new_n16997_;
  assign new_n16999_ = ~new_n16885_ & ~new_n16998_;
  assign new_n17000_ = \b[10]  & ~new_n16874_;
  assign new_n17001_ = ~new_n16872_ & new_n17000_;
  assign new_n17002_ = ~new_n16876_ & ~new_n17001_;
  assign new_n17003_ = ~new_n16999_ & new_n17002_;
  assign new_n17004_ = ~new_n16876_ & ~new_n17003_;
  assign new_n17005_ = \b[11]  & ~new_n16865_;
  assign new_n17006_ = ~new_n16863_ & new_n17005_;
  assign new_n17007_ = ~new_n16867_ & ~new_n17006_;
  assign new_n17008_ = ~new_n17004_ & new_n17007_;
  assign new_n17009_ = ~new_n16867_ & ~new_n17008_;
  assign new_n17010_ = \b[12]  & ~new_n16856_;
  assign new_n17011_ = ~new_n16854_ & new_n17010_;
  assign new_n17012_ = ~new_n16858_ & ~new_n17011_;
  assign new_n17013_ = ~new_n17009_ & new_n17012_;
  assign new_n17014_ = ~new_n16858_ & ~new_n17013_;
  assign new_n17015_ = \b[13]  & ~new_n16847_;
  assign new_n17016_ = ~new_n16845_ & new_n17015_;
  assign new_n17017_ = ~new_n16849_ & ~new_n17016_;
  assign new_n17018_ = ~new_n17014_ & new_n17017_;
  assign new_n17019_ = ~new_n16849_ & ~new_n17018_;
  assign new_n17020_ = \b[14]  & ~new_n16838_;
  assign new_n17021_ = ~new_n16836_ & new_n17020_;
  assign new_n17022_ = ~new_n16840_ & ~new_n17021_;
  assign new_n17023_ = ~new_n17019_ & new_n17022_;
  assign new_n17024_ = ~new_n16840_ & ~new_n17023_;
  assign new_n17025_ = \b[15]  & ~new_n16829_;
  assign new_n17026_ = ~new_n16827_ & new_n17025_;
  assign new_n17027_ = ~new_n16831_ & ~new_n17026_;
  assign new_n17028_ = ~new_n17024_ & new_n17027_;
  assign new_n17029_ = ~new_n16831_ & ~new_n17028_;
  assign new_n17030_ = \b[16]  & ~new_n16820_;
  assign new_n17031_ = ~new_n16818_ & new_n17030_;
  assign new_n17032_ = ~new_n16822_ & ~new_n17031_;
  assign new_n17033_ = ~new_n17029_ & new_n17032_;
  assign new_n17034_ = ~new_n16822_ & ~new_n17033_;
  assign new_n17035_ = \b[17]  & ~new_n16811_;
  assign new_n17036_ = ~new_n16809_ & new_n17035_;
  assign new_n17037_ = ~new_n16813_ & ~new_n17036_;
  assign new_n17038_ = ~new_n17034_ & new_n17037_;
  assign new_n17039_ = ~new_n16813_ & ~new_n17038_;
  assign new_n17040_ = \b[18]  & ~new_n16802_;
  assign new_n17041_ = ~new_n16800_ & new_n17040_;
  assign new_n17042_ = ~new_n16804_ & ~new_n17041_;
  assign new_n17043_ = ~new_n17039_ & new_n17042_;
  assign new_n17044_ = ~new_n16804_ & ~new_n17043_;
  assign new_n17045_ = \b[19]  & ~new_n16793_;
  assign new_n17046_ = ~new_n16791_ & new_n17045_;
  assign new_n17047_ = ~new_n16795_ & ~new_n17046_;
  assign new_n17048_ = ~new_n17044_ & new_n17047_;
  assign new_n17049_ = ~new_n16795_ & ~new_n17048_;
  assign new_n17050_ = \b[20]  & ~new_n16784_;
  assign new_n17051_ = ~new_n16782_ & new_n17050_;
  assign new_n17052_ = ~new_n16786_ & ~new_n17051_;
  assign new_n17053_ = ~new_n17049_ & new_n17052_;
  assign new_n17054_ = ~new_n16786_ & ~new_n17053_;
  assign new_n17055_ = \b[21]  & ~new_n16775_;
  assign new_n17056_ = ~new_n16773_ & new_n17055_;
  assign new_n17057_ = ~new_n16777_ & ~new_n17056_;
  assign new_n17058_ = ~new_n17054_ & new_n17057_;
  assign new_n17059_ = ~new_n16777_ & ~new_n17058_;
  assign new_n17060_ = \b[22]  & ~new_n16766_;
  assign new_n17061_ = ~new_n16764_ & new_n17060_;
  assign new_n17062_ = ~new_n16768_ & ~new_n17061_;
  assign new_n17063_ = ~new_n17059_ & new_n17062_;
  assign new_n17064_ = ~new_n16768_ & ~new_n17063_;
  assign new_n17065_ = \b[23]  & ~new_n16757_;
  assign new_n17066_ = ~new_n16755_ & new_n17065_;
  assign new_n17067_ = ~new_n16759_ & ~new_n17066_;
  assign new_n17068_ = ~new_n17064_ & new_n17067_;
  assign new_n17069_ = ~new_n16759_ & ~new_n17068_;
  assign new_n17070_ = \b[24]  & ~new_n16748_;
  assign new_n17071_ = ~new_n16746_ & new_n17070_;
  assign new_n17072_ = ~new_n16750_ & ~new_n17071_;
  assign new_n17073_ = ~new_n17069_ & new_n17072_;
  assign new_n17074_ = ~new_n16750_ & ~new_n17073_;
  assign new_n17075_ = \b[25]  & ~new_n16739_;
  assign new_n17076_ = ~new_n16737_ & new_n17075_;
  assign new_n17077_ = ~new_n16741_ & ~new_n17076_;
  assign new_n17078_ = ~new_n17074_ & new_n17077_;
  assign new_n17079_ = ~new_n16741_ & ~new_n17078_;
  assign new_n17080_ = \b[26]  & ~new_n16730_;
  assign new_n17081_ = ~new_n16728_ & new_n17080_;
  assign new_n17082_ = ~new_n16732_ & ~new_n17081_;
  assign new_n17083_ = ~new_n17079_ & new_n17082_;
  assign new_n17084_ = ~new_n16732_ & ~new_n17083_;
  assign new_n17085_ = \b[27]  & ~new_n16721_;
  assign new_n17086_ = ~new_n16719_ & new_n17085_;
  assign new_n17087_ = ~new_n16723_ & ~new_n17086_;
  assign new_n17088_ = ~new_n17084_ & new_n17087_;
  assign new_n17089_ = ~new_n16723_ & ~new_n17088_;
  assign new_n17090_ = \b[28]  & ~new_n16712_;
  assign new_n17091_ = ~new_n16710_ & new_n17090_;
  assign new_n17092_ = ~new_n16714_ & ~new_n17091_;
  assign new_n17093_ = ~new_n17089_ & new_n17092_;
  assign new_n17094_ = ~new_n16714_ & ~new_n17093_;
  assign new_n17095_ = \b[29]  & ~new_n16703_;
  assign new_n17096_ = ~new_n16701_ & new_n17095_;
  assign new_n17097_ = ~new_n16705_ & ~new_n17096_;
  assign new_n17098_ = ~new_n17094_ & new_n17097_;
  assign new_n17099_ = ~new_n16705_ & ~new_n17098_;
  assign new_n17100_ = \b[30]  & ~new_n16694_;
  assign new_n17101_ = ~new_n16692_ & new_n17100_;
  assign new_n17102_ = ~new_n16696_ & ~new_n17101_;
  assign new_n17103_ = ~new_n17099_ & new_n17102_;
  assign new_n17104_ = ~new_n16696_ & ~new_n17103_;
  assign new_n17105_ = \b[31]  & ~new_n16685_;
  assign new_n17106_ = ~new_n16683_ & new_n17105_;
  assign new_n17107_ = ~new_n16687_ & ~new_n17106_;
  assign new_n17108_ = ~new_n17104_ & new_n17107_;
  assign new_n17109_ = ~new_n16687_ & ~new_n17108_;
  assign new_n17110_ = \b[32]  & ~new_n16676_;
  assign new_n17111_ = ~new_n16674_ & new_n17110_;
  assign new_n17112_ = ~new_n16678_ & ~new_n17111_;
  assign new_n17113_ = ~new_n17109_ & new_n17112_;
  assign new_n17114_ = ~new_n16678_ & ~new_n17113_;
  assign new_n17115_ = \b[33]  & ~new_n16667_;
  assign new_n17116_ = ~new_n16665_ & new_n17115_;
  assign new_n17117_ = ~new_n16669_ & ~new_n17116_;
  assign new_n17118_ = ~new_n17114_ & new_n17117_;
  assign new_n17119_ = ~new_n16669_ & ~new_n17118_;
  assign new_n17120_ = \b[34]  & ~new_n16658_;
  assign new_n17121_ = ~new_n16656_ & new_n17120_;
  assign new_n17122_ = ~new_n16660_ & ~new_n17121_;
  assign new_n17123_ = ~new_n17119_ & new_n17122_;
  assign new_n17124_ = ~new_n16660_ & ~new_n17123_;
  assign new_n17125_ = \b[35]  & ~new_n16649_;
  assign new_n17126_ = ~new_n16647_ & new_n17125_;
  assign new_n17127_ = ~new_n16651_ & ~new_n17126_;
  assign new_n17128_ = ~new_n17124_ & new_n17127_;
  assign new_n17129_ = ~new_n16651_ & ~new_n17128_;
  assign new_n17130_ = \b[36]  & ~new_n16640_;
  assign new_n17131_ = ~new_n16638_ & new_n17130_;
  assign new_n17132_ = ~new_n16642_ & ~new_n17131_;
  assign new_n17133_ = ~new_n17129_ & new_n17132_;
  assign new_n17134_ = ~new_n16642_ & ~new_n17133_;
  assign new_n17135_ = \b[37]  & ~new_n16631_;
  assign new_n17136_ = ~new_n16629_ & new_n17135_;
  assign new_n17137_ = ~new_n16633_ & ~new_n17136_;
  assign new_n17138_ = ~new_n17134_ & new_n17137_;
  assign new_n17139_ = ~new_n16633_ & ~new_n17138_;
  assign new_n17140_ = \b[38]  & ~new_n16622_;
  assign new_n17141_ = ~new_n16620_ & new_n17140_;
  assign new_n17142_ = ~new_n16624_ & ~new_n17141_;
  assign new_n17143_ = ~new_n17139_ & new_n17142_;
  assign new_n17144_ = ~new_n16624_ & ~new_n17143_;
  assign new_n17145_ = \b[39]  & ~new_n16613_;
  assign new_n17146_ = ~new_n16611_ & new_n17145_;
  assign new_n17147_ = ~new_n16615_ & ~new_n17146_;
  assign new_n17148_ = ~new_n17144_ & new_n17147_;
  assign new_n17149_ = ~new_n16615_ & ~new_n17148_;
  assign new_n17150_ = \b[40]  & ~new_n16604_;
  assign new_n17151_ = ~new_n16602_ & new_n17150_;
  assign new_n17152_ = ~new_n16606_ & ~new_n17151_;
  assign new_n17153_ = ~new_n17149_ & new_n17152_;
  assign new_n17154_ = ~new_n16606_ & ~new_n17153_;
  assign new_n17155_ = \b[41]  & ~new_n16595_;
  assign new_n17156_ = ~new_n16593_ & new_n17155_;
  assign new_n17157_ = ~new_n16597_ & ~new_n17156_;
  assign new_n17158_ = ~new_n17154_ & new_n17157_;
  assign new_n17159_ = ~new_n16597_ & ~new_n17158_;
  assign new_n17160_ = \b[42]  & ~new_n16586_;
  assign new_n17161_ = ~new_n16584_ & new_n17160_;
  assign new_n17162_ = ~new_n16588_ & ~new_n17161_;
  assign new_n17163_ = ~new_n17159_ & new_n17162_;
  assign new_n17164_ = ~new_n16588_ & ~new_n17163_;
  assign new_n17165_ = \b[43]  & ~new_n16577_;
  assign new_n17166_ = ~new_n16575_ & new_n17165_;
  assign new_n17167_ = ~new_n16579_ & ~new_n17166_;
  assign new_n17168_ = ~new_n17164_ & new_n17167_;
  assign new_n17169_ = ~new_n16579_ & ~new_n17168_;
  assign new_n17170_ = \b[44]  & ~new_n16568_;
  assign new_n17171_ = ~new_n16566_ & new_n17170_;
  assign new_n17172_ = ~new_n16570_ & ~new_n17171_;
  assign new_n17173_ = ~new_n17169_ & new_n17172_;
  assign new_n17174_ = ~new_n16570_ & ~new_n17173_;
  assign new_n17175_ = \b[45]  & ~new_n16559_;
  assign new_n17176_ = ~new_n16557_ & new_n17175_;
  assign new_n17177_ = ~new_n16561_ & ~new_n17176_;
  assign new_n17178_ = ~new_n17174_ & new_n17177_;
  assign new_n17179_ = ~new_n16561_ & ~new_n17178_;
  assign new_n17180_ = \b[46]  & ~new_n16550_;
  assign new_n17181_ = ~new_n16548_ & new_n17180_;
  assign new_n17182_ = ~new_n16552_ & ~new_n17181_;
  assign new_n17183_ = ~new_n17179_ & new_n17182_;
  assign new_n17184_ = ~new_n16552_ & ~new_n17183_;
  assign new_n17185_ = \b[47]  & ~new_n16530_;
  assign new_n17186_ = ~new_n16528_ & new_n17185_;
  assign new_n17187_ = ~new_n16543_ & ~new_n17186_;
  assign new_n17188_ = ~new_n17184_ & new_n17187_;
  assign new_n17189_ = ~new_n16543_ & ~new_n17188_;
  assign new_n17190_ = \b[48]  & ~new_n16540_;
  assign new_n17191_ = ~new_n16538_ & new_n17190_;
  assign new_n17192_ = ~new_n16542_ & ~new_n17191_;
  assign new_n17193_ = ~new_n17189_ & new_n17192_;
  assign new_n17194_ = ~new_n16542_ & ~new_n17193_;
  assign \quotient[15]  = new_n408_ & ~new_n17194_;
  assign new_n17196_ = ~new_n16531_ & ~\quotient[15] ;
  assign new_n17197_ = ~new_n16552_ & new_n17187_;
  assign new_n17198_ = ~new_n17183_ & new_n17197_;
  assign new_n17199_ = ~new_n17184_ & ~new_n17187_;
  assign new_n17200_ = ~new_n17198_ & ~new_n17199_;
  assign new_n17201_ = new_n408_ & ~new_n17200_;
  assign new_n17202_ = ~new_n17194_ & new_n17201_;
  assign new_n17203_ = ~new_n17196_ & ~new_n17202_;
  assign new_n17204_ = ~\b[48]  & ~new_n17203_;
  assign new_n17205_ = ~new_n16551_ & ~\quotient[15] ;
  assign new_n17206_ = ~new_n16561_ & new_n17182_;
  assign new_n17207_ = ~new_n17178_ & new_n17206_;
  assign new_n17208_ = ~new_n17179_ & ~new_n17182_;
  assign new_n17209_ = ~new_n17207_ & ~new_n17208_;
  assign new_n17210_ = new_n408_ & ~new_n17209_;
  assign new_n17211_ = ~new_n17194_ & new_n17210_;
  assign new_n17212_ = ~new_n17205_ & ~new_n17211_;
  assign new_n17213_ = ~\b[47]  & ~new_n17212_;
  assign new_n17214_ = ~new_n16560_ & ~\quotient[15] ;
  assign new_n17215_ = ~new_n16570_ & new_n17177_;
  assign new_n17216_ = ~new_n17173_ & new_n17215_;
  assign new_n17217_ = ~new_n17174_ & ~new_n17177_;
  assign new_n17218_ = ~new_n17216_ & ~new_n17217_;
  assign new_n17219_ = new_n408_ & ~new_n17218_;
  assign new_n17220_ = ~new_n17194_ & new_n17219_;
  assign new_n17221_ = ~new_n17214_ & ~new_n17220_;
  assign new_n17222_ = ~\b[46]  & ~new_n17221_;
  assign new_n17223_ = ~new_n16569_ & ~\quotient[15] ;
  assign new_n17224_ = ~new_n16579_ & new_n17172_;
  assign new_n17225_ = ~new_n17168_ & new_n17224_;
  assign new_n17226_ = ~new_n17169_ & ~new_n17172_;
  assign new_n17227_ = ~new_n17225_ & ~new_n17226_;
  assign new_n17228_ = new_n408_ & ~new_n17227_;
  assign new_n17229_ = ~new_n17194_ & new_n17228_;
  assign new_n17230_ = ~new_n17223_ & ~new_n17229_;
  assign new_n17231_ = ~\b[45]  & ~new_n17230_;
  assign new_n17232_ = ~new_n16578_ & ~\quotient[15] ;
  assign new_n17233_ = ~new_n16588_ & new_n17167_;
  assign new_n17234_ = ~new_n17163_ & new_n17233_;
  assign new_n17235_ = ~new_n17164_ & ~new_n17167_;
  assign new_n17236_ = ~new_n17234_ & ~new_n17235_;
  assign new_n17237_ = new_n408_ & ~new_n17236_;
  assign new_n17238_ = ~new_n17194_ & new_n17237_;
  assign new_n17239_ = ~new_n17232_ & ~new_n17238_;
  assign new_n17240_ = ~\b[44]  & ~new_n17239_;
  assign new_n17241_ = ~new_n16587_ & ~\quotient[15] ;
  assign new_n17242_ = ~new_n16597_ & new_n17162_;
  assign new_n17243_ = ~new_n17158_ & new_n17242_;
  assign new_n17244_ = ~new_n17159_ & ~new_n17162_;
  assign new_n17245_ = ~new_n17243_ & ~new_n17244_;
  assign new_n17246_ = new_n408_ & ~new_n17245_;
  assign new_n17247_ = ~new_n17194_ & new_n17246_;
  assign new_n17248_ = ~new_n17241_ & ~new_n17247_;
  assign new_n17249_ = ~\b[43]  & ~new_n17248_;
  assign new_n17250_ = ~new_n16596_ & ~\quotient[15] ;
  assign new_n17251_ = ~new_n16606_ & new_n17157_;
  assign new_n17252_ = ~new_n17153_ & new_n17251_;
  assign new_n17253_ = ~new_n17154_ & ~new_n17157_;
  assign new_n17254_ = ~new_n17252_ & ~new_n17253_;
  assign new_n17255_ = new_n408_ & ~new_n17254_;
  assign new_n17256_ = ~new_n17194_ & new_n17255_;
  assign new_n17257_ = ~new_n17250_ & ~new_n17256_;
  assign new_n17258_ = ~\b[42]  & ~new_n17257_;
  assign new_n17259_ = ~new_n16605_ & ~\quotient[15] ;
  assign new_n17260_ = ~new_n16615_ & new_n17152_;
  assign new_n17261_ = ~new_n17148_ & new_n17260_;
  assign new_n17262_ = ~new_n17149_ & ~new_n17152_;
  assign new_n17263_ = ~new_n17261_ & ~new_n17262_;
  assign new_n17264_ = new_n408_ & ~new_n17263_;
  assign new_n17265_ = ~new_n17194_ & new_n17264_;
  assign new_n17266_ = ~new_n17259_ & ~new_n17265_;
  assign new_n17267_ = ~\b[41]  & ~new_n17266_;
  assign new_n17268_ = ~new_n16614_ & ~\quotient[15] ;
  assign new_n17269_ = ~new_n16624_ & new_n17147_;
  assign new_n17270_ = ~new_n17143_ & new_n17269_;
  assign new_n17271_ = ~new_n17144_ & ~new_n17147_;
  assign new_n17272_ = ~new_n17270_ & ~new_n17271_;
  assign new_n17273_ = new_n408_ & ~new_n17272_;
  assign new_n17274_ = ~new_n17194_ & new_n17273_;
  assign new_n17275_ = ~new_n17268_ & ~new_n17274_;
  assign new_n17276_ = ~\b[40]  & ~new_n17275_;
  assign new_n17277_ = ~new_n16623_ & ~\quotient[15] ;
  assign new_n17278_ = ~new_n16633_ & new_n17142_;
  assign new_n17279_ = ~new_n17138_ & new_n17278_;
  assign new_n17280_ = ~new_n17139_ & ~new_n17142_;
  assign new_n17281_ = ~new_n17279_ & ~new_n17280_;
  assign new_n17282_ = new_n408_ & ~new_n17281_;
  assign new_n17283_ = ~new_n17194_ & new_n17282_;
  assign new_n17284_ = ~new_n17277_ & ~new_n17283_;
  assign new_n17285_ = ~\b[39]  & ~new_n17284_;
  assign new_n17286_ = ~new_n16632_ & ~\quotient[15] ;
  assign new_n17287_ = ~new_n16642_ & new_n17137_;
  assign new_n17288_ = ~new_n17133_ & new_n17287_;
  assign new_n17289_ = ~new_n17134_ & ~new_n17137_;
  assign new_n17290_ = ~new_n17288_ & ~new_n17289_;
  assign new_n17291_ = new_n408_ & ~new_n17290_;
  assign new_n17292_ = ~new_n17194_ & new_n17291_;
  assign new_n17293_ = ~new_n17286_ & ~new_n17292_;
  assign new_n17294_ = ~\b[38]  & ~new_n17293_;
  assign new_n17295_ = ~new_n16641_ & ~\quotient[15] ;
  assign new_n17296_ = ~new_n16651_ & new_n17132_;
  assign new_n17297_ = ~new_n17128_ & new_n17296_;
  assign new_n17298_ = ~new_n17129_ & ~new_n17132_;
  assign new_n17299_ = ~new_n17297_ & ~new_n17298_;
  assign new_n17300_ = new_n408_ & ~new_n17299_;
  assign new_n17301_ = ~new_n17194_ & new_n17300_;
  assign new_n17302_ = ~new_n17295_ & ~new_n17301_;
  assign new_n17303_ = ~\b[37]  & ~new_n17302_;
  assign new_n17304_ = ~new_n16650_ & ~\quotient[15] ;
  assign new_n17305_ = ~new_n16660_ & new_n17127_;
  assign new_n17306_ = ~new_n17123_ & new_n17305_;
  assign new_n17307_ = ~new_n17124_ & ~new_n17127_;
  assign new_n17308_ = ~new_n17306_ & ~new_n17307_;
  assign new_n17309_ = new_n408_ & ~new_n17308_;
  assign new_n17310_ = ~new_n17194_ & new_n17309_;
  assign new_n17311_ = ~new_n17304_ & ~new_n17310_;
  assign new_n17312_ = ~\b[36]  & ~new_n17311_;
  assign new_n17313_ = ~new_n16659_ & ~\quotient[15] ;
  assign new_n17314_ = ~new_n16669_ & new_n17122_;
  assign new_n17315_ = ~new_n17118_ & new_n17314_;
  assign new_n17316_ = ~new_n17119_ & ~new_n17122_;
  assign new_n17317_ = ~new_n17315_ & ~new_n17316_;
  assign new_n17318_ = new_n408_ & ~new_n17317_;
  assign new_n17319_ = ~new_n17194_ & new_n17318_;
  assign new_n17320_ = ~new_n17313_ & ~new_n17319_;
  assign new_n17321_ = ~\b[35]  & ~new_n17320_;
  assign new_n17322_ = ~new_n16668_ & ~\quotient[15] ;
  assign new_n17323_ = ~new_n16678_ & new_n17117_;
  assign new_n17324_ = ~new_n17113_ & new_n17323_;
  assign new_n17325_ = ~new_n17114_ & ~new_n17117_;
  assign new_n17326_ = ~new_n17324_ & ~new_n17325_;
  assign new_n17327_ = new_n408_ & ~new_n17326_;
  assign new_n17328_ = ~new_n17194_ & new_n17327_;
  assign new_n17329_ = ~new_n17322_ & ~new_n17328_;
  assign new_n17330_ = ~\b[34]  & ~new_n17329_;
  assign new_n17331_ = ~new_n16677_ & ~\quotient[15] ;
  assign new_n17332_ = ~new_n16687_ & new_n17112_;
  assign new_n17333_ = ~new_n17108_ & new_n17332_;
  assign new_n17334_ = ~new_n17109_ & ~new_n17112_;
  assign new_n17335_ = ~new_n17333_ & ~new_n17334_;
  assign new_n17336_ = new_n408_ & ~new_n17335_;
  assign new_n17337_ = ~new_n17194_ & new_n17336_;
  assign new_n17338_ = ~new_n17331_ & ~new_n17337_;
  assign new_n17339_ = ~\b[33]  & ~new_n17338_;
  assign new_n17340_ = ~new_n16686_ & ~\quotient[15] ;
  assign new_n17341_ = ~new_n16696_ & new_n17107_;
  assign new_n17342_ = ~new_n17103_ & new_n17341_;
  assign new_n17343_ = ~new_n17104_ & ~new_n17107_;
  assign new_n17344_ = ~new_n17342_ & ~new_n17343_;
  assign new_n17345_ = new_n408_ & ~new_n17344_;
  assign new_n17346_ = ~new_n17194_ & new_n17345_;
  assign new_n17347_ = ~new_n17340_ & ~new_n17346_;
  assign new_n17348_ = ~\b[32]  & ~new_n17347_;
  assign new_n17349_ = ~new_n16695_ & ~\quotient[15] ;
  assign new_n17350_ = ~new_n16705_ & new_n17102_;
  assign new_n17351_ = ~new_n17098_ & new_n17350_;
  assign new_n17352_ = ~new_n17099_ & ~new_n17102_;
  assign new_n17353_ = ~new_n17351_ & ~new_n17352_;
  assign new_n17354_ = new_n408_ & ~new_n17353_;
  assign new_n17355_ = ~new_n17194_ & new_n17354_;
  assign new_n17356_ = ~new_n17349_ & ~new_n17355_;
  assign new_n17357_ = ~\b[31]  & ~new_n17356_;
  assign new_n17358_ = ~new_n16704_ & ~\quotient[15] ;
  assign new_n17359_ = ~new_n16714_ & new_n17097_;
  assign new_n17360_ = ~new_n17093_ & new_n17359_;
  assign new_n17361_ = ~new_n17094_ & ~new_n17097_;
  assign new_n17362_ = ~new_n17360_ & ~new_n17361_;
  assign new_n17363_ = new_n408_ & ~new_n17362_;
  assign new_n17364_ = ~new_n17194_ & new_n17363_;
  assign new_n17365_ = ~new_n17358_ & ~new_n17364_;
  assign new_n17366_ = ~\b[30]  & ~new_n17365_;
  assign new_n17367_ = ~new_n16713_ & ~\quotient[15] ;
  assign new_n17368_ = ~new_n16723_ & new_n17092_;
  assign new_n17369_ = ~new_n17088_ & new_n17368_;
  assign new_n17370_ = ~new_n17089_ & ~new_n17092_;
  assign new_n17371_ = ~new_n17369_ & ~new_n17370_;
  assign new_n17372_ = new_n408_ & ~new_n17371_;
  assign new_n17373_ = ~new_n17194_ & new_n17372_;
  assign new_n17374_ = ~new_n17367_ & ~new_n17373_;
  assign new_n17375_ = ~\b[29]  & ~new_n17374_;
  assign new_n17376_ = ~new_n16722_ & ~\quotient[15] ;
  assign new_n17377_ = ~new_n16732_ & new_n17087_;
  assign new_n17378_ = ~new_n17083_ & new_n17377_;
  assign new_n17379_ = ~new_n17084_ & ~new_n17087_;
  assign new_n17380_ = ~new_n17378_ & ~new_n17379_;
  assign new_n17381_ = new_n408_ & ~new_n17380_;
  assign new_n17382_ = ~new_n17194_ & new_n17381_;
  assign new_n17383_ = ~new_n17376_ & ~new_n17382_;
  assign new_n17384_ = ~\b[28]  & ~new_n17383_;
  assign new_n17385_ = ~new_n16731_ & ~\quotient[15] ;
  assign new_n17386_ = ~new_n16741_ & new_n17082_;
  assign new_n17387_ = ~new_n17078_ & new_n17386_;
  assign new_n17388_ = ~new_n17079_ & ~new_n17082_;
  assign new_n17389_ = ~new_n17387_ & ~new_n17388_;
  assign new_n17390_ = new_n408_ & ~new_n17389_;
  assign new_n17391_ = ~new_n17194_ & new_n17390_;
  assign new_n17392_ = ~new_n17385_ & ~new_n17391_;
  assign new_n17393_ = ~\b[27]  & ~new_n17392_;
  assign new_n17394_ = ~new_n16740_ & ~\quotient[15] ;
  assign new_n17395_ = ~new_n16750_ & new_n17077_;
  assign new_n17396_ = ~new_n17073_ & new_n17395_;
  assign new_n17397_ = ~new_n17074_ & ~new_n17077_;
  assign new_n17398_ = ~new_n17396_ & ~new_n17397_;
  assign new_n17399_ = new_n408_ & ~new_n17398_;
  assign new_n17400_ = ~new_n17194_ & new_n17399_;
  assign new_n17401_ = ~new_n17394_ & ~new_n17400_;
  assign new_n17402_ = ~\b[26]  & ~new_n17401_;
  assign new_n17403_ = ~new_n16749_ & ~\quotient[15] ;
  assign new_n17404_ = ~new_n16759_ & new_n17072_;
  assign new_n17405_ = ~new_n17068_ & new_n17404_;
  assign new_n17406_ = ~new_n17069_ & ~new_n17072_;
  assign new_n17407_ = ~new_n17405_ & ~new_n17406_;
  assign new_n17408_ = new_n408_ & ~new_n17407_;
  assign new_n17409_ = ~new_n17194_ & new_n17408_;
  assign new_n17410_ = ~new_n17403_ & ~new_n17409_;
  assign new_n17411_ = ~\b[25]  & ~new_n17410_;
  assign new_n17412_ = ~new_n16758_ & ~\quotient[15] ;
  assign new_n17413_ = ~new_n16768_ & new_n17067_;
  assign new_n17414_ = ~new_n17063_ & new_n17413_;
  assign new_n17415_ = ~new_n17064_ & ~new_n17067_;
  assign new_n17416_ = ~new_n17414_ & ~new_n17415_;
  assign new_n17417_ = new_n408_ & ~new_n17416_;
  assign new_n17418_ = ~new_n17194_ & new_n17417_;
  assign new_n17419_ = ~new_n17412_ & ~new_n17418_;
  assign new_n17420_ = ~\b[24]  & ~new_n17419_;
  assign new_n17421_ = ~new_n16767_ & ~\quotient[15] ;
  assign new_n17422_ = ~new_n16777_ & new_n17062_;
  assign new_n17423_ = ~new_n17058_ & new_n17422_;
  assign new_n17424_ = ~new_n17059_ & ~new_n17062_;
  assign new_n17425_ = ~new_n17423_ & ~new_n17424_;
  assign new_n17426_ = new_n408_ & ~new_n17425_;
  assign new_n17427_ = ~new_n17194_ & new_n17426_;
  assign new_n17428_ = ~new_n17421_ & ~new_n17427_;
  assign new_n17429_ = ~\b[23]  & ~new_n17428_;
  assign new_n17430_ = ~new_n16776_ & ~\quotient[15] ;
  assign new_n17431_ = ~new_n16786_ & new_n17057_;
  assign new_n17432_ = ~new_n17053_ & new_n17431_;
  assign new_n17433_ = ~new_n17054_ & ~new_n17057_;
  assign new_n17434_ = ~new_n17432_ & ~new_n17433_;
  assign new_n17435_ = new_n408_ & ~new_n17434_;
  assign new_n17436_ = ~new_n17194_ & new_n17435_;
  assign new_n17437_ = ~new_n17430_ & ~new_n17436_;
  assign new_n17438_ = ~\b[22]  & ~new_n17437_;
  assign new_n17439_ = ~new_n16785_ & ~\quotient[15] ;
  assign new_n17440_ = ~new_n16795_ & new_n17052_;
  assign new_n17441_ = ~new_n17048_ & new_n17440_;
  assign new_n17442_ = ~new_n17049_ & ~new_n17052_;
  assign new_n17443_ = ~new_n17441_ & ~new_n17442_;
  assign new_n17444_ = new_n408_ & ~new_n17443_;
  assign new_n17445_ = ~new_n17194_ & new_n17444_;
  assign new_n17446_ = ~new_n17439_ & ~new_n17445_;
  assign new_n17447_ = ~\b[21]  & ~new_n17446_;
  assign new_n17448_ = ~new_n16794_ & ~\quotient[15] ;
  assign new_n17449_ = ~new_n16804_ & new_n17047_;
  assign new_n17450_ = ~new_n17043_ & new_n17449_;
  assign new_n17451_ = ~new_n17044_ & ~new_n17047_;
  assign new_n17452_ = ~new_n17450_ & ~new_n17451_;
  assign new_n17453_ = new_n408_ & ~new_n17452_;
  assign new_n17454_ = ~new_n17194_ & new_n17453_;
  assign new_n17455_ = ~new_n17448_ & ~new_n17454_;
  assign new_n17456_ = ~\b[20]  & ~new_n17455_;
  assign new_n17457_ = ~new_n16803_ & ~\quotient[15] ;
  assign new_n17458_ = ~new_n16813_ & new_n17042_;
  assign new_n17459_ = ~new_n17038_ & new_n17458_;
  assign new_n17460_ = ~new_n17039_ & ~new_n17042_;
  assign new_n17461_ = ~new_n17459_ & ~new_n17460_;
  assign new_n17462_ = new_n408_ & ~new_n17461_;
  assign new_n17463_ = ~new_n17194_ & new_n17462_;
  assign new_n17464_ = ~new_n17457_ & ~new_n17463_;
  assign new_n17465_ = ~\b[19]  & ~new_n17464_;
  assign new_n17466_ = ~new_n16812_ & ~\quotient[15] ;
  assign new_n17467_ = ~new_n16822_ & new_n17037_;
  assign new_n17468_ = ~new_n17033_ & new_n17467_;
  assign new_n17469_ = ~new_n17034_ & ~new_n17037_;
  assign new_n17470_ = ~new_n17468_ & ~new_n17469_;
  assign new_n17471_ = new_n408_ & ~new_n17470_;
  assign new_n17472_ = ~new_n17194_ & new_n17471_;
  assign new_n17473_ = ~new_n17466_ & ~new_n17472_;
  assign new_n17474_ = ~\b[18]  & ~new_n17473_;
  assign new_n17475_ = ~new_n16821_ & ~\quotient[15] ;
  assign new_n17476_ = ~new_n16831_ & new_n17032_;
  assign new_n17477_ = ~new_n17028_ & new_n17476_;
  assign new_n17478_ = ~new_n17029_ & ~new_n17032_;
  assign new_n17479_ = ~new_n17477_ & ~new_n17478_;
  assign new_n17480_ = new_n408_ & ~new_n17479_;
  assign new_n17481_ = ~new_n17194_ & new_n17480_;
  assign new_n17482_ = ~new_n17475_ & ~new_n17481_;
  assign new_n17483_ = ~\b[17]  & ~new_n17482_;
  assign new_n17484_ = ~new_n16830_ & ~\quotient[15] ;
  assign new_n17485_ = ~new_n16840_ & new_n17027_;
  assign new_n17486_ = ~new_n17023_ & new_n17485_;
  assign new_n17487_ = ~new_n17024_ & ~new_n17027_;
  assign new_n17488_ = ~new_n17486_ & ~new_n17487_;
  assign new_n17489_ = new_n408_ & ~new_n17488_;
  assign new_n17490_ = ~new_n17194_ & new_n17489_;
  assign new_n17491_ = ~new_n17484_ & ~new_n17490_;
  assign new_n17492_ = ~\b[16]  & ~new_n17491_;
  assign new_n17493_ = ~new_n16839_ & ~\quotient[15] ;
  assign new_n17494_ = ~new_n16849_ & new_n17022_;
  assign new_n17495_ = ~new_n17018_ & new_n17494_;
  assign new_n17496_ = ~new_n17019_ & ~new_n17022_;
  assign new_n17497_ = ~new_n17495_ & ~new_n17496_;
  assign new_n17498_ = new_n408_ & ~new_n17497_;
  assign new_n17499_ = ~new_n17194_ & new_n17498_;
  assign new_n17500_ = ~new_n17493_ & ~new_n17499_;
  assign new_n17501_ = ~\b[15]  & ~new_n17500_;
  assign new_n17502_ = ~new_n16848_ & ~\quotient[15] ;
  assign new_n17503_ = ~new_n16858_ & new_n17017_;
  assign new_n17504_ = ~new_n17013_ & new_n17503_;
  assign new_n17505_ = ~new_n17014_ & ~new_n17017_;
  assign new_n17506_ = ~new_n17504_ & ~new_n17505_;
  assign new_n17507_ = new_n408_ & ~new_n17506_;
  assign new_n17508_ = ~new_n17194_ & new_n17507_;
  assign new_n17509_ = ~new_n17502_ & ~new_n17508_;
  assign new_n17510_ = ~\b[14]  & ~new_n17509_;
  assign new_n17511_ = ~new_n16857_ & ~\quotient[15] ;
  assign new_n17512_ = ~new_n16867_ & new_n17012_;
  assign new_n17513_ = ~new_n17008_ & new_n17512_;
  assign new_n17514_ = ~new_n17009_ & ~new_n17012_;
  assign new_n17515_ = ~new_n17513_ & ~new_n17514_;
  assign new_n17516_ = new_n408_ & ~new_n17515_;
  assign new_n17517_ = ~new_n17194_ & new_n17516_;
  assign new_n17518_ = ~new_n17511_ & ~new_n17517_;
  assign new_n17519_ = ~\b[13]  & ~new_n17518_;
  assign new_n17520_ = ~new_n16866_ & ~\quotient[15] ;
  assign new_n17521_ = ~new_n16876_ & new_n17007_;
  assign new_n17522_ = ~new_n17003_ & new_n17521_;
  assign new_n17523_ = ~new_n17004_ & ~new_n17007_;
  assign new_n17524_ = ~new_n17522_ & ~new_n17523_;
  assign new_n17525_ = new_n408_ & ~new_n17524_;
  assign new_n17526_ = ~new_n17194_ & new_n17525_;
  assign new_n17527_ = ~new_n17520_ & ~new_n17526_;
  assign new_n17528_ = ~\b[12]  & ~new_n17527_;
  assign new_n17529_ = ~new_n16875_ & ~\quotient[15] ;
  assign new_n17530_ = ~new_n16885_ & new_n17002_;
  assign new_n17531_ = ~new_n16998_ & new_n17530_;
  assign new_n17532_ = ~new_n16999_ & ~new_n17002_;
  assign new_n17533_ = ~new_n17531_ & ~new_n17532_;
  assign new_n17534_ = new_n408_ & ~new_n17533_;
  assign new_n17535_ = ~new_n17194_ & new_n17534_;
  assign new_n17536_ = ~new_n17529_ & ~new_n17535_;
  assign new_n17537_ = ~\b[11]  & ~new_n17536_;
  assign new_n17538_ = ~new_n16884_ & ~\quotient[15] ;
  assign new_n17539_ = ~new_n16894_ & new_n16997_;
  assign new_n17540_ = ~new_n16993_ & new_n17539_;
  assign new_n17541_ = ~new_n16994_ & ~new_n16997_;
  assign new_n17542_ = ~new_n17540_ & ~new_n17541_;
  assign new_n17543_ = new_n408_ & ~new_n17542_;
  assign new_n17544_ = ~new_n17194_ & new_n17543_;
  assign new_n17545_ = ~new_n17538_ & ~new_n17544_;
  assign new_n17546_ = ~\b[10]  & ~new_n17545_;
  assign new_n17547_ = ~new_n16893_ & ~\quotient[15] ;
  assign new_n17548_ = ~new_n16903_ & new_n16992_;
  assign new_n17549_ = ~new_n16988_ & new_n17548_;
  assign new_n17550_ = ~new_n16989_ & ~new_n16992_;
  assign new_n17551_ = ~new_n17549_ & ~new_n17550_;
  assign new_n17552_ = new_n408_ & ~new_n17551_;
  assign new_n17553_ = ~new_n17194_ & new_n17552_;
  assign new_n17554_ = ~new_n17547_ & ~new_n17553_;
  assign new_n17555_ = ~\b[9]  & ~new_n17554_;
  assign new_n17556_ = ~new_n16902_ & ~\quotient[15] ;
  assign new_n17557_ = ~new_n16912_ & new_n16987_;
  assign new_n17558_ = ~new_n16983_ & new_n17557_;
  assign new_n17559_ = ~new_n16984_ & ~new_n16987_;
  assign new_n17560_ = ~new_n17558_ & ~new_n17559_;
  assign new_n17561_ = new_n408_ & ~new_n17560_;
  assign new_n17562_ = ~new_n17194_ & new_n17561_;
  assign new_n17563_ = ~new_n17556_ & ~new_n17562_;
  assign new_n17564_ = ~\b[8]  & ~new_n17563_;
  assign new_n17565_ = ~new_n16911_ & ~\quotient[15] ;
  assign new_n17566_ = ~new_n16921_ & new_n16982_;
  assign new_n17567_ = ~new_n16978_ & new_n17566_;
  assign new_n17568_ = ~new_n16979_ & ~new_n16982_;
  assign new_n17569_ = ~new_n17567_ & ~new_n17568_;
  assign new_n17570_ = new_n408_ & ~new_n17569_;
  assign new_n17571_ = ~new_n17194_ & new_n17570_;
  assign new_n17572_ = ~new_n17565_ & ~new_n17571_;
  assign new_n17573_ = ~\b[7]  & ~new_n17572_;
  assign new_n17574_ = ~new_n16920_ & ~\quotient[15] ;
  assign new_n17575_ = ~new_n16930_ & new_n16977_;
  assign new_n17576_ = ~new_n16973_ & new_n17575_;
  assign new_n17577_ = ~new_n16974_ & ~new_n16977_;
  assign new_n17578_ = ~new_n17576_ & ~new_n17577_;
  assign new_n17579_ = new_n408_ & ~new_n17578_;
  assign new_n17580_ = ~new_n17194_ & new_n17579_;
  assign new_n17581_ = ~new_n17574_ & ~new_n17580_;
  assign new_n17582_ = ~\b[6]  & ~new_n17581_;
  assign new_n17583_ = ~new_n16929_ & ~\quotient[15] ;
  assign new_n17584_ = ~new_n16939_ & new_n16972_;
  assign new_n17585_ = ~new_n16968_ & new_n17584_;
  assign new_n17586_ = ~new_n16969_ & ~new_n16972_;
  assign new_n17587_ = ~new_n17585_ & ~new_n17586_;
  assign new_n17588_ = new_n408_ & ~new_n17587_;
  assign new_n17589_ = ~new_n17194_ & new_n17588_;
  assign new_n17590_ = ~new_n17583_ & ~new_n17589_;
  assign new_n17591_ = ~\b[5]  & ~new_n17590_;
  assign new_n17592_ = ~new_n16938_ & ~\quotient[15] ;
  assign new_n17593_ = ~new_n16947_ & new_n16967_;
  assign new_n17594_ = ~new_n16963_ & new_n17593_;
  assign new_n17595_ = ~new_n16964_ & ~new_n16967_;
  assign new_n17596_ = ~new_n17594_ & ~new_n17595_;
  assign new_n17597_ = new_n408_ & ~new_n17596_;
  assign new_n17598_ = ~new_n17194_ & new_n17597_;
  assign new_n17599_ = ~new_n17592_ & ~new_n17598_;
  assign new_n17600_ = ~\b[4]  & ~new_n17599_;
  assign new_n17601_ = ~new_n16946_ & ~\quotient[15] ;
  assign new_n17602_ = ~new_n16958_ & new_n16962_;
  assign new_n17603_ = ~new_n16957_ & new_n17602_;
  assign new_n17604_ = ~new_n16959_ & ~new_n16962_;
  assign new_n17605_ = ~new_n17603_ & ~new_n17604_;
  assign new_n17606_ = new_n408_ & ~new_n17605_;
  assign new_n17607_ = ~new_n17194_ & new_n17606_;
  assign new_n17608_ = ~new_n17601_ & ~new_n17607_;
  assign new_n17609_ = ~\b[3]  & ~new_n17608_;
  assign new_n17610_ = ~new_n16951_ & ~\quotient[15] ;
  assign new_n17611_ = ~new_n16954_ & new_n16956_;
  assign new_n17612_ = ~new_n16952_ & new_n17611_;
  assign new_n17613_ = new_n408_ & ~new_n17612_;
  assign new_n17614_ = ~new_n16957_ & new_n17613_;
  assign new_n17615_ = ~new_n17194_ & new_n17614_;
  assign new_n17616_ = ~new_n17610_ & ~new_n17615_;
  assign new_n17617_ = ~\b[2]  & ~new_n17616_;
  assign new_n17618_ = \b[0]  & ~\b[49] ;
  assign new_n17619_ = new_n297_ & new_n17618_;
  assign new_n17620_ = new_n286_ & new_n17619_;
  assign new_n17621_ = new_n337_ & new_n17620_;
  assign new_n17622_ = ~new_n17194_ & new_n17621_;
  assign new_n17623_ = \a[15]  & ~new_n17622_;
  assign new_n17624_ = new_n400_ & new_n16956_;
  assign new_n17625_ = new_n595_ & new_n17624_;
  assign new_n17626_ = ~new_n17194_ & new_n17625_;
  assign new_n17627_ = ~new_n17623_ & ~new_n17626_;
  assign new_n17628_ = \b[1]  & ~new_n17627_;
  assign new_n17629_ = ~\b[1]  & ~new_n17626_;
  assign new_n17630_ = ~new_n17623_ & new_n17629_;
  assign new_n17631_ = ~new_n17628_ & ~new_n17630_;
  assign new_n17632_ = ~\a[14]  & \b[0] ;
  assign new_n17633_ = ~new_n17631_ & ~new_n17632_;
  assign new_n17634_ = ~\b[1]  & ~new_n17627_;
  assign new_n17635_ = ~new_n17633_ & ~new_n17634_;
  assign new_n17636_ = \b[2]  & ~new_n17615_;
  assign new_n17637_ = ~new_n17610_ & new_n17636_;
  assign new_n17638_ = ~new_n17617_ & ~new_n17637_;
  assign new_n17639_ = ~new_n17635_ & new_n17638_;
  assign new_n17640_ = ~new_n17617_ & ~new_n17639_;
  assign new_n17641_ = \b[3]  & ~new_n17607_;
  assign new_n17642_ = ~new_n17601_ & new_n17641_;
  assign new_n17643_ = ~new_n17609_ & ~new_n17642_;
  assign new_n17644_ = ~new_n17640_ & new_n17643_;
  assign new_n17645_ = ~new_n17609_ & ~new_n17644_;
  assign new_n17646_ = \b[4]  & ~new_n17598_;
  assign new_n17647_ = ~new_n17592_ & new_n17646_;
  assign new_n17648_ = ~new_n17600_ & ~new_n17647_;
  assign new_n17649_ = ~new_n17645_ & new_n17648_;
  assign new_n17650_ = ~new_n17600_ & ~new_n17649_;
  assign new_n17651_ = \b[5]  & ~new_n17589_;
  assign new_n17652_ = ~new_n17583_ & new_n17651_;
  assign new_n17653_ = ~new_n17591_ & ~new_n17652_;
  assign new_n17654_ = ~new_n17650_ & new_n17653_;
  assign new_n17655_ = ~new_n17591_ & ~new_n17654_;
  assign new_n17656_ = \b[6]  & ~new_n17580_;
  assign new_n17657_ = ~new_n17574_ & new_n17656_;
  assign new_n17658_ = ~new_n17582_ & ~new_n17657_;
  assign new_n17659_ = ~new_n17655_ & new_n17658_;
  assign new_n17660_ = ~new_n17582_ & ~new_n17659_;
  assign new_n17661_ = \b[7]  & ~new_n17571_;
  assign new_n17662_ = ~new_n17565_ & new_n17661_;
  assign new_n17663_ = ~new_n17573_ & ~new_n17662_;
  assign new_n17664_ = ~new_n17660_ & new_n17663_;
  assign new_n17665_ = ~new_n17573_ & ~new_n17664_;
  assign new_n17666_ = \b[8]  & ~new_n17562_;
  assign new_n17667_ = ~new_n17556_ & new_n17666_;
  assign new_n17668_ = ~new_n17564_ & ~new_n17667_;
  assign new_n17669_ = ~new_n17665_ & new_n17668_;
  assign new_n17670_ = ~new_n17564_ & ~new_n17669_;
  assign new_n17671_ = \b[9]  & ~new_n17553_;
  assign new_n17672_ = ~new_n17547_ & new_n17671_;
  assign new_n17673_ = ~new_n17555_ & ~new_n17672_;
  assign new_n17674_ = ~new_n17670_ & new_n17673_;
  assign new_n17675_ = ~new_n17555_ & ~new_n17674_;
  assign new_n17676_ = \b[10]  & ~new_n17544_;
  assign new_n17677_ = ~new_n17538_ & new_n17676_;
  assign new_n17678_ = ~new_n17546_ & ~new_n17677_;
  assign new_n17679_ = ~new_n17675_ & new_n17678_;
  assign new_n17680_ = ~new_n17546_ & ~new_n17679_;
  assign new_n17681_ = \b[11]  & ~new_n17535_;
  assign new_n17682_ = ~new_n17529_ & new_n17681_;
  assign new_n17683_ = ~new_n17537_ & ~new_n17682_;
  assign new_n17684_ = ~new_n17680_ & new_n17683_;
  assign new_n17685_ = ~new_n17537_ & ~new_n17684_;
  assign new_n17686_ = \b[12]  & ~new_n17526_;
  assign new_n17687_ = ~new_n17520_ & new_n17686_;
  assign new_n17688_ = ~new_n17528_ & ~new_n17687_;
  assign new_n17689_ = ~new_n17685_ & new_n17688_;
  assign new_n17690_ = ~new_n17528_ & ~new_n17689_;
  assign new_n17691_ = \b[13]  & ~new_n17517_;
  assign new_n17692_ = ~new_n17511_ & new_n17691_;
  assign new_n17693_ = ~new_n17519_ & ~new_n17692_;
  assign new_n17694_ = ~new_n17690_ & new_n17693_;
  assign new_n17695_ = ~new_n17519_ & ~new_n17694_;
  assign new_n17696_ = \b[14]  & ~new_n17508_;
  assign new_n17697_ = ~new_n17502_ & new_n17696_;
  assign new_n17698_ = ~new_n17510_ & ~new_n17697_;
  assign new_n17699_ = ~new_n17695_ & new_n17698_;
  assign new_n17700_ = ~new_n17510_ & ~new_n17699_;
  assign new_n17701_ = \b[15]  & ~new_n17499_;
  assign new_n17702_ = ~new_n17493_ & new_n17701_;
  assign new_n17703_ = ~new_n17501_ & ~new_n17702_;
  assign new_n17704_ = ~new_n17700_ & new_n17703_;
  assign new_n17705_ = ~new_n17501_ & ~new_n17704_;
  assign new_n17706_ = \b[16]  & ~new_n17490_;
  assign new_n17707_ = ~new_n17484_ & new_n17706_;
  assign new_n17708_ = ~new_n17492_ & ~new_n17707_;
  assign new_n17709_ = ~new_n17705_ & new_n17708_;
  assign new_n17710_ = ~new_n17492_ & ~new_n17709_;
  assign new_n17711_ = \b[17]  & ~new_n17481_;
  assign new_n17712_ = ~new_n17475_ & new_n17711_;
  assign new_n17713_ = ~new_n17483_ & ~new_n17712_;
  assign new_n17714_ = ~new_n17710_ & new_n17713_;
  assign new_n17715_ = ~new_n17483_ & ~new_n17714_;
  assign new_n17716_ = \b[18]  & ~new_n17472_;
  assign new_n17717_ = ~new_n17466_ & new_n17716_;
  assign new_n17718_ = ~new_n17474_ & ~new_n17717_;
  assign new_n17719_ = ~new_n17715_ & new_n17718_;
  assign new_n17720_ = ~new_n17474_ & ~new_n17719_;
  assign new_n17721_ = \b[19]  & ~new_n17463_;
  assign new_n17722_ = ~new_n17457_ & new_n17721_;
  assign new_n17723_ = ~new_n17465_ & ~new_n17722_;
  assign new_n17724_ = ~new_n17720_ & new_n17723_;
  assign new_n17725_ = ~new_n17465_ & ~new_n17724_;
  assign new_n17726_ = \b[20]  & ~new_n17454_;
  assign new_n17727_ = ~new_n17448_ & new_n17726_;
  assign new_n17728_ = ~new_n17456_ & ~new_n17727_;
  assign new_n17729_ = ~new_n17725_ & new_n17728_;
  assign new_n17730_ = ~new_n17456_ & ~new_n17729_;
  assign new_n17731_ = \b[21]  & ~new_n17445_;
  assign new_n17732_ = ~new_n17439_ & new_n17731_;
  assign new_n17733_ = ~new_n17447_ & ~new_n17732_;
  assign new_n17734_ = ~new_n17730_ & new_n17733_;
  assign new_n17735_ = ~new_n17447_ & ~new_n17734_;
  assign new_n17736_ = \b[22]  & ~new_n17436_;
  assign new_n17737_ = ~new_n17430_ & new_n17736_;
  assign new_n17738_ = ~new_n17438_ & ~new_n17737_;
  assign new_n17739_ = ~new_n17735_ & new_n17738_;
  assign new_n17740_ = ~new_n17438_ & ~new_n17739_;
  assign new_n17741_ = \b[23]  & ~new_n17427_;
  assign new_n17742_ = ~new_n17421_ & new_n17741_;
  assign new_n17743_ = ~new_n17429_ & ~new_n17742_;
  assign new_n17744_ = ~new_n17740_ & new_n17743_;
  assign new_n17745_ = ~new_n17429_ & ~new_n17744_;
  assign new_n17746_ = \b[24]  & ~new_n17418_;
  assign new_n17747_ = ~new_n17412_ & new_n17746_;
  assign new_n17748_ = ~new_n17420_ & ~new_n17747_;
  assign new_n17749_ = ~new_n17745_ & new_n17748_;
  assign new_n17750_ = ~new_n17420_ & ~new_n17749_;
  assign new_n17751_ = \b[25]  & ~new_n17409_;
  assign new_n17752_ = ~new_n17403_ & new_n17751_;
  assign new_n17753_ = ~new_n17411_ & ~new_n17752_;
  assign new_n17754_ = ~new_n17750_ & new_n17753_;
  assign new_n17755_ = ~new_n17411_ & ~new_n17754_;
  assign new_n17756_ = \b[26]  & ~new_n17400_;
  assign new_n17757_ = ~new_n17394_ & new_n17756_;
  assign new_n17758_ = ~new_n17402_ & ~new_n17757_;
  assign new_n17759_ = ~new_n17755_ & new_n17758_;
  assign new_n17760_ = ~new_n17402_ & ~new_n17759_;
  assign new_n17761_ = \b[27]  & ~new_n17391_;
  assign new_n17762_ = ~new_n17385_ & new_n17761_;
  assign new_n17763_ = ~new_n17393_ & ~new_n17762_;
  assign new_n17764_ = ~new_n17760_ & new_n17763_;
  assign new_n17765_ = ~new_n17393_ & ~new_n17764_;
  assign new_n17766_ = \b[28]  & ~new_n17382_;
  assign new_n17767_ = ~new_n17376_ & new_n17766_;
  assign new_n17768_ = ~new_n17384_ & ~new_n17767_;
  assign new_n17769_ = ~new_n17765_ & new_n17768_;
  assign new_n17770_ = ~new_n17384_ & ~new_n17769_;
  assign new_n17771_ = \b[29]  & ~new_n17373_;
  assign new_n17772_ = ~new_n17367_ & new_n17771_;
  assign new_n17773_ = ~new_n17375_ & ~new_n17772_;
  assign new_n17774_ = ~new_n17770_ & new_n17773_;
  assign new_n17775_ = ~new_n17375_ & ~new_n17774_;
  assign new_n17776_ = \b[30]  & ~new_n17364_;
  assign new_n17777_ = ~new_n17358_ & new_n17776_;
  assign new_n17778_ = ~new_n17366_ & ~new_n17777_;
  assign new_n17779_ = ~new_n17775_ & new_n17778_;
  assign new_n17780_ = ~new_n17366_ & ~new_n17779_;
  assign new_n17781_ = \b[31]  & ~new_n17355_;
  assign new_n17782_ = ~new_n17349_ & new_n17781_;
  assign new_n17783_ = ~new_n17357_ & ~new_n17782_;
  assign new_n17784_ = ~new_n17780_ & new_n17783_;
  assign new_n17785_ = ~new_n17357_ & ~new_n17784_;
  assign new_n17786_ = \b[32]  & ~new_n17346_;
  assign new_n17787_ = ~new_n17340_ & new_n17786_;
  assign new_n17788_ = ~new_n17348_ & ~new_n17787_;
  assign new_n17789_ = ~new_n17785_ & new_n17788_;
  assign new_n17790_ = ~new_n17348_ & ~new_n17789_;
  assign new_n17791_ = \b[33]  & ~new_n17337_;
  assign new_n17792_ = ~new_n17331_ & new_n17791_;
  assign new_n17793_ = ~new_n17339_ & ~new_n17792_;
  assign new_n17794_ = ~new_n17790_ & new_n17793_;
  assign new_n17795_ = ~new_n17339_ & ~new_n17794_;
  assign new_n17796_ = \b[34]  & ~new_n17328_;
  assign new_n17797_ = ~new_n17322_ & new_n17796_;
  assign new_n17798_ = ~new_n17330_ & ~new_n17797_;
  assign new_n17799_ = ~new_n17795_ & new_n17798_;
  assign new_n17800_ = ~new_n17330_ & ~new_n17799_;
  assign new_n17801_ = \b[35]  & ~new_n17319_;
  assign new_n17802_ = ~new_n17313_ & new_n17801_;
  assign new_n17803_ = ~new_n17321_ & ~new_n17802_;
  assign new_n17804_ = ~new_n17800_ & new_n17803_;
  assign new_n17805_ = ~new_n17321_ & ~new_n17804_;
  assign new_n17806_ = \b[36]  & ~new_n17310_;
  assign new_n17807_ = ~new_n17304_ & new_n17806_;
  assign new_n17808_ = ~new_n17312_ & ~new_n17807_;
  assign new_n17809_ = ~new_n17805_ & new_n17808_;
  assign new_n17810_ = ~new_n17312_ & ~new_n17809_;
  assign new_n17811_ = \b[37]  & ~new_n17301_;
  assign new_n17812_ = ~new_n17295_ & new_n17811_;
  assign new_n17813_ = ~new_n17303_ & ~new_n17812_;
  assign new_n17814_ = ~new_n17810_ & new_n17813_;
  assign new_n17815_ = ~new_n17303_ & ~new_n17814_;
  assign new_n17816_ = \b[38]  & ~new_n17292_;
  assign new_n17817_ = ~new_n17286_ & new_n17816_;
  assign new_n17818_ = ~new_n17294_ & ~new_n17817_;
  assign new_n17819_ = ~new_n17815_ & new_n17818_;
  assign new_n17820_ = ~new_n17294_ & ~new_n17819_;
  assign new_n17821_ = \b[39]  & ~new_n17283_;
  assign new_n17822_ = ~new_n17277_ & new_n17821_;
  assign new_n17823_ = ~new_n17285_ & ~new_n17822_;
  assign new_n17824_ = ~new_n17820_ & new_n17823_;
  assign new_n17825_ = ~new_n17285_ & ~new_n17824_;
  assign new_n17826_ = \b[40]  & ~new_n17274_;
  assign new_n17827_ = ~new_n17268_ & new_n17826_;
  assign new_n17828_ = ~new_n17276_ & ~new_n17827_;
  assign new_n17829_ = ~new_n17825_ & new_n17828_;
  assign new_n17830_ = ~new_n17276_ & ~new_n17829_;
  assign new_n17831_ = \b[41]  & ~new_n17265_;
  assign new_n17832_ = ~new_n17259_ & new_n17831_;
  assign new_n17833_ = ~new_n17267_ & ~new_n17832_;
  assign new_n17834_ = ~new_n17830_ & new_n17833_;
  assign new_n17835_ = ~new_n17267_ & ~new_n17834_;
  assign new_n17836_ = \b[42]  & ~new_n17256_;
  assign new_n17837_ = ~new_n17250_ & new_n17836_;
  assign new_n17838_ = ~new_n17258_ & ~new_n17837_;
  assign new_n17839_ = ~new_n17835_ & new_n17838_;
  assign new_n17840_ = ~new_n17258_ & ~new_n17839_;
  assign new_n17841_ = \b[43]  & ~new_n17247_;
  assign new_n17842_ = ~new_n17241_ & new_n17841_;
  assign new_n17843_ = ~new_n17249_ & ~new_n17842_;
  assign new_n17844_ = ~new_n17840_ & new_n17843_;
  assign new_n17845_ = ~new_n17249_ & ~new_n17844_;
  assign new_n17846_ = \b[44]  & ~new_n17238_;
  assign new_n17847_ = ~new_n17232_ & new_n17846_;
  assign new_n17848_ = ~new_n17240_ & ~new_n17847_;
  assign new_n17849_ = ~new_n17845_ & new_n17848_;
  assign new_n17850_ = ~new_n17240_ & ~new_n17849_;
  assign new_n17851_ = \b[45]  & ~new_n17229_;
  assign new_n17852_ = ~new_n17223_ & new_n17851_;
  assign new_n17853_ = ~new_n17231_ & ~new_n17852_;
  assign new_n17854_ = ~new_n17850_ & new_n17853_;
  assign new_n17855_ = ~new_n17231_ & ~new_n17854_;
  assign new_n17856_ = \b[46]  & ~new_n17220_;
  assign new_n17857_ = ~new_n17214_ & new_n17856_;
  assign new_n17858_ = ~new_n17222_ & ~new_n17857_;
  assign new_n17859_ = ~new_n17855_ & new_n17858_;
  assign new_n17860_ = ~new_n17222_ & ~new_n17859_;
  assign new_n17861_ = \b[47]  & ~new_n17211_;
  assign new_n17862_ = ~new_n17205_ & new_n17861_;
  assign new_n17863_ = ~new_n17213_ & ~new_n17862_;
  assign new_n17864_ = ~new_n17860_ & new_n17863_;
  assign new_n17865_ = ~new_n17213_ & ~new_n17864_;
  assign new_n17866_ = \b[48]  & ~new_n17202_;
  assign new_n17867_ = ~new_n17196_ & new_n17866_;
  assign new_n17868_ = ~new_n17204_ & ~new_n17867_;
  assign new_n17869_ = ~new_n17865_ & new_n17868_;
  assign new_n17870_ = ~new_n17204_ & ~new_n17869_;
  assign new_n17871_ = ~new_n16541_ & ~\quotient[15] ;
  assign new_n17872_ = ~new_n16543_ & new_n17192_;
  assign new_n17873_ = ~new_n17188_ & new_n17872_;
  assign new_n17874_ = ~new_n17189_ & ~new_n17192_;
  assign new_n17875_ = ~new_n17873_ & ~new_n17874_;
  assign new_n17876_ = \quotient[15]  & ~new_n17875_;
  assign new_n17877_ = ~new_n17871_ & ~new_n17876_;
  assign new_n17878_ = ~\b[49]  & ~new_n17877_;
  assign new_n17879_ = \b[49]  & ~new_n17871_;
  assign new_n17880_ = ~new_n17876_ & new_n17879_;
  assign new_n17881_ = new_n286_ & new_n297_;
  assign new_n17882_ = new_n337_ & new_n17881_;
  assign new_n17883_ = ~new_n17880_ & new_n17882_;
  assign new_n17884_ = ~new_n17878_ & new_n17883_;
  assign new_n17885_ = ~new_n17870_ & new_n17884_;
  assign new_n17886_ = new_n408_ & ~new_n17877_;
  assign \quotient[14]  = new_n17885_ | new_n17886_;
  assign new_n17888_ = ~new_n17213_ & new_n17868_;
  assign new_n17889_ = ~new_n17864_ & new_n17888_;
  assign new_n17890_ = ~new_n17865_ & ~new_n17868_;
  assign new_n17891_ = ~new_n17889_ & ~new_n17890_;
  assign new_n17892_ = \quotient[14]  & ~new_n17891_;
  assign new_n17893_ = ~new_n17203_ & ~new_n17886_;
  assign new_n17894_ = ~new_n17885_ & new_n17893_;
  assign new_n17895_ = ~new_n17892_ & ~new_n17894_;
  assign new_n17896_ = ~\b[49]  & ~new_n17895_;
  assign new_n17897_ = ~new_n17222_ & new_n17863_;
  assign new_n17898_ = ~new_n17859_ & new_n17897_;
  assign new_n17899_ = ~new_n17860_ & ~new_n17863_;
  assign new_n17900_ = ~new_n17898_ & ~new_n17899_;
  assign new_n17901_ = \quotient[14]  & ~new_n17900_;
  assign new_n17902_ = ~new_n17212_ & ~new_n17886_;
  assign new_n17903_ = ~new_n17885_ & new_n17902_;
  assign new_n17904_ = ~new_n17901_ & ~new_n17903_;
  assign new_n17905_ = ~\b[48]  & ~new_n17904_;
  assign new_n17906_ = ~new_n17231_ & new_n17858_;
  assign new_n17907_ = ~new_n17854_ & new_n17906_;
  assign new_n17908_ = ~new_n17855_ & ~new_n17858_;
  assign new_n17909_ = ~new_n17907_ & ~new_n17908_;
  assign new_n17910_ = \quotient[14]  & ~new_n17909_;
  assign new_n17911_ = ~new_n17221_ & ~new_n17886_;
  assign new_n17912_ = ~new_n17885_ & new_n17911_;
  assign new_n17913_ = ~new_n17910_ & ~new_n17912_;
  assign new_n17914_ = ~\b[47]  & ~new_n17913_;
  assign new_n17915_ = ~new_n17240_ & new_n17853_;
  assign new_n17916_ = ~new_n17849_ & new_n17915_;
  assign new_n17917_ = ~new_n17850_ & ~new_n17853_;
  assign new_n17918_ = ~new_n17916_ & ~new_n17917_;
  assign new_n17919_ = \quotient[14]  & ~new_n17918_;
  assign new_n17920_ = ~new_n17230_ & ~new_n17886_;
  assign new_n17921_ = ~new_n17885_ & new_n17920_;
  assign new_n17922_ = ~new_n17919_ & ~new_n17921_;
  assign new_n17923_ = ~\b[46]  & ~new_n17922_;
  assign new_n17924_ = ~new_n17249_ & new_n17848_;
  assign new_n17925_ = ~new_n17844_ & new_n17924_;
  assign new_n17926_ = ~new_n17845_ & ~new_n17848_;
  assign new_n17927_ = ~new_n17925_ & ~new_n17926_;
  assign new_n17928_ = \quotient[14]  & ~new_n17927_;
  assign new_n17929_ = ~new_n17239_ & ~new_n17886_;
  assign new_n17930_ = ~new_n17885_ & new_n17929_;
  assign new_n17931_ = ~new_n17928_ & ~new_n17930_;
  assign new_n17932_ = ~\b[45]  & ~new_n17931_;
  assign new_n17933_ = ~new_n17258_ & new_n17843_;
  assign new_n17934_ = ~new_n17839_ & new_n17933_;
  assign new_n17935_ = ~new_n17840_ & ~new_n17843_;
  assign new_n17936_ = ~new_n17934_ & ~new_n17935_;
  assign new_n17937_ = \quotient[14]  & ~new_n17936_;
  assign new_n17938_ = ~new_n17248_ & ~new_n17886_;
  assign new_n17939_ = ~new_n17885_ & new_n17938_;
  assign new_n17940_ = ~new_n17937_ & ~new_n17939_;
  assign new_n17941_ = ~\b[44]  & ~new_n17940_;
  assign new_n17942_ = ~new_n17267_ & new_n17838_;
  assign new_n17943_ = ~new_n17834_ & new_n17942_;
  assign new_n17944_ = ~new_n17835_ & ~new_n17838_;
  assign new_n17945_ = ~new_n17943_ & ~new_n17944_;
  assign new_n17946_ = \quotient[14]  & ~new_n17945_;
  assign new_n17947_ = ~new_n17257_ & ~new_n17886_;
  assign new_n17948_ = ~new_n17885_ & new_n17947_;
  assign new_n17949_ = ~new_n17946_ & ~new_n17948_;
  assign new_n17950_ = ~\b[43]  & ~new_n17949_;
  assign new_n17951_ = ~new_n17276_ & new_n17833_;
  assign new_n17952_ = ~new_n17829_ & new_n17951_;
  assign new_n17953_ = ~new_n17830_ & ~new_n17833_;
  assign new_n17954_ = ~new_n17952_ & ~new_n17953_;
  assign new_n17955_ = \quotient[14]  & ~new_n17954_;
  assign new_n17956_ = ~new_n17266_ & ~new_n17886_;
  assign new_n17957_ = ~new_n17885_ & new_n17956_;
  assign new_n17958_ = ~new_n17955_ & ~new_n17957_;
  assign new_n17959_ = ~\b[42]  & ~new_n17958_;
  assign new_n17960_ = ~new_n17285_ & new_n17828_;
  assign new_n17961_ = ~new_n17824_ & new_n17960_;
  assign new_n17962_ = ~new_n17825_ & ~new_n17828_;
  assign new_n17963_ = ~new_n17961_ & ~new_n17962_;
  assign new_n17964_ = \quotient[14]  & ~new_n17963_;
  assign new_n17965_ = ~new_n17275_ & ~new_n17886_;
  assign new_n17966_ = ~new_n17885_ & new_n17965_;
  assign new_n17967_ = ~new_n17964_ & ~new_n17966_;
  assign new_n17968_ = ~\b[41]  & ~new_n17967_;
  assign new_n17969_ = ~new_n17294_ & new_n17823_;
  assign new_n17970_ = ~new_n17819_ & new_n17969_;
  assign new_n17971_ = ~new_n17820_ & ~new_n17823_;
  assign new_n17972_ = ~new_n17970_ & ~new_n17971_;
  assign new_n17973_ = \quotient[14]  & ~new_n17972_;
  assign new_n17974_ = ~new_n17284_ & ~new_n17886_;
  assign new_n17975_ = ~new_n17885_ & new_n17974_;
  assign new_n17976_ = ~new_n17973_ & ~new_n17975_;
  assign new_n17977_ = ~\b[40]  & ~new_n17976_;
  assign new_n17978_ = ~new_n17303_ & new_n17818_;
  assign new_n17979_ = ~new_n17814_ & new_n17978_;
  assign new_n17980_ = ~new_n17815_ & ~new_n17818_;
  assign new_n17981_ = ~new_n17979_ & ~new_n17980_;
  assign new_n17982_ = \quotient[14]  & ~new_n17981_;
  assign new_n17983_ = ~new_n17293_ & ~new_n17886_;
  assign new_n17984_ = ~new_n17885_ & new_n17983_;
  assign new_n17985_ = ~new_n17982_ & ~new_n17984_;
  assign new_n17986_ = ~\b[39]  & ~new_n17985_;
  assign new_n17987_ = ~new_n17312_ & new_n17813_;
  assign new_n17988_ = ~new_n17809_ & new_n17987_;
  assign new_n17989_ = ~new_n17810_ & ~new_n17813_;
  assign new_n17990_ = ~new_n17988_ & ~new_n17989_;
  assign new_n17991_ = \quotient[14]  & ~new_n17990_;
  assign new_n17992_ = ~new_n17302_ & ~new_n17886_;
  assign new_n17993_ = ~new_n17885_ & new_n17992_;
  assign new_n17994_ = ~new_n17991_ & ~new_n17993_;
  assign new_n17995_ = ~\b[38]  & ~new_n17994_;
  assign new_n17996_ = ~new_n17321_ & new_n17808_;
  assign new_n17997_ = ~new_n17804_ & new_n17996_;
  assign new_n17998_ = ~new_n17805_ & ~new_n17808_;
  assign new_n17999_ = ~new_n17997_ & ~new_n17998_;
  assign new_n18000_ = \quotient[14]  & ~new_n17999_;
  assign new_n18001_ = ~new_n17311_ & ~new_n17886_;
  assign new_n18002_ = ~new_n17885_ & new_n18001_;
  assign new_n18003_ = ~new_n18000_ & ~new_n18002_;
  assign new_n18004_ = ~\b[37]  & ~new_n18003_;
  assign new_n18005_ = ~new_n17330_ & new_n17803_;
  assign new_n18006_ = ~new_n17799_ & new_n18005_;
  assign new_n18007_ = ~new_n17800_ & ~new_n17803_;
  assign new_n18008_ = ~new_n18006_ & ~new_n18007_;
  assign new_n18009_ = \quotient[14]  & ~new_n18008_;
  assign new_n18010_ = ~new_n17320_ & ~new_n17886_;
  assign new_n18011_ = ~new_n17885_ & new_n18010_;
  assign new_n18012_ = ~new_n18009_ & ~new_n18011_;
  assign new_n18013_ = ~\b[36]  & ~new_n18012_;
  assign new_n18014_ = ~new_n17339_ & new_n17798_;
  assign new_n18015_ = ~new_n17794_ & new_n18014_;
  assign new_n18016_ = ~new_n17795_ & ~new_n17798_;
  assign new_n18017_ = ~new_n18015_ & ~new_n18016_;
  assign new_n18018_ = \quotient[14]  & ~new_n18017_;
  assign new_n18019_ = ~new_n17329_ & ~new_n17886_;
  assign new_n18020_ = ~new_n17885_ & new_n18019_;
  assign new_n18021_ = ~new_n18018_ & ~new_n18020_;
  assign new_n18022_ = ~\b[35]  & ~new_n18021_;
  assign new_n18023_ = ~new_n17348_ & new_n17793_;
  assign new_n18024_ = ~new_n17789_ & new_n18023_;
  assign new_n18025_ = ~new_n17790_ & ~new_n17793_;
  assign new_n18026_ = ~new_n18024_ & ~new_n18025_;
  assign new_n18027_ = \quotient[14]  & ~new_n18026_;
  assign new_n18028_ = ~new_n17338_ & ~new_n17886_;
  assign new_n18029_ = ~new_n17885_ & new_n18028_;
  assign new_n18030_ = ~new_n18027_ & ~new_n18029_;
  assign new_n18031_ = ~\b[34]  & ~new_n18030_;
  assign new_n18032_ = ~new_n17357_ & new_n17788_;
  assign new_n18033_ = ~new_n17784_ & new_n18032_;
  assign new_n18034_ = ~new_n17785_ & ~new_n17788_;
  assign new_n18035_ = ~new_n18033_ & ~new_n18034_;
  assign new_n18036_ = \quotient[14]  & ~new_n18035_;
  assign new_n18037_ = ~new_n17347_ & ~new_n17886_;
  assign new_n18038_ = ~new_n17885_ & new_n18037_;
  assign new_n18039_ = ~new_n18036_ & ~new_n18038_;
  assign new_n18040_ = ~\b[33]  & ~new_n18039_;
  assign new_n18041_ = ~new_n17366_ & new_n17783_;
  assign new_n18042_ = ~new_n17779_ & new_n18041_;
  assign new_n18043_ = ~new_n17780_ & ~new_n17783_;
  assign new_n18044_ = ~new_n18042_ & ~new_n18043_;
  assign new_n18045_ = \quotient[14]  & ~new_n18044_;
  assign new_n18046_ = ~new_n17356_ & ~new_n17886_;
  assign new_n18047_ = ~new_n17885_ & new_n18046_;
  assign new_n18048_ = ~new_n18045_ & ~new_n18047_;
  assign new_n18049_ = ~\b[32]  & ~new_n18048_;
  assign new_n18050_ = ~new_n17375_ & new_n17778_;
  assign new_n18051_ = ~new_n17774_ & new_n18050_;
  assign new_n18052_ = ~new_n17775_ & ~new_n17778_;
  assign new_n18053_ = ~new_n18051_ & ~new_n18052_;
  assign new_n18054_ = \quotient[14]  & ~new_n18053_;
  assign new_n18055_ = ~new_n17365_ & ~new_n17886_;
  assign new_n18056_ = ~new_n17885_ & new_n18055_;
  assign new_n18057_ = ~new_n18054_ & ~new_n18056_;
  assign new_n18058_ = ~\b[31]  & ~new_n18057_;
  assign new_n18059_ = ~new_n17384_ & new_n17773_;
  assign new_n18060_ = ~new_n17769_ & new_n18059_;
  assign new_n18061_ = ~new_n17770_ & ~new_n17773_;
  assign new_n18062_ = ~new_n18060_ & ~new_n18061_;
  assign new_n18063_ = \quotient[14]  & ~new_n18062_;
  assign new_n18064_ = ~new_n17374_ & ~new_n17886_;
  assign new_n18065_ = ~new_n17885_ & new_n18064_;
  assign new_n18066_ = ~new_n18063_ & ~new_n18065_;
  assign new_n18067_ = ~\b[30]  & ~new_n18066_;
  assign new_n18068_ = ~new_n17393_ & new_n17768_;
  assign new_n18069_ = ~new_n17764_ & new_n18068_;
  assign new_n18070_ = ~new_n17765_ & ~new_n17768_;
  assign new_n18071_ = ~new_n18069_ & ~new_n18070_;
  assign new_n18072_ = \quotient[14]  & ~new_n18071_;
  assign new_n18073_ = ~new_n17383_ & ~new_n17886_;
  assign new_n18074_ = ~new_n17885_ & new_n18073_;
  assign new_n18075_ = ~new_n18072_ & ~new_n18074_;
  assign new_n18076_ = ~\b[29]  & ~new_n18075_;
  assign new_n18077_ = ~new_n17402_ & new_n17763_;
  assign new_n18078_ = ~new_n17759_ & new_n18077_;
  assign new_n18079_ = ~new_n17760_ & ~new_n17763_;
  assign new_n18080_ = ~new_n18078_ & ~new_n18079_;
  assign new_n18081_ = \quotient[14]  & ~new_n18080_;
  assign new_n18082_ = ~new_n17392_ & ~new_n17886_;
  assign new_n18083_ = ~new_n17885_ & new_n18082_;
  assign new_n18084_ = ~new_n18081_ & ~new_n18083_;
  assign new_n18085_ = ~\b[28]  & ~new_n18084_;
  assign new_n18086_ = ~new_n17411_ & new_n17758_;
  assign new_n18087_ = ~new_n17754_ & new_n18086_;
  assign new_n18088_ = ~new_n17755_ & ~new_n17758_;
  assign new_n18089_ = ~new_n18087_ & ~new_n18088_;
  assign new_n18090_ = \quotient[14]  & ~new_n18089_;
  assign new_n18091_ = ~new_n17401_ & ~new_n17886_;
  assign new_n18092_ = ~new_n17885_ & new_n18091_;
  assign new_n18093_ = ~new_n18090_ & ~new_n18092_;
  assign new_n18094_ = ~\b[27]  & ~new_n18093_;
  assign new_n18095_ = ~new_n17420_ & new_n17753_;
  assign new_n18096_ = ~new_n17749_ & new_n18095_;
  assign new_n18097_ = ~new_n17750_ & ~new_n17753_;
  assign new_n18098_ = ~new_n18096_ & ~new_n18097_;
  assign new_n18099_ = \quotient[14]  & ~new_n18098_;
  assign new_n18100_ = ~new_n17410_ & ~new_n17886_;
  assign new_n18101_ = ~new_n17885_ & new_n18100_;
  assign new_n18102_ = ~new_n18099_ & ~new_n18101_;
  assign new_n18103_ = ~\b[26]  & ~new_n18102_;
  assign new_n18104_ = ~new_n17429_ & new_n17748_;
  assign new_n18105_ = ~new_n17744_ & new_n18104_;
  assign new_n18106_ = ~new_n17745_ & ~new_n17748_;
  assign new_n18107_ = ~new_n18105_ & ~new_n18106_;
  assign new_n18108_ = \quotient[14]  & ~new_n18107_;
  assign new_n18109_ = ~new_n17419_ & ~new_n17886_;
  assign new_n18110_ = ~new_n17885_ & new_n18109_;
  assign new_n18111_ = ~new_n18108_ & ~new_n18110_;
  assign new_n18112_ = ~\b[25]  & ~new_n18111_;
  assign new_n18113_ = ~new_n17438_ & new_n17743_;
  assign new_n18114_ = ~new_n17739_ & new_n18113_;
  assign new_n18115_ = ~new_n17740_ & ~new_n17743_;
  assign new_n18116_ = ~new_n18114_ & ~new_n18115_;
  assign new_n18117_ = \quotient[14]  & ~new_n18116_;
  assign new_n18118_ = ~new_n17428_ & ~new_n17886_;
  assign new_n18119_ = ~new_n17885_ & new_n18118_;
  assign new_n18120_ = ~new_n18117_ & ~new_n18119_;
  assign new_n18121_ = ~\b[24]  & ~new_n18120_;
  assign new_n18122_ = ~new_n17447_ & new_n17738_;
  assign new_n18123_ = ~new_n17734_ & new_n18122_;
  assign new_n18124_ = ~new_n17735_ & ~new_n17738_;
  assign new_n18125_ = ~new_n18123_ & ~new_n18124_;
  assign new_n18126_ = \quotient[14]  & ~new_n18125_;
  assign new_n18127_ = ~new_n17437_ & ~new_n17886_;
  assign new_n18128_ = ~new_n17885_ & new_n18127_;
  assign new_n18129_ = ~new_n18126_ & ~new_n18128_;
  assign new_n18130_ = ~\b[23]  & ~new_n18129_;
  assign new_n18131_ = ~new_n17456_ & new_n17733_;
  assign new_n18132_ = ~new_n17729_ & new_n18131_;
  assign new_n18133_ = ~new_n17730_ & ~new_n17733_;
  assign new_n18134_ = ~new_n18132_ & ~new_n18133_;
  assign new_n18135_ = \quotient[14]  & ~new_n18134_;
  assign new_n18136_ = ~new_n17446_ & ~new_n17886_;
  assign new_n18137_ = ~new_n17885_ & new_n18136_;
  assign new_n18138_ = ~new_n18135_ & ~new_n18137_;
  assign new_n18139_ = ~\b[22]  & ~new_n18138_;
  assign new_n18140_ = ~new_n17465_ & new_n17728_;
  assign new_n18141_ = ~new_n17724_ & new_n18140_;
  assign new_n18142_ = ~new_n17725_ & ~new_n17728_;
  assign new_n18143_ = ~new_n18141_ & ~new_n18142_;
  assign new_n18144_ = \quotient[14]  & ~new_n18143_;
  assign new_n18145_ = ~new_n17455_ & ~new_n17886_;
  assign new_n18146_ = ~new_n17885_ & new_n18145_;
  assign new_n18147_ = ~new_n18144_ & ~new_n18146_;
  assign new_n18148_ = ~\b[21]  & ~new_n18147_;
  assign new_n18149_ = ~new_n17474_ & new_n17723_;
  assign new_n18150_ = ~new_n17719_ & new_n18149_;
  assign new_n18151_ = ~new_n17720_ & ~new_n17723_;
  assign new_n18152_ = ~new_n18150_ & ~new_n18151_;
  assign new_n18153_ = \quotient[14]  & ~new_n18152_;
  assign new_n18154_ = ~new_n17464_ & ~new_n17886_;
  assign new_n18155_ = ~new_n17885_ & new_n18154_;
  assign new_n18156_ = ~new_n18153_ & ~new_n18155_;
  assign new_n18157_ = ~\b[20]  & ~new_n18156_;
  assign new_n18158_ = ~new_n17483_ & new_n17718_;
  assign new_n18159_ = ~new_n17714_ & new_n18158_;
  assign new_n18160_ = ~new_n17715_ & ~new_n17718_;
  assign new_n18161_ = ~new_n18159_ & ~new_n18160_;
  assign new_n18162_ = \quotient[14]  & ~new_n18161_;
  assign new_n18163_ = ~new_n17473_ & ~new_n17886_;
  assign new_n18164_ = ~new_n17885_ & new_n18163_;
  assign new_n18165_ = ~new_n18162_ & ~new_n18164_;
  assign new_n18166_ = ~\b[19]  & ~new_n18165_;
  assign new_n18167_ = ~new_n17492_ & new_n17713_;
  assign new_n18168_ = ~new_n17709_ & new_n18167_;
  assign new_n18169_ = ~new_n17710_ & ~new_n17713_;
  assign new_n18170_ = ~new_n18168_ & ~new_n18169_;
  assign new_n18171_ = \quotient[14]  & ~new_n18170_;
  assign new_n18172_ = ~new_n17482_ & ~new_n17886_;
  assign new_n18173_ = ~new_n17885_ & new_n18172_;
  assign new_n18174_ = ~new_n18171_ & ~new_n18173_;
  assign new_n18175_ = ~\b[18]  & ~new_n18174_;
  assign new_n18176_ = ~new_n17501_ & new_n17708_;
  assign new_n18177_ = ~new_n17704_ & new_n18176_;
  assign new_n18178_ = ~new_n17705_ & ~new_n17708_;
  assign new_n18179_ = ~new_n18177_ & ~new_n18178_;
  assign new_n18180_ = \quotient[14]  & ~new_n18179_;
  assign new_n18181_ = ~new_n17491_ & ~new_n17886_;
  assign new_n18182_ = ~new_n17885_ & new_n18181_;
  assign new_n18183_ = ~new_n18180_ & ~new_n18182_;
  assign new_n18184_ = ~\b[17]  & ~new_n18183_;
  assign new_n18185_ = ~new_n17510_ & new_n17703_;
  assign new_n18186_ = ~new_n17699_ & new_n18185_;
  assign new_n18187_ = ~new_n17700_ & ~new_n17703_;
  assign new_n18188_ = ~new_n18186_ & ~new_n18187_;
  assign new_n18189_ = \quotient[14]  & ~new_n18188_;
  assign new_n18190_ = ~new_n17500_ & ~new_n17886_;
  assign new_n18191_ = ~new_n17885_ & new_n18190_;
  assign new_n18192_ = ~new_n18189_ & ~new_n18191_;
  assign new_n18193_ = ~\b[16]  & ~new_n18192_;
  assign new_n18194_ = ~new_n17519_ & new_n17698_;
  assign new_n18195_ = ~new_n17694_ & new_n18194_;
  assign new_n18196_ = ~new_n17695_ & ~new_n17698_;
  assign new_n18197_ = ~new_n18195_ & ~new_n18196_;
  assign new_n18198_ = \quotient[14]  & ~new_n18197_;
  assign new_n18199_ = ~new_n17509_ & ~new_n17886_;
  assign new_n18200_ = ~new_n17885_ & new_n18199_;
  assign new_n18201_ = ~new_n18198_ & ~new_n18200_;
  assign new_n18202_ = ~\b[15]  & ~new_n18201_;
  assign new_n18203_ = ~new_n17528_ & new_n17693_;
  assign new_n18204_ = ~new_n17689_ & new_n18203_;
  assign new_n18205_ = ~new_n17690_ & ~new_n17693_;
  assign new_n18206_ = ~new_n18204_ & ~new_n18205_;
  assign new_n18207_ = \quotient[14]  & ~new_n18206_;
  assign new_n18208_ = ~new_n17518_ & ~new_n17886_;
  assign new_n18209_ = ~new_n17885_ & new_n18208_;
  assign new_n18210_ = ~new_n18207_ & ~new_n18209_;
  assign new_n18211_ = ~\b[14]  & ~new_n18210_;
  assign new_n18212_ = ~new_n17537_ & new_n17688_;
  assign new_n18213_ = ~new_n17684_ & new_n18212_;
  assign new_n18214_ = ~new_n17685_ & ~new_n17688_;
  assign new_n18215_ = ~new_n18213_ & ~new_n18214_;
  assign new_n18216_ = \quotient[14]  & ~new_n18215_;
  assign new_n18217_ = ~new_n17527_ & ~new_n17886_;
  assign new_n18218_ = ~new_n17885_ & new_n18217_;
  assign new_n18219_ = ~new_n18216_ & ~new_n18218_;
  assign new_n18220_ = ~\b[13]  & ~new_n18219_;
  assign new_n18221_ = ~new_n17546_ & new_n17683_;
  assign new_n18222_ = ~new_n17679_ & new_n18221_;
  assign new_n18223_ = ~new_n17680_ & ~new_n17683_;
  assign new_n18224_ = ~new_n18222_ & ~new_n18223_;
  assign new_n18225_ = \quotient[14]  & ~new_n18224_;
  assign new_n18226_ = ~new_n17536_ & ~new_n17886_;
  assign new_n18227_ = ~new_n17885_ & new_n18226_;
  assign new_n18228_ = ~new_n18225_ & ~new_n18227_;
  assign new_n18229_ = ~\b[12]  & ~new_n18228_;
  assign new_n18230_ = ~new_n17555_ & new_n17678_;
  assign new_n18231_ = ~new_n17674_ & new_n18230_;
  assign new_n18232_ = ~new_n17675_ & ~new_n17678_;
  assign new_n18233_ = ~new_n18231_ & ~new_n18232_;
  assign new_n18234_ = \quotient[14]  & ~new_n18233_;
  assign new_n18235_ = ~new_n17545_ & ~new_n17886_;
  assign new_n18236_ = ~new_n17885_ & new_n18235_;
  assign new_n18237_ = ~new_n18234_ & ~new_n18236_;
  assign new_n18238_ = ~\b[11]  & ~new_n18237_;
  assign new_n18239_ = ~new_n17564_ & new_n17673_;
  assign new_n18240_ = ~new_n17669_ & new_n18239_;
  assign new_n18241_ = ~new_n17670_ & ~new_n17673_;
  assign new_n18242_ = ~new_n18240_ & ~new_n18241_;
  assign new_n18243_ = \quotient[14]  & ~new_n18242_;
  assign new_n18244_ = ~new_n17554_ & ~new_n17886_;
  assign new_n18245_ = ~new_n17885_ & new_n18244_;
  assign new_n18246_ = ~new_n18243_ & ~new_n18245_;
  assign new_n18247_ = ~\b[10]  & ~new_n18246_;
  assign new_n18248_ = ~new_n17573_ & new_n17668_;
  assign new_n18249_ = ~new_n17664_ & new_n18248_;
  assign new_n18250_ = ~new_n17665_ & ~new_n17668_;
  assign new_n18251_ = ~new_n18249_ & ~new_n18250_;
  assign new_n18252_ = \quotient[14]  & ~new_n18251_;
  assign new_n18253_ = ~new_n17563_ & ~new_n17886_;
  assign new_n18254_ = ~new_n17885_ & new_n18253_;
  assign new_n18255_ = ~new_n18252_ & ~new_n18254_;
  assign new_n18256_ = ~\b[9]  & ~new_n18255_;
  assign new_n18257_ = ~new_n17582_ & new_n17663_;
  assign new_n18258_ = ~new_n17659_ & new_n18257_;
  assign new_n18259_ = ~new_n17660_ & ~new_n17663_;
  assign new_n18260_ = ~new_n18258_ & ~new_n18259_;
  assign new_n18261_ = \quotient[14]  & ~new_n18260_;
  assign new_n18262_ = ~new_n17572_ & ~new_n17886_;
  assign new_n18263_ = ~new_n17885_ & new_n18262_;
  assign new_n18264_ = ~new_n18261_ & ~new_n18263_;
  assign new_n18265_ = ~\b[8]  & ~new_n18264_;
  assign new_n18266_ = ~new_n17591_ & new_n17658_;
  assign new_n18267_ = ~new_n17654_ & new_n18266_;
  assign new_n18268_ = ~new_n17655_ & ~new_n17658_;
  assign new_n18269_ = ~new_n18267_ & ~new_n18268_;
  assign new_n18270_ = \quotient[14]  & ~new_n18269_;
  assign new_n18271_ = ~new_n17581_ & ~new_n17886_;
  assign new_n18272_ = ~new_n17885_ & new_n18271_;
  assign new_n18273_ = ~new_n18270_ & ~new_n18272_;
  assign new_n18274_ = ~\b[7]  & ~new_n18273_;
  assign new_n18275_ = ~new_n17600_ & new_n17653_;
  assign new_n18276_ = ~new_n17649_ & new_n18275_;
  assign new_n18277_ = ~new_n17650_ & ~new_n17653_;
  assign new_n18278_ = ~new_n18276_ & ~new_n18277_;
  assign new_n18279_ = \quotient[14]  & ~new_n18278_;
  assign new_n18280_ = ~new_n17590_ & ~new_n17886_;
  assign new_n18281_ = ~new_n17885_ & new_n18280_;
  assign new_n18282_ = ~new_n18279_ & ~new_n18281_;
  assign new_n18283_ = ~\b[6]  & ~new_n18282_;
  assign new_n18284_ = ~new_n17609_ & new_n17648_;
  assign new_n18285_ = ~new_n17644_ & new_n18284_;
  assign new_n18286_ = ~new_n17645_ & ~new_n17648_;
  assign new_n18287_ = ~new_n18285_ & ~new_n18286_;
  assign new_n18288_ = \quotient[14]  & ~new_n18287_;
  assign new_n18289_ = ~new_n17599_ & ~new_n17886_;
  assign new_n18290_ = ~new_n17885_ & new_n18289_;
  assign new_n18291_ = ~new_n18288_ & ~new_n18290_;
  assign new_n18292_ = ~\b[5]  & ~new_n18291_;
  assign new_n18293_ = ~new_n17617_ & new_n17643_;
  assign new_n18294_ = ~new_n17639_ & new_n18293_;
  assign new_n18295_ = ~new_n17640_ & ~new_n17643_;
  assign new_n18296_ = ~new_n18294_ & ~new_n18295_;
  assign new_n18297_ = \quotient[14]  & ~new_n18296_;
  assign new_n18298_ = ~new_n17608_ & ~new_n17886_;
  assign new_n18299_ = ~new_n17885_ & new_n18298_;
  assign new_n18300_ = ~new_n18297_ & ~new_n18299_;
  assign new_n18301_ = ~\b[4]  & ~new_n18300_;
  assign new_n18302_ = ~new_n17634_ & new_n17638_;
  assign new_n18303_ = ~new_n17633_ & new_n18302_;
  assign new_n18304_ = ~new_n17635_ & ~new_n17638_;
  assign new_n18305_ = ~new_n18303_ & ~new_n18304_;
  assign new_n18306_ = \quotient[14]  & ~new_n18305_;
  assign new_n18307_ = ~new_n17616_ & ~new_n17886_;
  assign new_n18308_ = ~new_n17885_ & new_n18307_;
  assign new_n18309_ = ~new_n18306_ & ~new_n18308_;
  assign new_n18310_ = ~\b[3]  & ~new_n18309_;
  assign new_n18311_ = ~new_n17630_ & new_n17632_;
  assign new_n18312_ = ~new_n17628_ & new_n18311_;
  assign new_n18313_ = ~new_n17633_ & ~new_n18312_;
  assign new_n18314_ = \quotient[14]  & new_n18313_;
  assign new_n18315_ = ~new_n17627_ & ~new_n17886_;
  assign new_n18316_ = ~new_n17885_ & new_n18315_;
  assign new_n18317_ = ~new_n18314_ & ~new_n18316_;
  assign new_n18318_ = ~\b[2]  & ~new_n18317_;
  assign new_n18319_ = \b[0]  & \quotient[14] ;
  assign new_n18320_ = \a[14]  & ~new_n18319_;
  assign new_n18321_ = new_n17632_ & \quotient[14] ;
  assign new_n18322_ = ~new_n18320_ & ~new_n18321_;
  assign new_n18323_ = \b[1]  & ~new_n18322_;
  assign new_n18324_ = ~\b[1]  & ~new_n18321_;
  assign new_n18325_ = ~new_n18320_ & new_n18324_;
  assign new_n18326_ = ~new_n18323_ & ~new_n18325_;
  assign new_n18327_ = ~\a[13]  & \b[0] ;
  assign new_n18328_ = ~new_n18326_ & ~new_n18327_;
  assign new_n18329_ = ~\b[1]  & ~new_n18322_;
  assign new_n18330_ = ~new_n18328_ & ~new_n18329_;
  assign new_n18331_ = \b[2]  & ~new_n18316_;
  assign new_n18332_ = ~new_n18314_ & new_n18331_;
  assign new_n18333_ = ~new_n18318_ & ~new_n18332_;
  assign new_n18334_ = ~new_n18330_ & new_n18333_;
  assign new_n18335_ = ~new_n18318_ & ~new_n18334_;
  assign new_n18336_ = \b[3]  & ~new_n18308_;
  assign new_n18337_ = ~new_n18306_ & new_n18336_;
  assign new_n18338_ = ~new_n18310_ & ~new_n18337_;
  assign new_n18339_ = ~new_n18335_ & new_n18338_;
  assign new_n18340_ = ~new_n18310_ & ~new_n18339_;
  assign new_n18341_ = \b[4]  & ~new_n18299_;
  assign new_n18342_ = ~new_n18297_ & new_n18341_;
  assign new_n18343_ = ~new_n18301_ & ~new_n18342_;
  assign new_n18344_ = ~new_n18340_ & new_n18343_;
  assign new_n18345_ = ~new_n18301_ & ~new_n18344_;
  assign new_n18346_ = \b[5]  & ~new_n18290_;
  assign new_n18347_ = ~new_n18288_ & new_n18346_;
  assign new_n18348_ = ~new_n18292_ & ~new_n18347_;
  assign new_n18349_ = ~new_n18345_ & new_n18348_;
  assign new_n18350_ = ~new_n18292_ & ~new_n18349_;
  assign new_n18351_ = \b[6]  & ~new_n18281_;
  assign new_n18352_ = ~new_n18279_ & new_n18351_;
  assign new_n18353_ = ~new_n18283_ & ~new_n18352_;
  assign new_n18354_ = ~new_n18350_ & new_n18353_;
  assign new_n18355_ = ~new_n18283_ & ~new_n18354_;
  assign new_n18356_ = \b[7]  & ~new_n18272_;
  assign new_n18357_ = ~new_n18270_ & new_n18356_;
  assign new_n18358_ = ~new_n18274_ & ~new_n18357_;
  assign new_n18359_ = ~new_n18355_ & new_n18358_;
  assign new_n18360_ = ~new_n18274_ & ~new_n18359_;
  assign new_n18361_ = \b[8]  & ~new_n18263_;
  assign new_n18362_ = ~new_n18261_ & new_n18361_;
  assign new_n18363_ = ~new_n18265_ & ~new_n18362_;
  assign new_n18364_ = ~new_n18360_ & new_n18363_;
  assign new_n18365_ = ~new_n18265_ & ~new_n18364_;
  assign new_n18366_ = \b[9]  & ~new_n18254_;
  assign new_n18367_ = ~new_n18252_ & new_n18366_;
  assign new_n18368_ = ~new_n18256_ & ~new_n18367_;
  assign new_n18369_ = ~new_n18365_ & new_n18368_;
  assign new_n18370_ = ~new_n18256_ & ~new_n18369_;
  assign new_n18371_ = \b[10]  & ~new_n18245_;
  assign new_n18372_ = ~new_n18243_ & new_n18371_;
  assign new_n18373_ = ~new_n18247_ & ~new_n18372_;
  assign new_n18374_ = ~new_n18370_ & new_n18373_;
  assign new_n18375_ = ~new_n18247_ & ~new_n18374_;
  assign new_n18376_ = \b[11]  & ~new_n18236_;
  assign new_n18377_ = ~new_n18234_ & new_n18376_;
  assign new_n18378_ = ~new_n18238_ & ~new_n18377_;
  assign new_n18379_ = ~new_n18375_ & new_n18378_;
  assign new_n18380_ = ~new_n18238_ & ~new_n18379_;
  assign new_n18381_ = \b[12]  & ~new_n18227_;
  assign new_n18382_ = ~new_n18225_ & new_n18381_;
  assign new_n18383_ = ~new_n18229_ & ~new_n18382_;
  assign new_n18384_ = ~new_n18380_ & new_n18383_;
  assign new_n18385_ = ~new_n18229_ & ~new_n18384_;
  assign new_n18386_ = \b[13]  & ~new_n18218_;
  assign new_n18387_ = ~new_n18216_ & new_n18386_;
  assign new_n18388_ = ~new_n18220_ & ~new_n18387_;
  assign new_n18389_ = ~new_n18385_ & new_n18388_;
  assign new_n18390_ = ~new_n18220_ & ~new_n18389_;
  assign new_n18391_ = \b[14]  & ~new_n18209_;
  assign new_n18392_ = ~new_n18207_ & new_n18391_;
  assign new_n18393_ = ~new_n18211_ & ~new_n18392_;
  assign new_n18394_ = ~new_n18390_ & new_n18393_;
  assign new_n18395_ = ~new_n18211_ & ~new_n18394_;
  assign new_n18396_ = \b[15]  & ~new_n18200_;
  assign new_n18397_ = ~new_n18198_ & new_n18396_;
  assign new_n18398_ = ~new_n18202_ & ~new_n18397_;
  assign new_n18399_ = ~new_n18395_ & new_n18398_;
  assign new_n18400_ = ~new_n18202_ & ~new_n18399_;
  assign new_n18401_ = \b[16]  & ~new_n18191_;
  assign new_n18402_ = ~new_n18189_ & new_n18401_;
  assign new_n18403_ = ~new_n18193_ & ~new_n18402_;
  assign new_n18404_ = ~new_n18400_ & new_n18403_;
  assign new_n18405_ = ~new_n18193_ & ~new_n18404_;
  assign new_n18406_ = \b[17]  & ~new_n18182_;
  assign new_n18407_ = ~new_n18180_ & new_n18406_;
  assign new_n18408_ = ~new_n18184_ & ~new_n18407_;
  assign new_n18409_ = ~new_n18405_ & new_n18408_;
  assign new_n18410_ = ~new_n18184_ & ~new_n18409_;
  assign new_n18411_ = \b[18]  & ~new_n18173_;
  assign new_n18412_ = ~new_n18171_ & new_n18411_;
  assign new_n18413_ = ~new_n18175_ & ~new_n18412_;
  assign new_n18414_ = ~new_n18410_ & new_n18413_;
  assign new_n18415_ = ~new_n18175_ & ~new_n18414_;
  assign new_n18416_ = \b[19]  & ~new_n18164_;
  assign new_n18417_ = ~new_n18162_ & new_n18416_;
  assign new_n18418_ = ~new_n18166_ & ~new_n18417_;
  assign new_n18419_ = ~new_n18415_ & new_n18418_;
  assign new_n18420_ = ~new_n18166_ & ~new_n18419_;
  assign new_n18421_ = \b[20]  & ~new_n18155_;
  assign new_n18422_ = ~new_n18153_ & new_n18421_;
  assign new_n18423_ = ~new_n18157_ & ~new_n18422_;
  assign new_n18424_ = ~new_n18420_ & new_n18423_;
  assign new_n18425_ = ~new_n18157_ & ~new_n18424_;
  assign new_n18426_ = \b[21]  & ~new_n18146_;
  assign new_n18427_ = ~new_n18144_ & new_n18426_;
  assign new_n18428_ = ~new_n18148_ & ~new_n18427_;
  assign new_n18429_ = ~new_n18425_ & new_n18428_;
  assign new_n18430_ = ~new_n18148_ & ~new_n18429_;
  assign new_n18431_ = \b[22]  & ~new_n18137_;
  assign new_n18432_ = ~new_n18135_ & new_n18431_;
  assign new_n18433_ = ~new_n18139_ & ~new_n18432_;
  assign new_n18434_ = ~new_n18430_ & new_n18433_;
  assign new_n18435_ = ~new_n18139_ & ~new_n18434_;
  assign new_n18436_ = \b[23]  & ~new_n18128_;
  assign new_n18437_ = ~new_n18126_ & new_n18436_;
  assign new_n18438_ = ~new_n18130_ & ~new_n18437_;
  assign new_n18439_ = ~new_n18435_ & new_n18438_;
  assign new_n18440_ = ~new_n18130_ & ~new_n18439_;
  assign new_n18441_ = \b[24]  & ~new_n18119_;
  assign new_n18442_ = ~new_n18117_ & new_n18441_;
  assign new_n18443_ = ~new_n18121_ & ~new_n18442_;
  assign new_n18444_ = ~new_n18440_ & new_n18443_;
  assign new_n18445_ = ~new_n18121_ & ~new_n18444_;
  assign new_n18446_ = \b[25]  & ~new_n18110_;
  assign new_n18447_ = ~new_n18108_ & new_n18446_;
  assign new_n18448_ = ~new_n18112_ & ~new_n18447_;
  assign new_n18449_ = ~new_n18445_ & new_n18448_;
  assign new_n18450_ = ~new_n18112_ & ~new_n18449_;
  assign new_n18451_ = \b[26]  & ~new_n18101_;
  assign new_n18452_ = ~new_n18099_ & new_n18451_;
  assign new_n18453_ = ~new_n18103_ & ~new_n18452_;
  assign new_n18454_ = ~new_n18450_ & new_n18453_;
  assign new_n18455_ = ~new_n18103_ & ~new_n18454_;
  assign new_n18456_ = \b[27]  & ~new_n18092_;
  assign new_n18457_ = ~new_n18090_ & new_n18456_;
  assign new_n18458_ = ~new_n18094_ & ~new_n18457_;
  assign new_n18459_ = ~new_n18455_ & new_n18458_;
  assign new_n18460_ = ~new_n18094_ & ~new_n18459_;
  assign new_n18461_ = \b[28]  & ~new_n18083_;
  assign new_n18462_ = ~new_n18081_ & new_n18461_;
  assign new_n18463_ = ~new_n18085_ & ~new_n18462_;
  assign new_n18464_ = ~new_n18460_ & new_n18463_;
  assign new_n18465_ = ~new_n18085_ & ~new_n18464_;
  assign new_n18466_ = \b[29]  & ~new_n18074_;
  assign new_n18467_ = ~new_n18072_ & new_n18466_;
  assign new_n18468_ = ~new_n18076_ & ~new_n18467_;
  assign new_n18469_ = ~new_n18465_ & new_n18468_;
  assign new_n18470_ = ~new_n18076_ & ~new_n18469_;
  assign new_n18471_ = \b[30]  & ~new_n18065_;
  assign new_n18472_ = ~new_n18063_ & new_n18471_;
  assign new_n18473_ = ~new_n18067_ & ~new_n18472_;
  assign new_n18474_ = ~new_n18470_ & new_n18473_;
  assign new_n18475_ = ~new_n18067_ & ~new_n18474_;
  assign new_n18476_ = \b[31]  & ~new_n18056_;
  assign new_n18477_ = ~new_n18054_ & new_n18476_;
  assign new_n18478_ = ~new_n18058_ & ~new_n18477_;
  assign new_n18479_ = ~new_n18475_ & new_n18478_;
  assign new_n18480_ = ~new_n18058_ & ~new_n18479_;
  assign new_n18481_ = \b[32]  & ~new_n18047_;
  assign new_n18482_ = ~new_n18045_ & new_n18481_;
  assign new_n18483_ = ~new_n18049_ & ~new_n18482_;
  assign new_n18484_ = ~new_n18480_ & new_n18483_;
  assign new_n18485_ = ~new_n18049_ & ~new_n18484_;
  assign new_n18486_ = \b[33]  & ~new_n18038_;
  assign new_n18487_ = ~new_n18036_ & new_n18486_;
  assign new_n18488_ = ~new_n18040_ & ~new_n18487_;
  assign new_n18489_ = ~new_n18485_ & new_n18488_;
  assign new_n18490_ = ~new_n18040_ & ~new_n18489_;
  assign new_n18491_ = \b[34]  & ~new_n18029_;
  assign new_n18492_ = ~new_n18027_ & new_n18491_;
  assign new_n18493_ = ~new_n18031_ & ~new_n18492_;
  assign new_n18494_ = ~new_n18490_ & new_n18493_;
  assign new_n18495_ = ~new_n18031_ & ~new_n18494_;
  assign new_n18496_ = \b[35]  & ~new_n18020_;
  assign new_n18497_ = ~new_n18018_ & new_n18496_;
  assign new_n18498_ = ~new_n18022_ & ~new_n18497_;
  assign new_n18499_ = ~new_n18495_ & new_n18498_;
  assign new_n18500_ = ~new_n18022_ & ~new_n18499_;
  assign new_n18501_ = \b[36]  & ~new_n18011_;
  assign new_n18502_ = ~new_n18009_ & new_n18501_;
  assign new_n18503_ = ~new_n18013_ & ~new_n18502_;
  assign new_n18504_ = ~new_n18500_ & new_n18503_;
  assign new_n18505_ = ~new_n18013_ & ~new_n18504_;
  assign new_n18506_ = \b[37]  & ~new_n18002_;
  assign new_n18507_ = ~new_n18000_ & new_n18506_;
  assign new_n18508_ = ~new_n18004_ & ~new_n18507_;
  assign new_n18509_ = ~new_n18505_ & new_n18508_;
  assign new_n18510_ = ~new_n18004_ & ~new_n18509_;
  assign new_n18511_ = \b[38]  & ~new_n17993_;
  assign new_n18512_ = ~new_n17991_ & new_n18511_;
  assign new_n18513_ = ~new_n17995_ & ~new_n18512_;
  assign new_n18514_ = ~new_n18510_ & new_n18513_;
  assign new_n18515_ = ~new_n17995_ & ~new_n18514_;
  assign new_n18516_ = \b[39]  & ~new_n17984_;
  assign new_n18517_ = ~new_n17982_ & new_n18516_;
  assign new_n18518_ = ~new_n17986_ & ~new_n18517_;
  assign new_n18519_ = ~new_n18515_ & new_n18518_;
  assign new_n18520_ = ~new_n17986_ & ~new_n18519_;
  assign new_n18521_ = \b[40]  & ~new_n17975_;
  assign new_n18522_ = ~new_n17973_ & new_n18521_;
  assign new_n18523_ = ~new_n17977_ & ~new_n18522_;
  assign new_n18524_ = ~new_n18520_ & new_n18523_;
  assign new_n18525_ = ~new_n17977_ & ~new_n18524_;
  assign new_n18526_ = \b[41]  & ~new_n17966_;
  assign new_n18527_ = ~new_n17964_ & new_n18526_;
  assign new_n18528_ = ~new_n17968_ & ~new_n18527_;
  assign new_n18529_ = ~new_n18525_ & new_n18528_;
  assign new_n18530_ = ~new_n17968_ & ~new_n18529_;
  assign new_n18531_ = \b[42]  & ~new_n17957_;
  assign new_n18532_ = ~new_n17955_ & new_n18531_;
  assign new_n18533_ = ~new_n17959_ & ~new_n18532_;
  assign new_n18534_ = ~new_n18530_ & new_n18533_;
  assign new_n18535_ = ~new_n17959_ & ~new_n18534_;
  assign new_n18536_ = \b[43]  & ~new_n17948_;
  assign new_n18537_ = ~new_n17946_ & new_n18536_;
  assign new_n18538_ = ~new_n17950_ & ~new_n18537_;
  assign new_n18539_ = ~new_n18535_ & new_n18538_;
  assign new_n18540_ = ~new_n17950_ & ~new_n18539_;
  assign new_n18541_ = \b[44]  & ~new_n17939_;
  assign new_n18542_ = ~new_n17937_ & new_n18541_;
  assign new_n18543_ = ~new_n17941_ & ~new_n18542_;
  assign new_n18544_ = ~new_n18540_ & new_n18543_;
  assign new_n18545_ = ~new_n17941_ & ~new_n18544_;
  assign new_n18546_ = \b[45]  & ~new_n17930_;
  assign new_n18547_ = ~new_n17928_ & new_n18546_;
  assign new_n18548_ = ~new_n17932_ & ~new_n18547_;
  assign new_n18549_ = ~new_n18545_ & new_n18548_;
  assign new_n18550_ = ~new_n17932_ & ~new_n18549_;
  assign new_n18551_ = \b[46]  & ~new_n17921_;
  assign new_n18552_ = ~new_n17919_ & new_n18551_;
  assign new_n18553_ = ~new_n17923_ & ~new_n18552_;
  assign new_n18554_ = ~new_n18550_ & new_n18553_;
  assign new_n18555_ = ~new_n17923_ & ~new_n18554_;
  assign new_n18556_ = \b[47]  & ~new_n17912_;
  assign new_n18557_ = ~new_n17910_ & new_n18556_;
  assign new_n18558_ = ~new_n17914_ & ~new_n18557_;
  assign new_n18559_ = ~new_n18555_ & new_n18558_;
  assign new_n18560_ = ~new_n17914_ & ~new_n18559_;
  assign new_n18561_ = \b[48]  & ~new_n17903_;
  assign new_n18562_ = ~new_n17901_ & new_n18561_;
  assign new_n18563_ = ~new_n17905_ & ~new_n18562_;
  assign new_n18564_ = ~new_n18560_ & new_n18563_;
  assign new_n18565_ = ~new_n17905_ & ~new_n18564_;
  assign new_n18566_ = \b[49]  & ~new_n17894_;
  assign new_n18567_ = ~new_n17892_ & new_n18566_;
  assign new_n18568_ = ~new_n17896_ & ~new_n18567_;
  assign new_n18569_ = ~new_n18565_ & new_n18568_;
  assign new_n18570_ = ~new_n17896_ & ~new_n18569_;
  assign new_n18571_ = ~new_n17204_ & ~new_n17880_;
  assign new_n18572_ = ~new_n17878_ & new_n18571_;
  assign new_n18573_ = ~new_n17869_ & new_n18572_;
  assign new_n18574_ = ~new_n17878_ & ~new_n17880_;
  assign new_n18575_ = ~new_n17870_ & ~new_n18574_;
  assign new_n18576_ = ~new_n18573_ & ~new_n18575_;
  assign new_n18577_ = \quotient[14]  & ~new_n18576_;
  assign new_n18578_ = ~new_n17877_ & ~new_n17886_;
  assign new_n18579_ = ~new_n17885_ & new_n18578_;
  assign new_n18580_ = ~new_n18577_ & ~new_n18579_;
  assign new_n18581_ = ~\b[50]  & ~new_n18580_;
  assign new_n18582_ = \b[50]  & ~new_n18579_;
  assign new_n18583_ = ~new_n18577_ & new_n18582_;
  assign new_n18584_ = new_n397_ & new_n399_;
  assign new_n18585_ = new_n407_ & new_n18584_;
  assign new_n18586_ = ~new_n18583_ & new_n18585_;
  assign new_n18587_ = ~new_n18581_ & new_n18586_;
  assign new_n18588_ = ~new_n18570_ & new_n18587_;
  assign new_n18589_ = new_n17882_ & ~new_n18580_;
  assign \quotient[13]  = new_n18588_ | new_n18589_;
  assign new_n18591_ = ~new_n17905_ & new_n18568_;
  assign new_n18592_ = ~new_n18564_ & new_n18591_;
  assign new_n18593_ = ~new_n18565_ & ~new_n18568_;
  assign new_n18594_ = ~new_n18592_ & ~new_n18593_;
  assign new_n18595_ = \quotient[13]  & ~new_n18594_;
  assign new_n18596_ = ~new_n17895_ & ~new_n18589_;
  assign new_n18597_ = ~new_n18588_ & new_n18596_;
  assign new_n18598_ = ~new_n18595_ & ~new_n18597_;
  assign new_n18599_ = ~new_n17896_ & ~new_n18583_;
  assign new_n18600_ = ~new_n18581_ & new_n18599_;
  assign new_n18601_ = ~new_n18569_ & new_n18600_;
  assign new_n18602_ = ~new_n18581_ & ~new_n18583_;
  assign new_n18603_ = ~new_n18570_ & ~new_n18602_;
  assign new_n18604_ = ~new_n18601_ & ~new_n18603_;
  assign new_n18605_ = \quotient[13]  & ~new_n18604_;
  assign new_n18606_ = ~new_n18580_ & ~new_n18589_;
  assign new_n18607_ = ~new_n18588_ & new_n18606_;
  assign new_n18608_ = ~new_n18605_ & ~new_n18607_;
  assign new_n18609_ = ~\b[51]  & ~new_n18608_;
  assign new_n18610_ = ~\b[50]  & ~new_n18598_;
  assign new_n18611_ = ~new_n17914_ & new_n18563_;
  assign new_n18612_ = ~new_n18559_ & new_n18611_;
  assign new_n18613_ = ~new_n18560_ & ~new_n18563_;
  assign new_n18614_ = ~new_n18612_ & ~new_n18613_;
  assign new_n18615_ = \quotient[13]  & ~new_n18614_;
  assign new_n18616_ = ~new_n17904_ & ~new_n18589_;
  assign new_n18617_ = ~new_n18588_ & new_n18616_;
  assign new_n18618_ = ~new_n18615_ & ~new_n18617_;
  assign new_n18619_ = ~\b[49]  & ~new_n18618_;
  assign new_n18620_ = ~new_n17923_ & new_n18558_;
  assign new_n18621_ = ~new_n18554_ & new_n18620_;
  assign new_n18622_ = ~new_n18555_ & ~new_n18558_;
  assign new_n18623_ = ~new_n18621_ & ~new_n18622_;
  assign new_n18624_ = \quotient[13]  & ~new_n18623_;
  assign new_n18625_ = ~new_n17913_ & ~new_n18589_;
  assign new_n18626_ = ~new_n18588_ & new_n18625_;
  assign new_n18627_ = ~new_n18624_ & ~new_n18626_;
  assign new_n18628_ = ~\b[48]  & ~new_n18627_;
  assign new_n18629_ = ~new_n17932_ & new_n18553_;
  assign new_n18630_ = ~new_n18549_ & new_n18629_;
  assign new_n18631_ = ~new_n18550_ & ~new_n18553_;
  assign new_n18632_ = ~new_n18630_ & ~new_n18631_;
  assign new_n18633_ = \quotient[13]  & ~new_n18632_;
  assign new_n18634_ = ~new_n17922_ & ~new_n18589_;
  assign new_n18635_ = ~new_n18588_ & new_n18634_;
  assign new_n18636_ = ~new_n18633_ & ~new_n18635_;
  assign new_n18637_ = ~\b[47]  & ~new_n18636_;
  assign new_n18638_ = ~new_n17941_ & new_n18548_;
  assign new_n18639_ = ~new_n18544_ & new_n18638_;
  assign new_n18640_ = ~new_n18545_ & ~new_n18548_;
  assign new_n18641_ = ~new_n18639_ & ~new_n18640_;
  assign new_n18642_ = \quotient[13]  & ~new_n18641_;
  assign new_n18643_ = ~new_n17931_ & ~new_n18589_;
  assign new_n18644_ = ~new_n18588_ & new_n18643_;
  assign new_n18645_ = ~new_n18642_ & ~new_n18644_;
  assign new_n18646_ = ~\b[46]  & ~new_n18645_;
  assign new_n18647_ = ~new_n17950_ & new_n18543_;
  assign new_n18648_ = ~new_n18539_ & new_n18647_;
  assign new_n18649_ = ~new_n18540_ & ~new_n18543_;
  assign new_n18650_ = ~new_n18648_ & ~new_n18649_;
  assign new_n18651_ = \quotient[13]  & ~new_n18650_;
  assign new_n18652_ = ~new_n17940_ & ~new_n18589_;
  assign new_n18653_ = ~new_n18588_ & new_n18652_;
  assign new_n18654_ = ~new_n18651_ & ~new_n18653_;
  assign new_n18655_ = ~\b[45]  & ~new_n18654_;
  assign new_n18656_ = ~new_n17959_ & new_n18538_;
  assign new_n18657_ = ~new_n18534_ & new_n18656_;
  assign new_n18658_ = ~new_n18535_ & ~new_n18538_;
  assign new_n18659_ = ~new_n18657_ & ~new_n18658_;
  assign new_n18660_ = \quotient[13]  & ~new_n18659_;
  assign new_n18661_ = ~new_n17949_ & ~new_n18589_;
  assign new_n18662_ = ~new_n18588_ & new_n18661_;
  assign new_n18663_ = ~new_n18660_ & ~new_n18662_;
  assign new_n18664_ = ~\b[44]  & ~new_n18663_;
  assign new_n18665_ = ~new_n17968_ & new_n18533_;
  assign new_n18666_ = ~new_n18529_ & new_n18665_;
  assign new_n18667_ = ~new_n18530_ & ~new_n18533_;
  assign new_n18668_ = ~new_n18666_ & ~new_n18667_;
  assign new_n18669_ = \quotient[13]  & ~new_n18668_;
  assign new_n18670_ = ~new_n17958_ & ~new_n18589_;
  assign new_n18671_ = ~new_n18588_ & new_n18670_;
  assign new_n18672_ = ~new_n18669_ & ~new_n18671_;
  assign new_n18673_ = ~\b[43]  & ~new_n18672_;
  assign new_n18674_ = ~new_n17977_ & new_n18528_;
  assign new_n18675_ = ~new_n18524_ & new_n18674_;
  assign new_n18676_ = ~new_n18525_ & ~new_n18528_;
  assign new_n18677_ = ~new_n18675_ & ~new_n18676_;
  assign new_n18678_ = \quotient[13]  & ~new_n18677_;
  assign new_n18679_ = ~new_n17967_ & ~new_n18589_;
  assign new_n18680_ = ~new_n18588_ & new_n18679_;
  assign new_n18681_ = ~new_n18678_ & ~new_n18680_;
  assign new_n18682_ = ~\b[42]  & ~new_n18681_;
  assign new_n18683_ = ~new_n17986_ & new_n18523_;
  assign new_n18684_ = ~new_n18519_ & new_n18683_;
  assign new_n18685_ = ~new_n18520_ & ~new_n18523_;
  assign new_n18686_ = ~new_n18684_ & ~new_n18685_;
  assign new_n18687_ = \quotient[13]  & ~new_n18686_;
  assign new_n18688_ = ~new_n17976_ & ~new_n18589_;
  assign new_n18689_ = ~new_n18588_ & new_n18688_;
  assign new_n18690_ = ~new_n18687_ & ~new_n18689_;
  assign new_n18691_ = ~\b[41]  & ~new_n18690_;
  assign new_n18692_ = ~new_n17995_ & new_n18518_;
  assign new_n18693_ = ~new_n18514_ & new_n18692_;
  assign new_n18694_ = ~new_n18515_ & ~new_n18518_;
  assign new_n18695_ = ~new_n18693_ & ~new_n18694_;
  assign new_n18696_ = \quotient[13]  & ~new_n18695_;
  assign new_n18697_ = ~new_n17985_ & ~new_n18589_;
  assign new_n18698_ = ~new_n18588_ & new_n18697_;
  assign new_n18699_ = ~new_n18696_ & ~new_n18698_;
  assign new_n18700_ = ~\b[40]  & ~new_n18699_;
  assign new_n18701_ = ~new_n18004_ & new_n18513_;
  assign new_n18702_ = ~new_n18509_ & new_n18701_;
  assign new_n18703_ = ~new_n18510_ & ~new_n18513_;
  assign new_n18704_ = ~new_n18702_ & ~new_n18703_;
  assign new_n18705_ = \quotient[13]  & ~new_n18704_;
  assign new_n18706_ = ~new_n17994_ & ~new_n18589_;
  assign new_n18707_ = ~new_n18588_ & new_n18706_;
  assign new_n18708_ = ~new_n18705_ & ~new_n18707_;
  assign new_n18709_ = ~\b[39]  & ~new_n18708_;
  assign new_n18710_ = ~new_n18013_ & new_n18508_;
  assign new_n18711_ = ~new_n18504_ & new_n18710_;
  assign new_n18712_ = ~new_n18505_ & ~new_n18508_;
  assign new_n18713_ = ~new_n18711_ & ~new_n18712_;
  assign new_n18714_ = \quotient[13]  & ~new_n18713_;
  assign new_n18715_ = ~new_n18003_ & ~new_n18589_;
  assign new_n18716_ = ~new_n18588_ & new_n18715_;
  assign new_n18717_ = ~new_n18714_ & ~new_n18716_;
  assign new_n18718_ = ~\b[38]  & ~new_n18717_;
  assign new_n18719_ = ~new_n18022_ & new_n18503_;
  assign new_n18720_ = ~new_n18499_ & new_n18719_;
  assign new_n18721_ = ~new_n18500_ & ~new_n18503_;
  assign new_n18722_ = ~new_n18720_ & ~new_n18721_;
  assign new_n18723_ = \quotient[13]  & ~new_n18722_;
  assign new_n18724_ = ~new_n18012_ & ~new_n18589_;
  assign new_n18725_ = ~new_n18588_ & new_n18724_;
  assign new_n18726_ = ~new_n18723_ & ~new_n18725_;
  assign new_n18727_ = ~\b[37]  & ~new_n18726_;
  assign new_n18728_ = ~new_n18031_ & new_n18498_;
  assign new_n18729_ = ~new_n18494_ & new_n18728_;
  assign new_n18730_ = ~new_n18495_ & ~new_n18498_;
  assign new_n18731_ = ~new_n18729_ & ~new_n18730_;
  assign new_n18732_ = \quotient[13]  & ~new_n18731_;
  assign new_n18733_ = ~new_n18021_ & ~new_n18589_;
  assign new_n18734_ = ~new_n18588_ & new_n18733_;
  assign new_n18735_ = ~new_n18732_ & ~new_n18734_;
  assign new_n18736_ = ~\b[36]  & ~new_n18735_;
  assign new_n18737_ = ~new_n18040_ & new_n18493_;
  assign new_n18738_ = ~new_n18489_ & new_n18737_;
  assign new_n18739_ = ~new_n18490_ & ~new_n18493_;
  assign new_n18740_ = ~new_n18738_ & ~new_n18739_;
  assign new_n18741_ = \quotient[13]  & ~new_n18740_;
  assign new_n18742_ = ~new_n18030_ & ~new_n18589_;
  assign new_n18743_ = ~new_n18588_ & new_n18742_;
  assign new_n18744_ = ~new_n18741_ & ~new_n18743_;
  assign new_n18745_ = ~\b[35]  & ~new_n18744_;
  assign new_n18746_ = ~new_n18049_ & new_n18488_;
  assign new_n18747_ = ~new_n18484_ & new_n18746_;
  assign new_n18748_ = ~new_n18485_ & ~new_n18488_;
  assign new_n18749_ = ~new_n18747_ & ~new_n18748_;
  assign new_n18750_ = \quotient[13]  & ~new_n18749_;
  assign new_n18751_ = ~new_n18039_ & ~new_n18589_;
  assign new_n18752_ = ~new_n18588_ & new_n18751_;
  assign new_n18753_ = ~new_n18750_ & ~new_n18752_;
  assign new_n18754_ = ~\b[34]  & ~new_n18753_;
  assign new_n18755_ = ~new_n18058_ & new_n18483_;
  assign new_n18756_ = ~new_n18479_ & new_n18755_;
  assign new_n18757_ = ~new_n18480_ & ~new_n18483_;
  assign new_n18758_ = ~new_n18756_ & ~new_n18757_;
  assign new_n18759_ = \quotient[13]  & ~new_n18758_;
  assign new_n18760_ = ~new_n18048_ & ~new_n18589_;
  assign new_n18761_ = ~new_n18588_ & new_n18760_;
  assign new_n18762_ = ~new_n18759_ & ~new_n18761_;
  assign new_n18763_ = ~\b[33]  & ~new_n18762_;
  assign new_n18764_ = ~new_n18067_ & new_n18478_;
  assign new_n18765_ = ~new_n18474_ & new_n18764_;
  assign new_n18766_ = ~new_n18475_ & ~new_n18478_;
  assign new_n18767_ = ~new_n18765_ & ~new_n18766_;
  assign new_n18768_ = \quotient[13]  & ~new_n18767_;
  assign new_n18769_ = ~new_n18057_ & ~new_n18589_;
  assign new_n18770_ = ~new_n18588_ & new_n18769_;
  assign new_n18771_ = ~new_n18768_ & ~new_n18770_;
  assign new_n18772_ = ~\b[32]  & ~new_n18771_;
  assign new_n18773_ = ~new_n18076_ & new_n18473_;
  assign new_n18774_ = ~new_n18469_ & new_n18773_;
  assign new_n18775_ = ~new_n18470_ & ~new_n18473_;
  assign new_n18776_ = ~new_n18774_ & ~new_n18775_;
  assign new_n18777_ = \quotient[13]  & ~new_n18776_;
  assign new_n18778_ = ~new_n18066_ & ~new_n18589_;
  assign new_n18779_ = ~new_n18588_ & new_n18778_;
  assign new_n18780_ = ~new_n18777_ & ~new_n18779_;
  assign new_n18781_ = ~\b[31]  & ~new_n18780_;
  assign new_n18782_ = ~new_n18085_ & new_n18468_;
  assign new_n18783_ = ~new_n18464_ & new_n18782_;
  assign new_n18784_ = ~new_n18465_ & ~new_n18468_;
  assign new_n18785_ = ~new_n18783_ & ~new_n18784_;
  assign new_n18786_ = \quotient[13]  & ~new_n18785_;
  assign new_n18787_ = ~new_n18075_ & ~new_n18589_;
  assign new_n18788_ = ~new_n18588_ & new_n18787_;
  assign new_n18789_ = ~new_n18786_ & ~new_n18788_;
  assign new_n18790_ = ~\b[30]  & ~new_n18789_;
  assign new_n18791_ = ~new_n18094_ & new_n18463_;
  assign new_n18792_ = ~new_n18459_ & new_n18791_;
  assign new_n18793_ = ~new_n18460_ & ~new_n18463_;
  assign new_n18794_ = ~new_n18792_ & ~new_n18793_;
  assign new_n18795_ = \quotient[13]  & ~new_n18794_;
  assign new_n18796_ = ~new_n18084_ & ~new_n18589_;
  assign new_n18797_ = ~new_n18588_ & new_n18796_;
  assign new_n18798_ = ~new_n18795_ & ~new_n18797_;
  assign new_n18799_ = ~\b[29]  & ~new_n18798_;
  assign new_n18800_ = ~new_n18103_ & new_n18458_;
  assign new_n18801_ = ~new_n18454_ & new_n18800_;
  assign new_n18802_ = ~new_n18455_ & ~new_n18458_;
  assign new_n18803_ = ~new_n18801_ & ~new_n18802_;
  assign new_n18804_ = \quotient[13]  & ~new_n18803_;
  assign new_n18805_ = ~new_n18093_ & ~new_n18589_;
  assign new_n18806_ = ~new_n18588_ & new_n18805_;
  assign new_n18807_ = ~new_n18804_ & ~new_n18806_;
  assign new_n18808_ = ~\b[28]  & ~new_n18807_;
  assign new_n18809_ = ~new_n18112_ & new_n18453_;
  assign new_n18810_ = ~new_n18449_ & new_n18809_;
  assign new_n18811_ = ~new_n18450_ & ~new_n18453_;
  assign new_n18812_ = ~new_n18810_ & ~new_n18811_;
  assign new_n18813_ = \quotient[13]  & ~new_n18812_;
  assign new_n18814_ = ~new_n18102_ & ~new_n18589_;
  assign new_n18815_ = ~new_n18588_ & new_n18814_;
  assign new_n18816_ = ~new_n18813_ & ~new_n18815_;
  assign new_n18817_ = ~\b[27]  & ~new_n18816_;
  assign new_n18818_ = ~new_n18121_ & new_n18448_;
  assign new_n18819_ = ~new_n18444_ & new_n18818_;
  assign new_n18820_ = ~new_n18445_ & ~new_n18448_;
  assign new_n18821_ = ~new_n18819_ & ~new_n18820_;
  assign new_n18822_ = \quotient[13]  & ~new_n18821_;
  assign new_n18823_ = ~new_n18111_ & ~new_n18589_;
  assign new_n18824_ = ~new_n18588_ & new_n18823_;
  assign new_n18825_ = ~new_n18822_ & ~new_n18824_;
  assign new_n18826_ = ~\b[26]  & ~new_n18825_;
  assign new_n18827_ = ~new_n18130_ & new_n18443_;
  assign new_n18828_ = ~new_n18439_ & new_n18827_;
  assign new_n18829_ = ~new_n18440_ & ~new_n18443_;
  assign new_n18830_ = ~new_n18828_ & ~new_n18829_;
  assign new_n18831_ = \quotient[13]  & ~new_n18830_;
  assign new_n18832_ = ~new_n18120_ & ~new_n18589_;
  assign new_n18833_ = ~new_n18588_ & new_n18832_;
  assign new_n18834_ = ~new_n18831_ & ~new_n18833_;
  assign new_n18835_ = ~\b[25]  & ~new_n18834_;
  assign new_n18836_ = ~new_n18139_ & new_n18438_;
  assign new_n18837_ = ~new_n18434_ & new_n18836_;
  assign new_n18838_ = ~new_n18435_ & ~new_n18438_;
  assign new_n18839_ = ~new_n18837_ & ~new_n18838_;
  assign new_n18840_ = \quotient[13]  & ~new_n18839_;
  assign new_n18841_ = ~new_n18129_ & ~new_n18589_;
  assign new_n18842_ = ~new_n18588_ & new_n18841_;
  assign new_n18843_ = ~new_n18840_ & ~new_n18842_;
  assign new_n18844_ = ~\b[24]  & ~new_n18843_;
  assign new_n18845_ = ~new_n18148_ & new_n18433_;
  assign new_n18846_ = ~new_n18429_ & new_n18845_;
  assign new_n18847_ = ~new_n18430_ & ~new_n18433_;
  assign new_n18848_ = ~new_n18846_ & ~new_n18847_;
  assign new_n18849_ = \quotient[13]  & ~new_n18848_;
  assign new_n18850_ = ~new_n18138_ & ~new_n18589_;
  assign new_n18851_ = ~new_n18588_ & new_n18850_;
  assign new_n18852_ = ~new_n18849_ & ~new_n18851_;
  assign new_n18853_ = ~\b[23]  & ~new_n18852_;
  assign new_n18854_ = ~new_n18157_ & new_n18428_;
  assign new_n18855_ = ~new_n18424_ & new_n18854_;
  assign new_n18856_ = ~new_n18425_ & ~new_n18428_;
  assign new_n18857_ = ~new_n18855_ & ~new_n18856_;
  assign new_n18858_ = \quotient[13]  & ~new_n18857_;
  assign new_n18859_ = ~new_n18147_ & ~new_n18589_;
  assign new_n18860_ = ~new_n18588_ & new_n18859_;
  assign new_n18861_ = ~new_n18858_ & ~new_n18860_;
  assign new_n18862_ = ~\b[22]  & ~new_n18861_;
  assign new_n18863_ = ~new_n18166_ & new_n18423_;
  assign new_n18864_ = ~new_n18419_ & new_n18863_;
  assign new_n18865_ = ~new_n18420_ & ~new_n18423_;
  assign new_n18866_ = ~new_n18864_ & ~new_n18865_;
  assign new_n18867_ = \quotient[13]  & ~new_n18866_;
  assign new_n18868_ = ~new_n18156_ & ~new_n18589_;
  assign new_n18869_ = ~new_n18588_ & new_n18868_;
  assign new_n18870_ = ~new_n18867_ & ~new_n18869_;
  assign new_n18871_ = ~\b[21]  & ~new_n18870_;
  assign new_n18872_ = ~new_n18175_ & new_n18418_;
  assign new_n18873_ = ~new_n18414_ & new_n18872_;
  assign new_n18874_ = ~new_n18415_ & ~new_n18418_;
  assign new_n18875_ = ~new_n18873_ & ~new_n18874_;
  assign new_n18876_ = \quotient[13]  & ~new_n18875_;
  assign new_n18877_ = ~new_n18165_ & ~new_n18589_;
  assign new_n18878_ = ~new_n18588_ & new_n18877_;
  assign new_n18879_ = ~new_n18876_ & ~new_n18878_;
  assign new_n18880_ = ~\b[20]  & ~new_n18879_;
  assign new_n18881_ = ~new_n18184_ & new_n18413_;
  assign new_n18882_ = ~new_n18409_ & new_n18881_;
  assign new_n18883_ = ~new_n18410_ & ~new_n18413_;
  assign new_n18884_ = ~new_n18882_ & ~new_n18883_;
  assign new_n18885_ = \quotient[13]  & ~new_n18884_;
  assign new_n18886_ = ~new_n18174_ & ~new_n18589_;
  assign new_n18887_ = ~new_n18588_ & new_n18886_;
  assign new_n18888_ = ~new_n18885_ & ~new_n18887_;
  assign new_n18889_ = ~\b[19]  & ~new_n18888_;
  assign new_n18890_ = ~new_n18193_ & new_n18408_;
  assign new_n18891_ = ~new_n18404_ & new_n18890_;
  assign new_n18892_ = ~new_n18405_ & ~new_n18408_;
  assign new_n18893_ = ~new_n18891_ & ~new_n18892_;
  assign new_n18894_ = \quotient[13]  & ~new_n18893_;
  assign new_n18895_ = ~new_n18183_ & ~new_n18589_;
  assign new_n18896_ = ~new_n18588_ & new_n18895_;
  assign new_n18897_ = ~new_n18894_ & ~new_n18896_;
  assign new_n18898_ = ~\b[18]  & ~new_n18897_;
  assign new_n18899_ = ~new_n18202_ & new_n18403_;
  assign new_n18900_ = ~new_n18399_ & new_n18899_;
  assign new_n18901_ = ~new_n18400_ & ~new_n18403_;
  assign new_n18902_ = ~new_n18900_ & ~new_n18901_;
  assign new_n18903_ = \quotient[13]  & ~new_n18902_;
  assign new_n18904_ = ~new_n18192_ & ~new_n18589_;
  assign new_n18905_ = ~new_n18588_ & new_n18904_;
  assign new_n18906_ = ~new_n18903_ & ~new_n18905_;
  assign new_n18907_ = ~\b[17]  & ~new_n18906_;
  assign new_n18908_ = ~new_n18211_ & new_n18398_;
  assign new_n18909_ = ~new_n18394_ & new_n18908_;
  assign new_n18910_ = ~new_n18395_ & ~new_n18398_;
  assign new_n18911_ = ~new_n18909_ & ~new_n18910_;
  assign new_n18912_ = \quotient[13]  & ~new_n18911_;
  assign new_n18913_ = ~new_n18201_ & ~new_n18589_;
  assign new_n18914_ = ~new_n18588_ & new_n18913_;
  assign new_n18915_ = ~new_n18912_ & ~new_n18914_;
  assign new_n18916_ = ~\b[16]  & ~new_n18915_;
  assign new_n18917_ = ~new_n18220_ & new_n18393_;
  assign new_n18918_ = ~new_n18389_ & new_n18917_;
  assign new_n18919_ = ~new_n18390_ & ~new_n18393_;
  assign new_n18920_ = ~new_n18918_ & ~new_n18919_;
  assign new_n18921_ = \quotient[13]  & ~new_n18920_;
  assign new_n18922_ = ~new_n18210_ & ~new_n18589_;
  assign new_n18923_ = ~new_n18588_ & new_n18922_;
  assign new_n18924_ = ~new_n18921_ & ~new_n18923_;
  assign new_n18925_ = ~\b[15]  & ~new_n18924_;
  assign new_n18926_ = ~new_n18229_ & new_n18388_;
  assign new_n18927_ = ~new_n18384_ & new_n18926_;
  assign new_n18928_ = ~new_n18385_ & ~new_n18388_;
  assign new_n18929_ = ~new_n18927_ & ~new_n18928_;
  assign new_n18930_ = \quotient[13]  & ~new_n18929_;
  assign new_n18931_ = ~new_n18219_ & ~new_n18589_;
  assign new_n18932_ = ~new_n18588_ & new_n18931_;
  assign new_n18933_ = ~new_n18930_ & ~new_n18932_;
  assign new_n18934_ = ~\b[14]  & ~new_n18933_;
  assign new_n18935_ = ~new_n18238_ & new_n18383_;
  assign new_n18936_ = ~new_n18379_ & new_n18935_;
  assign new_n18937_ = ~new_n18380_ & ~new_n18383_;
  assign new_n18938_ = ~new_n18936_ & ~new_n18937_;
  assign new_n18939_ = \quotient[13]  & ~new_n18938_;
  assign new_n18940_ = ~new_n18228_ & ~new_n18589_;
  assign new_n18941_ = ~new_n18588_ & new_n18940_;
  assign new_n18942_ = ~new_n18939_ & ~new_n18941_;
  assign new_n18943_ = ~\b[13]  & ~new_n18942_;
  assign new_n18944_ = ~new_n18247_ & new_n18378_;
  assign new_n18945_ = ~new_n18374_ & new_n18944_;
  assign new_n18946_ = ~new_n18375_ & ~new_n18378_;
  assign new_n18947_ = ~new_n18945_ & ~new_n18946_;
  assign new_n18948_ = \quotient[13]  & ~new_n18947_;
  assign new_n18949_ = ~new_n18237_ & ~new_n18589_;
  assign new_n18950_ = ~new_n18588_ & new_n18949_;
  assign new_n18951_ = ~new_n18948_ & ~new_n18950_;
  assign new_n18952_ = ~\b[12]  & ~new_n18951_;
  assign new_n18953_ = ~new_n18256_ & new_n18373_;
  assign new_n18954_ = ~new_n18369_ & new_n18953_;
  assign new_n18955_ = ~new_n18370_ & ~new_n18373_;
  assign new_n18956_ = ~new_n18954_ & ~new_n18955_;
  assign new_n18957_ = \quotient[13]  & ~new_n18956_;
  assign new_n18958_ = ~new_n18246_ & ~new_n18589_;
  assign new_n18959_ = ~new_n18588_ & new_n18958_;
  assign new_n18960_ = ~new_n18957_ & ~new_n18959_;
  assign new_n18961_ = ~\b[11]  & ~new_n18960_;
  assign new_n18962_ = ~new_n18265_ & new_n18368_;
  assign new_n18963_ = ~new_n18364_ & new_n18962_;
  assign new_n18964_ = ~new_n18365_ & ~new_n18368_;
  assign new_n18965_ = ~new_n18963_ & ~new_n18964_;
  assign new_n18966_ = \quotient[13]  & ~new_n18965_;
  assign new_n18967_ = ~new_n18255_ & ~new_n18589_;
  assign new_n18968_ = ~new_n18588_ & new_n18967_;
  assign new_n18969_ = ~new_n18966_ & ~new_n18968_;
  assign new_n18970_ = ~\b[10]  & ~new_n18969_;
  assign new_n18971_ = ~new_n18274_ & new_n18363_;
  assign new_n18972_ = ~new_n18359_ & new_n18971_;
  assign new_n18973_ = ~new_n18360_ & ~new_n18363_;
  assign new_n18974_ = ~new_n18972_ & ~new_n18973_;
  assign new_n18975_ = \quotient[13]  & ~new_n18974_;
  assign new_n18976_ = ~new_n18264_ & ~new_n18589_;
  assign new_n18977_ = ~new_n18588_ & new_n18976_;
  assign new_n18978_ = ~new_n18975_ & ~new_n18977_;
  assign new_n18979_ = ~\b[9]  & ~new_n18978_;
  assign new_n18980_ = ~new_n18283_ & new_n18358_;
  assign new_n18981_ = ~new_n18354_ & new_n18980_;
  assign new_n18982_ = ~new_n18355_ & ~new_n18358_;
  assign new_n18983_ = ~new_n18981_ & ~new_n18982_;
  assign new_n18984_ = \quotient[13]  & ~new_n18983_;
  assign new_n18985_ = ~new_n18273_ & ~new_n18589_;
  assign new_n18986_ = ~new_n18588_ & new_n18985_;
  assign new_n18987_ = ~new_n18984_ & ~new_n18986_;
  assign new_n18988_ = ~\b[8]  & ~new_n18987_;
  assign new_n18989_ = ~new_n18292_ & new_n18353_;
  assign new_n18990_ = ~new_n18349_ & new_n18989_;
  assign new_n18991_ = ~new_n18350_ & ~new_n18353_;
  assign new_n18992_ = ~new_n18990_ & ~new_n18991_;
  assign new_n18993_ = \quotient[13]  & ~new_n18992_;
  assign new_n18994_ = ~new_n18282_ & ~new_n18589_;
  assign new_n18995_ = ~new_n18588_ & new_n18994_;
  assign new_n18996_ = ~new_n18993_ & ~new_n18995_;
  assign new_n18997_ = ~\b[7]  & ~new_n18996_;
  assign new_n18998_ = ~new_n18301_ & new_n18348_;
  assign new_n18999_ = ~new_n18344_ & new_n18998_;
  assign new_n19000_ = ~new_n18345_ & ~new_n18348_;
  assign new_n19001_ = ~new_n18999_ & ~new_n19000_;
  assign new_n19002_ = \quotient[13]  & ~new_n19001_;
  assign new_n19003_ = ~new_n18291_ & ~new_n18589_;
  assign new_n19004_ = ~new_n18588_ & new_n19003_;
  assign new_n19005_ = ~new_n19002_ & ~new_n19004_;
  assign new_n19006_ = ~\b[6]  & ~new_n19005_;
  assign new_n19007_ = ~new_n18310_ & new_n18343_;
  assign new_n19008_ = ~new_n18339_ & new_n19007_;
  assign new_n19009_ = ~new_n18340_ & ~new_n18343_;
  assign new_n19010_ = ~new_n19008_ & ~new_n19009_;
  assign new_n19011_ = \quotient[13]  & ~new_n19010_;
  assign new_n19012_ = ~new_n18300_ & ~new_n18589_;
  assign new_n19013_ = ~new_n18588_ & new_n19012_;
  assign new_n19014_ = ~new_n19011_ & ~new_n19013_;
  assign new_n19015_ = ~\b[5]  & ~new_n19014_;
  assign new_n19016_ = ~new_n18318_ & new_n18338_;
  assign new_n19017_ = ~new_n18334_ & new_n19016_;
  assign new_n19018_ = ~new_n18335_ & ~new_n18338_;
  assign new_n19019_ = ~new_n19017_ & ~new_n19018_;
  assign new_n19020_ = \quotient[13]  & ~new_n19019_;
  assign new_n19021_ = ~new_n18309_ & ~new_n18589_;
  assign new_n19022_ = ~new_n18588_ & new_n19021_;
  assign new_n19023_ = ~new_n19020_ & ~new_n19022_;
  assign new_n19024_ = ~\b[4]  & ~new_n19023_;
  assign new_n19025_ = ~new_n18329_ & new_n18333_;
  assign new_n19026_ = ~new_n18328_ & new_n19025_;
  assign new_n19027_ = ~new_n18330_ & ~new_n18333_;
  assign new_n19028_ = ~new_n19026_ & ~new_n19027_;
  assign new_n19029_ = \quotient[13]  & ~new_n19028_;
  assign new_n19030_ = ~new_n18317_ & ~new_n18589_;
  assign new_n19031_ = ~new_n18588_ & new_n19030_;
  assign new_n19032_ = ~new_n19029_ & ~new_n19031_;
  assign new_n19033_ = ~\b[3]  & ~new_n19032_;
  assign new_n19034_ = ~new_n18325_ & new_n18327_;
  assign new_n19035_ = ~new_n18323_ & new_n19034_;
  assign new_n19036_ = ~new_n18328_ & ~new_n19035_;
  assign new_n19037_ = \quotient[13]  & new_n19036_;
  assign new_n19038_ = ~new_n18322_ & ~new_n18589_;
  assign new_n19039_ = ~new_n18588_ & new_n19038_;
  assign new_n19040_ = ~new_n19037_ & ~new_n19039_;
  assign new_n19041_ = ~\b[2]  & ~new_n19040_;
  assign new_n19042_ = \b[0]  & \quotient[13] ;
  assign new_n19043_ = \a[13]  & ~new_n19042_;
  assign new_n19044_ = new_n18327_ & \quotient[13] ;
  assign new_n19045_ = ~new_n19043_ & ~new_n19044_;
  assign new_n19046_ = \b[1]  & ~new_n19045_;
  assign new_n19047_ = ~\b[1]  & ~new_n19044_;
  assign new_n19048_ = ~new_n19043_ & new_n19047_;
  assign new_n19049_ = ~new_n19046_ & ~new_n19048_;
  assign new_n19050_ = ~\a[12]  & \b[0] ;
  assign new_n19051_ = ~new_n19049_ & ~new_n19050_;
  assign new_n19052_ = ~\b[1]  & ~new_n19045_;
  assign new_n19053_ = ~new_n19051_ & ~new_n19052_;
  assign new_n19054_ = \b[2]  & ~new_n19039_;
  assign new_n19055_ = ~new_n19037_ & new_n19054_;
  assign new_n19056_ = ~new_n19041_ & ~new_n19055_;
  assign new_n19057_ = ~new_n19053_ & new_n19056_;
  assign new_n19058_ = ~new_n19041_ & ~new_n19057_;
  assign new_n19059_ = \b[3]  & ~new_n19031_;
  assign new_n19060_ = ~new_n19029_ & new_n19059_;
  assign new_n19061_ = ~new_n19033_ & ~new_n19060_;
  assign new_n19062_ = ~new_n19058_ & new_n19061_;
  assign new_n19063_ = ~new_n19033_ & ~new_n19062_;
  assign new_n19064_ = \b[4]  & ~new_n19022_;
  assign new_n19065_ = ~new_n19020_ & new_n19064_;
  assign new_n19066_ = ~new_n19024_ & ~new_n19065_;
  assign new_n19067_ = ~new_n19063_ & new_n19066_;
  assign new_n19068_ = ~new_n19024_ & ~new_n19067_;
  assign new_n19069_ = \b[5]  & ~new_n19013_;
  assign new_n19070_ = ~new_n19011_ & new_n19069_;
  assign new_n19071_ = ~new_n19015_ & ~new_n19070_;
  assign new_n19072_ = ~new_n19068_ & new_n19071_;
  assign new_n19073_ = ~new_n19015_ & ~new_n19072_;
  assign new_n19074_ = \b[6]  & ~new_n19004_;
  assign new_n19075_ = ~new_n19002_ & new_n19074_;
  assign new_n19076_ = ~new_n19006_ & ~new_n19075_;
  assign new_n19077_ = ~new_n19073_ & new_n19076_;
  assign new_n19078_ = ~new_n19006_ & ~new_n19077_;
  assign new_n19079_ = \b[7]  & ~new_n18995_;
  assign new_n19080_ = ~new_n18993_ & new_n19079_;
  assign new_n19081_ = ~new_n18997_ & ~new_n19080_;
  assign new_n19082_ = ~new_n19078_ & new_n19081_;
  assign new_n19083_ = ~new_n18997_ & ~new_n19082_;
  assign new_n19084_ = \b[8]  & ~new_n18986_;
  assign new_n19085_ = ~new_n18984_ & new_n19084_;
  assign new_n19086_ = ~new_n18988_ & ~new_n19085_;
  assign new_n19087_ = ~new_n19083_ & new_n19086_;
  assign new_n19088_ = ~new_n18988_ & ~new_n19087_;
  assign new_n19089_ = \b[9]  & ~new_n18977_;
  assign new_n19090_ = ~new_n18975_ & new_n19089_;
  assign new_n19091_ = ~new_n18979_ & ~new_n19090_;
  assign new_n19092_ = ~new_n19088_ & new_n19091_;
  assign new_n19093_ = ~new_n18979_ & ~new_n19092_;
  assign new_n19094_ = \b[10]  & ~new_n18968_;
  assign new_n19095_ = ~new_n18966_ & new_n19094_;
  assign new_n19096_ = ~new_n18970_ & ~new_n19095_;
  assign new_n19097_ = ~new_n19093_ & new_n19096_;
  assign new_n19098_ = ~new_n18970_ & ~new_n19097_;
  assign new_n19099_ = \b[11]  & ~new_n18959_;
  assign new_n19100_ = ~new_n18957_ & new_n19099_;
  assign new_n19101_ = ~new_n18961_ & ~new_n19100_;
  assign new_n19102_ = ~new_n19098_ & new_n19101_;
  assign new_n19103_ = ~new_n18961_ & ~new_n19102_;
  assign new_n19104_ = \b[12]  & ~new_n18950_;
  assign new_n19105_ = ~new_n18948_ & new_n19104_;
  assign new_n19106_ = ~new_n18952_ & ~new_n19105_;
  assign new_n19107_ = ~new_n19103_ & new_n19106_;
  assign new_n19108_ = ~new_n18952_ & ~new_n19107_;
  assign new_n19109_ = \b[13]  & ~new_n18941_;
  assign new_n19110_ = ~new_n18939_ & new_n19109_;
  assign new_n19111_ = ~new_n18943_ & ~new_n19110_;
  assign new_n19112_ = ~new_n19108_ & new_n19111_;
  assign new_n19113_ = ~new_n18943_ & ~new_n19112_;
  assign new_n19114_ = \b[14]  & ~new_n18932_;
  assign new_n19115_ = ~new_n18930_ & new_n19114_;
  assign new_n19116_ = ~new_n18934_ & ~new_n19115_;
  assign new_n19117_ = ~new_n19113_ & new_n19116_;
  assign new_n19118_ = ~new_n18934_ & ~new_n19117_;
  assign new_n19119_ = \b[15]  & ~new_n18923_;
  assign new_n19120_ = ~new_n18921_ & new_n19119_;
  assign new_n19121_ = ~new_n18925_ & ~new_n19120_;
  assign new_n19122_ = ~new_n19118_ & new_n19121_;
  assign new_n19123_ = ~new_n18925_ & ~new_n19122_;
  assign new_n19124_ = \b[16]  & ~new_n18914_;
  assign new_n19125_ = ~new_n18912_ & new_n19124_;
  assign new_n19126_ = ~new_n18916_ & ~new_n19125_;
  assign new_n19127_ = ~new_n19123_ & new_n19126_;
  assign new_n19128_ = ~new_n18916_ & ~new_n19127_;
  assign new_n19129_ = \b[17]  & ~new_n18905_;
  assign new_n19130_ = ~new_n18903_ & new_n19129_;
  assign new_n19131_ = ~new_n18907_ & ~new_n19130_;
  assign new_n19132_ = ~new_n19128_ & new_n19131_;
  assign new_n19133_ = ~new_n18907_ & ~new_n19132_;
  assign new_n19134_ = \b[18]  & ~new_n18896_;
  assign new_n19135_ = ~new_n18894_ & new_n19134_;
  assign new_n19136_ = ~new_n18898_ & ~new_n19135_;
  assign new_n19137_ = ~new_n19133_ & new_n19136_;
  assign new_n19138_ = ~new_n18898_ & ~new_n19137_;
  assign new_n19139_ = \b[19]  & ~new_n18887_;
  assign new_n19140_ = ~new_n18885_ & new_n19139_;
  assign new_n19141_ = ~new_n18889_ & ~new_n19140_;
  assign new_n19142_ = ~new_n19138_ & new_n19141_;
  assign new_n19143_ = ~new_n18889_ & ~new_n19142_;
  assign new_n19144_ = \b[20]  & ~new_n18878_;
  assign new_n19145_ = ~new_n18876_ & new_n19144_;
  assign new_n19146_ = ~new_n18880_ & ~new_n19145_;
  assign new_n19147_ = ~new_n19143_ & new_n19146_;
  assign new_n19148_ = ~new_n18880_ & ~new_n19147_;
  assign new_n19149_ = \b[21]  & ~new_n18869_;
  assign new_n19150_ = ~new_n18867_ & new_n19149_;
  assign new_n19151_ = ~new_n18871_ & ~new_n19150_;
  assign new_n19152_ = ~new_n19148_ & new_n19151_;
  assign new_n19153_ = ~new_n18871_ & ~new_n19152_;
  assign new_n19154_ = \b[22]  & ~new_n18860_;
  assign new_n19155_ = ~new_n18858_ & new_n19154_;
  assign new_n19156_ = ~new_n18862_ & ~new_n19155_;
  assign new_n19157_ = ~new_n19153_ & new_n19156_;
  assign new_n19158_ = ~new_n18862_ & ~new_n19157_;
  assign new_n19159_ = \b[23]  & ~new_n18851_;
  assign new_n19160_ = ~new_n18849_ & new_n19159_;
  assign new_n19161_ = ~new_n18853_ & ~new_n19160_;
  assign new_n19162_ = ~new_n19158_ & new_n19161_;
  assign new_n19163_ = ~new_n18853_ & ~new_n19162_;
  assign new_n19164_ = \b[24]  & ~new_n18842_;
  assign new_n19165_ = ~new_n18840_ & new_n19164_;
  assign new_n19166_ = ~new_n18844_ & ~new_n19165_;
  assign new_n19167_ = ~new_n19163_ & new_n19166_;
  assign new_n19168_ = ~new_n18844_ & ~new_n19167_;
  assign new_n19169_ = \b[25]  & ~new_n18833_;
  assign new_n19170_ = ~new_n18831_ & new_n19169_;
  assign new_n19171_ = ~new_n18835_ & ~new_n19170_;
  assign new_n19172_ = ~new_n19168_ & new_n19171_;
  assign new_n19173_ = ~new_n18835_ & ~new_n19172_;
  assign new_n19174_ = \b[26]  & ~new_n18824_;
  assign new_n19175_ = ~new_n18822_ & new_n19174_;
  assign new_n19176_ = ~new_n18826_ & ~new_n19175_;
  assign new_n19177_ = ~new_n19173_ & new_n19176_;
  assign new_n19178_ = ~new_n18826_ & ~new_n19177_;
  assign new_n19179_ = \b[27]  & ~new_n18815_;
  assign new_n19180_ = ~new_n18813_ & new_n19179_;
  assign new_n19181_ = ~new_n18817_ & ~new_n19180_;
  assign new_n19182_ = ~new_n19178_ & new_n19181_;
  assign new_n19183_ = ~new_n18817_ & ~new_n19182_;
  assign new_n19184_ = \b[28]  & ~new_n18806_;
  assign new_n19185_ = ~new_n18804_ & new_n19184_;
  assign new_n19186_ = ~new_n18808_ & ~new_n19185_;
  assign new_n19187_ = ~new_n19183_ & new_n19186_;
  assign new_n19188_ = ~new_n18808_ & ~new_n19187_;
  assign new_n19189_ = \b[29]  & ~new_n18797_;
  assign new_n19190_ = ~new_n18795_ & new_n19189_;
  assign new_n19191_ = ~new_n18799_ & ~new_n19190_;
  assign new_n19192_ = ~new_n19188_ & new_n19191_;
  assign new_n19193_ = ~new_n18799_ & ~new_n19192_;
  assign new_n19194_ = \b[30]  & ~new_n18788_;
  assign new_n19195_ = ~new_n18786_ & new_n19194_;
  assign new_n19196_ = ~new_n18790_ & ~new_n19195_;
  assign new_n19197_ = ~new_n19193_ & new_n19196_;
  assign new_n19198_ = ~new_n18790_ & ~new_n19197_;
  assign new_n19199_ = \b[31]  & ~new_n18779_;
  assign new_n19200_ = ~new_n18777_ & new_n19199_;
  assign new_n19201_ = ~new_n18781_ & ~new_n19200_;
  assign new_n19202_ = ~new_n19198_ & new_n19201_;
  assign new_n19203_ = ~new_n18781_ & ~new_n19202_;
  assign new_n19204_ = \b[32]  & ~new_n18770_;
  assign new_n19205_ = ~new_n18768_ & new_n19204_;
  assign new_n19206_ = ~new_n18772_ & ~new_n19205_;
  assign new_n19207_ = ~new_n19203_ & new_n19206_;
  assign new_n19208_ = ~new_n18772_ & ~new_n19207_;
  assign new_n19209_ = \b[33]  & ~new_n18761_;
  assign new_n19210_ = ~new_n18759_ & new_n19209_;
  assign new_n19211_ = ~new_n18763_ & ~new_n19210_;
  assign new_n19212_ = ~new_n19208_ & new_n19211_;
  assign new_n19213_ = ~new_n18763_ & ~new_n19212_;
  assign new_n19214_ = \b[34]  & ~new_n18752_;
  assign new_n19215_ = ~new_n18750_ & new_n19214_;
  assign new_n19216_ = ~new_n18754_ & ~new_n19215_;
  assign new_n19217_ = ~new_n19213_ & new_n19216_;
  assign new_n19218_ = ~new_n18754_ & ~new_n19217_;
  assign new_n19219_ = \b[35]  & ~new_n18743_;
  assign new_n19220_ = ~new_n18741_ & new_n19219_;
  assign new_n19221_ = ~new_n18745_ & ~new_n19220_;
  assign new_n19222_ = ~new_n19218_ & new_n19221_;
  assign new_n19223_ = ~new_n18745_ & ~new_n19222_;
  assign new_n19224_ = \b[36]  & ~new_n18734_;
  assign new_n19225_ = ~new_n18732_ & new_n19224_;
  assign new_n19226_ = ~new_n18736_ & ~new_n19225_;
  assign new_n19227_ = ~new_n19223_ & new_n19226_;
  assign new_n19228_ = ~new_n18736_ & ~new_n19227_;
  assign new_n19229_ = \b[37]  & ~new_n18725_;
  assign new_n19230_ = ~new_n18723_ & new_n19229_;
  assign new_n19231_ = ~new_n18727_ & ~new_n19230_;
  assign new_n19232_ = ~new_n19228_ & new_n19231_;
  assign new_n19233_ = ~new_n18727_ & ~new_n19232_;
  assign new_n19234_ = \b[38]  & ~new_n18716_;
  assign new_n19235_ = ~new_n18714_ & new_n19234_;
  assign new_n19236_ = ~new_n18718_ & ~new_n19235_;
  assign new_n19237_ = ~new_n19233_ & new_n19236_;
  assign new_n19238_ = ~new_n18718_ & ~new_n19237_;
  assign new_n19239_ = \b[39]  & ~new_n18707_;
  assign new_n19240_ = ~new_n18705_ & new_n19239_;
  assign new_n19241_ = ~new_n18709_ & ~new_n19240_;
  assign new_n19242_ = ~new_n19238_ & new_n19241_;
  assign new_n19243_ = ~new_n18709_ & ~new_n19242_;
  assign new_n19244_ = \b[40]  & ~new_n18698_;
  assign new_n19245_ = ~new_n18696_ & new_n19244_;
  assign new_n19246_ = ~new_n18700_ & ~new_n19245_;
  assign new_n19247_ = ~new_n19243_ & new_n19246_;
  assign new_n19248_ = ~new_n18700_ & ~new_n19247_;
  assign new_n19249_ = \b[41]  & ~new_n18689_;
  assign new_n19250_ = ~new_n18687_ & new_n19249_;
  assign new_n19251_ = ~new_n18691_ & ~new_n19250_;
  assign new_n19252_ = ~new_n19248_ & new_n19251_;
  assign new_n19253_ = ~new_n18691_ & ~new_n19252_;
  assign new_n19254_ = \b[42]  & ~new_n18680_;
  assign new_n19255_ = ~new_n18678_ & new_n19254_;
  assign new_n19256_ = ~new_n18682_ & ~new_n19255_;
  assign new_n19257_ = ~new_n19253_ & new_n19256_;
  assign new_n19258_ = ~new_n18682_ & ~new_n19257_;
  assign new_n19259_ = \b[43]  & ~new_n18671_;
  assign new_n19260_ = ~new_n18669_ & new_n19259_;
  assign new_n19261_ = ~new_n18673_ & ~new_n19260_;
  assign new_n19262_ = ~new_n19258_ & new_n19261_;
  assign new_n19263_ = ~new_n18673_ & ~new_n19262_;
  assign new_n19264_ = \b[44]  & ~new_n18662_;
  assign new_n19265_ = ~new_n18660_ & new_n19264_;
  assign new_n19266_ = ~new_n18664_ & ~new_n19265_;
  assign new_n19267_ = ~new_n19263_ & new_n19266_;
  assign new_n19268_ = ~new_n18664_ & ~new_n19267_;
  assign new_n19269_ = \b[45]  & ~new_n18653_;
  assign new_n19270_ = ~new_n18651_ & new_n19269_;
  assign new_n19271_ = ~new_n18655_ & ~new_n19270_;
  assign new_n19272_ = ~new_n19268_ & new_n19271_;
  assign new_n19273_ = ~new_n18655_ & ~new_n19272_;
  assign new_n19274_ = \b[46]  & ~new_n18644_;
  assign new_n19275_ = ~new_n18642_ & new_n19274_;
  assign new_n19276_ = ~new_n18646_ & ~new_n19275_;
  assign new_n19277_ = ~new_n19273_ & new_n19276_;
  assign new_n19278_ = ~new_n18646_ & ~new_n19277_;
  assign new_n19279_ = \b[47]  & ~new_n18635_;
  assign new_n19280_ = ~new_n18633_ & new_n19279_;
  assign new_n19281_ = ~new_n18637_ & ~new_n19280_;
  assign new_n19282_ = ~new_n19278_ & new_n19281_;
  assign new_n19283_ = ~new_n18637_ & ~new_n19282_;
  assign new_n19284_ = \b[48]  & ~new_n18626_;
  assign new_n19285_ = ~new_n18624_ & new_n19284_;
  assign new_n19286_ = ~new_n18628_ & ~new_n19285_;
  assign new_n19287_ = ~new_n19283_ & new_n19286_;
  assign new_n19288_ = ~new_n18628_ & ~new_n19287_;
  assign new_n19289_ = \b[49]  & ~new_n18617_;
  assign new_n19290_ = ~new_n18615_ & new_n19289_;
  assign new_n19291_ = ~new_n18619_ & ~new_n19290_;
  assign new_n19292_ = ~new_n19288_ & new_n19291_;
  assign new_n19293_ = ~new_n18619_ & ~new_n19292_;
  assign new_n19294_ = \b[50]  & ~new_n18597_;
  assign new_n19295_ = ~new_n18595_ & new_n19294_;
  assign new_n19296_ = ~new_n18610_ & ~new_n19295_;
  assign new_n19297_ = ~new_n19293_ & new_n19296_;
  assign new_n19298_ = ~new_n18610_ & ~new_n19297_;
  assign new_n19299_ = \b[51]  & ~new_n18607_;
  assign new_n19300_ = ~new_n18605_ & new_n19299_;
  assign new_n19301_ = ~new_n18609_ & ~new_n19300_;
  assign new_n19302_ = ~new_n19298_ & new_n19301_;
  assign new_n19303_ = ~new_n18609_ & ~new_n19302_;
  assign \quotient[12]  = new_n288_ & ~new_n19303_;
  assign new_n19305_ = ~new_n18598_ & ~\quotient[12] ;
  assign new_n19306_ = ~new_n18619_ & new_n19296_;
  assign new_n19307_ = ~new_n19292_ & new_n19306_;
  assign new_n19308_ = ~new_n19293_ & ~new_n19296_;
  assign new_n19309_ = ~new_n19307_ & ~new_n19308_;
  assign new_n19310_ = new_n288_ & ~new_n19309_;
  assign new_n19311_ = ~new_n19303_ & new_n19310_;
  assign new_n19312_ = ~new_n19305_ & ~new_n19311_;
  assign new_n19313_ = ~\b[51]  & ~new_n19312_;
  assign new_n19314_ = ~new_n18618_ & ~\quotient[12] ;
  assign new_n19315_ = ~new_n18628_ & new_n19291_;
  assign new_n19316_ = ~new_n19287_ & new_n19315_;
  assign new_n19317_ = ~new_n19288_ & ~new_n19291_;
  assign new_n19318_ = ~new_n19316_ & ~new_n19317_;
  assign new_n19319_ = new_n288_ & ~new_n19318_;
  assign new_n19320_ = ~new_n19303_ & new_n19319_;
  assign new_n19321_ = ~new_n19314_ & ~new_n19320_;
  assign new_n19322_ = ~\b[50]  & ~new_n19321_;
  assign new_n19323_ = ~new_n18627_ & ~\quotient[12] ;
  assign new_n19324_ = ~new_n18637_ & new_n19286_;
  assign new_n19325_ = ~new_n19282_ & new_n19324_;
  assign new_n19326_ = ~new_n19283_ & ~new_n19286_;
  assign new_n19327_ = ~new_n19325_ & ~new_n19326_;
  assign new_n19328_ = new_n288_ & ~new_n19327_;
  assign new_n19329_ = ~new_n19303_ & new_n19328_;
  assign new_n19330_ = ~new_n19323_ & ~new_n19329_;
  assign new_n19331_ = ~\b[49]  & ~new_n19330_;
  assign new_n19332_ = ~new_n18636_ & ~\quotient[12] ;
  assign new_n19333_ = ~new_n18646_ & new_n19281_;
  assign new_n19334_ = ~new_n19277_ & new_n19333_;
  assign new_n19335_ = ~new_n19278_ & ~new_n19281_;
  assign new_n19336_ = ~new_n19334_ & ~new_n19335_;
  assign new_n19337_ = new_n288_ & ~new_n19336_;
  assign new_n19338_ = ~new_n19303_ & new_n19337_;
  assign new_n19339_ = ~new_n19332_ & ~new_n19338_;
  assign new_n19340_ = ~\b[48]  & ~new_n19339_;
  assign new_n19341_ = ~new_n18645_ & ~\quotient[12] ;
  assign new_n19342_ = ~new_n18655_ & new_n19276_;
  assign new_n19343_ = ~new_n19272_ & new_n19342_;
  assign new_n19344_ = ~new_n19273_ & ~new_n19276_;
  assign new_n19345_ = ~new_n19343_ & ~new_n19344_;
  assign new_n19346_ = new_n288_ & ~new_n19345_;
  assign new_n19347_ = ~new_n19303_ & new_n19346_;
  assign new_n19348_ = ~new_n19341_ & ~new_n19347_;
  assign new_n19349_ = ~\b[47]  & ~new_n19348_;
  assign new_n19350_ = ~new_n18654_ & ~\quotient[12] ;
  assign new_n19351_ = ~new_n18664_ & new_n19271_;
  assign new_n19352_ = ~new_n19267_ & new_n19351_;
  assign new_n19353_ = ~new_n19268_ & ~new_n19271_;
  assign new_n19354_ = ~new_n19352_ & ~new_n19353_;
  assign new_n19355_ = new_n288_ & ~new_n19354_;
  assign new_n19356_ = ~new_n19303_ & new_n19355_;
  assign new_n19357_ = ~new_n19350_ & ~new_n19356_;
  assign new_n19358_ = ~\b[46]  & ~new_n19357_;
  assign new_n19359_ = ~new_n18663_ & ~\quotient[12] ;
  assign new_n19360_ = ~new_n18673_ & new_n19266_;
  assign new_n19361_ = ~new_n19262_ & new_n19360_;
  assign new_n19362_ = ~new_n19263_ & ~new_n19266_;
  assign new_n19363_ = ~new_n19361_ & ~new_n19362_;
  assign new_n19364_ = new_n288_ & ~new_n19363_;
  assign new_n19365_ = ~new_n19303_ & new_n19364_;
  assign new_n19366_ = ~new_n19359_ & ~new_n19365_;
  assign new_n19367_ = ~\b[45]  & ~new_n19366_;
  assign new_n19368_ = ~new_n18672_ & ~\quotient[12] ;
  assign new_n19369_ = ~new_n18682_ & new_n19261_;
  assign new_n19370_ = ~new_n19257_ & new_n19369_;
  assign new_n19371_ = ~new_n19258_ & ~new_n19261_;
  assign new_n19372_ = ~new_n19370_ & ~new_n19371_;
  assign new_n19373_ = new_n288_ & ~new_n19372_;
  assign new_n19374_ = ~new_n19303_ & new_n19373_;
  assign new_n19375_ = ~new_n19368_ & ~new_n19374_;
  assign new_n19376_ = ~\b[44]  & ~new_n19375_;
  assign new_n19377_ = ~new_n18681_ & ~\quotient[12] ;
  assign new_n19378_ = ~new_n18691_ & new_n19256_;
  assign new_n19379_ = ~new_n19252_ & new_n19378_;
  assign new_n19380_ = ~new_n19253_ & ~new_n19256_;
  assign new_n19381_ = ~new_n19379_ & ~new_n19380_;
  assign new_n19382_ = new_n288_ & ~new_n19381_;
  assign new_n19383_ = ~new_n19303_ & new_n19382_;
  assign new_n19384_ = ~new_n19377_ & ~new_n19383_;
  assign new_n19385_ = ~\b[43]  & ~new_n19384_;
  assign new_n19386_ = ~new_n18690_ & ~\quotient[12] ;
  assign new_n19387_ = ~new_n18700_ & new_n19251_;
  assign new_n19388_ = ~new_n19247_ & new_n19387_;
  assign new_n19389_ = ~new_n19248_ & ~new_n19251_;
  assign new_n19390_ = ~new_n19388_ & ~new_n19389_;
  assign new_n19391_ = new_n288_ & ~new_n19390_;
  assign new_n19392_ = ~new_n19303_ & new_n19391_;
  assign new_n19393_ = ~new_n19386_ & ~new_n19392_;
  assign new_n19394_ = ~\b[42]  & ~new_n19393_;
  assign new_n19395_ = ~new_n18699_ & ~\quotient[12] ;
  assign new_n19396_ = ~new_n18709_ & new_n19246_;
  assign new_n19397_ = ~new_n19242_ & new_n19396_;
  assign new_n19398_ = ~new_n19243_ & ~new_n19246_;
  assign new_n19399_ = ~new_n19397_ & ~new_n19398_;
  assign new_n19400_ = new_n288_ & ~new_n19399_;
  assign new_n19401_ = ~new_n19303_ & new_n19400_;
  assign new_n19402_ = ~new_n19395_ & ~new_n19401_;
  assign new_n19403_ = ~\b[41]  & ~new_n19402_;
  assign new_n19404_ = ~new_n18708_ & ~\quotient[12] ;
  assign new_n19405_ = ~new_n18718_ & new_n19241_;
  assign new_n19406_ = ~new_n19237_ & new_n19405_;
  assign new_n19407_ = ~new_n19238_ & ~new_n19241_;
  assign new_n19408_ = ~new_n19406_ & ~new_n19407_;
  assign new_n19409_ = new_n288_ & ~new_n19408_;
  assign new_n19410_ = ~new_n19303_ & new_n19409_;
  assign new_n19411_ = ~new_n19404_ & ~new_n19410_;
  assign new_n19412_ = ~\b[40]  & ~new_n19411_;
  assign new_n19413_ = ~new_n18717_ & ~\quotient[12] ;
  assign new_n19414_ = ~new_n18727_ & new_n19236_;
  assign new_n19415_ = ~new_n19232_ & new_n19414_;
  assign new_n19416_ = ~new_n19233_ & ~new_n19236_;
  assign new_n19417_ = ~new_n19415_ & ~new_n19416_;
  assign new_n19418_ = new_n288_ & ~new_n19417_;
  assign new_n19419_ = ~new_n19303_ & new_n19418_;
  assign new_n19420_ = ~new_n19413_ & ~new_n19419_;
  assign new_n19421_ = ~\b[39]  & ~new_n19420_;
  assign new_n19422_ = ~new_n18726_ & ~\quotient[12] ;
  assign new_n19423_ = ~new_n18736_ & new_n19231_;
  assign new_n19424_ = ~new_n19227_ & new_n19423_;
  assign new_n19425_ = ~new_n19228_ & ~new_n19231_;
  assign new_n19426_ = ~new_n19424_ & ~new_n19425_;
  assign new_n19427_ = new_n288_ & ~new_n19426_;
  assign new_n19428_ = ~new_n19303_ & new_n19427_;
  assign new_n19429_ = ~new_n19422_ & ~new_n19428_;
  assign new_n19430_ = ~\b[38]  & ~new_n19429_;
  assign new_n19431_ = ~new_n18735_ & ~\quotient[12] ;
  assign new_n19432_ = ~new_n18745_ & new_n19226_;
  assign new_n19433_ = ~new_n19222_ & new_n19432_;
  assign new_n19434_ = ~new_n19223_ & ~new_n19226_;
  assign new_n19435_ = ~new_n19433_ & ~new_n19434_;
  assign new_n19436_ = new_n288_ & ~new_n19435_;
  assign new_n19437_ = ~new_n19303_ & new_n19436_;
  assign new_n19438_ = ~new_n19431_ & ~new_n19437_;
  assign new_n19439_ = ~\b[37]  & ~new_n19438_;
  assign new_n19440_ = ~new_n18744_ & ~\quotient[12] ;
  assign new_n19441_ = ~new_n18754_ & new_n19221_;
  assign new_n19442_ = ~new_n19217_ & new_n19441_;
  assign new_n19443_ = ~new_n19218_ & ~new_n19221_;
  assign new_n19444_ = ~new_n19442_ & ~new_n19443_;
  assign new_n19445_ = new_n288_ & ~new_n19444_;
  assign new_n19446_ = ~new_n19303_ & new_n19445_;
  assign new_n19447_ = ~new_n19440_ & ~new_n19446_;
  assign new_n19448_ = ~\b[36]  & ~new_n19447_;
  assign new_n19449_ = ~new_n18753_ & ~\quotient[12] ;
  assign new_n19450_ = ~new_n18763_ & new_n19216_;
  assign new_n19451_ = ~new_n19212_ & new_n19450_;
  assign new_n19452_ = ~new_n19213_ & ~new_n19216_;
  assign new_n19453_ = ~new_n19451_ & ~new_n19452_;
  assign new_n19454_ = new_n288_ & ~new_n19453_;
  assign new_n19455_ = ~new_n19303_ & new_n19454_;
  assign new_n19456_ = ~new_n19449_ & ~new_n19455_;
  assign new_n19457_ = ~\b[35]  & ~new_n19456_;
  assign new_n19458_ = ~new_n18762_ & ~\quotient[12] ;
  assign new_n19459_ = ~new_n18772_ & new_n19211_;
  assign new_n19460_ = ~new_n19207_ & new_n19459_;
  assign new_n19461_ = ~new_n19208_ & ~new_n19211_;
  assign new_n19462_ = ~new_n19460_ & ~new_n19461_;
  assign new_n19463_ = new_n288_ & ~new_n19462_;
  assign new_n19464_ = ~new_n19303_ & new_n19463_;
  assign new_n19465_ = ~new_n19458_ & ~new_n19464_;
  assign new_n19466_ = ~\b[34]  & ~new_n19465_;
  assign new_n19467_ = ~new_n18771_ & ~\quotient[12] ;
  assign new_n19468_ = ~new_n18781_ & new_n19206_;
  assign new_n19469_ = ~new_n19202_ & new_n19468_;
  assign new_n19470_ = ~new_n19203_ & ~new_n19206_;
  assign new_n19471_ = ~new_n19469_ & ~new_n19470_;
  assign new_n19472_ = new_n288_ & ~new_n19471_;
  assign new_n19473_ = ~new_n19303_ & new_n19472_;
  assign new_n19474_ = ~new_n19467_ & ~new_n19473_;
  assign new_n19475_ = ~\b[33]  & ~new_n19474_;
  assign new_n19476_ = ~new_n18780_ & ~\quotient[12] ;
  assign new_n19477_ = ~new_n18790_ & new_n19201_;
  assign new_n19478_ = ~new_n19197_ & new_n19477_;
  assign new_n19479_ = ~new_n19198_ & ~new_n19201_;
  assign new_n19480_ = ~new_n19478_ & ~new_n19479_;
  assign new_n19481_ = new_n288_ & ~new_n19480_;
  assign new_n19482_ = ~new_n19303_ & new_n19481_;
  assign new_n19483_ = ~new_n19476_ & ~new_n19482_;
  assign new_n19484_ = ~\b[32]  & ~new_n19483_;
  assign new_n19485_ = ~new_n18789_ & ~\quotient[12] ;
  assign new_n19486_ = ~new_n18799_ & new_n19196_;
  assign new_n19487_ = ~new_n19192_ & new_n19486_;
  assign new_n19488_ = ~new_n19193_ & ~new_n19196_;
  assign new_n19489_ = ~new_n19487_ & ~new_n19488_;
  assign new_n19490_ = new_n288_ & ~new_n19489_;
  assign new_n19491_ = ~new_n19303_ & new_n19490_;
  assign new_n19492_ = ~new_n19485_ & ~new_n19491_;
  assign new_n19493_ = ~\b[31]  & ~new_n19492_;
  assign new_n19494_ = ~new_n18798_ & ~\quotient[12] ;
  assign new_n19495_ = ~new_n18808_ & new_n19191_;
  assign new_n19496_ = ~new_n19187_ & new_n19495_;
  assign new_n19497_ = ~new_n19188_ & ~new_n19191_;
  assign new_n19498_ = ~new_n19496_ & ~new_n19497_;
  assign new_n19499_ = new_n288_ & ~new_n19498_;
  assign new_n19500_ = ~new_n19303_ & new_n19499_;
  assign new_n19501_ = ~new_n19494_ & ~new_n19500_;
  assign new_n19502_ = ~\b[30]  & ~new_n19501_;
  assign new_n19503_ = ~new_n18807_ & ~\quotient[12] ;
  assign new_n19504_ = ~new_n18817_ & new_n19186_;
  assign new_n19505_ = ~new_n19182_ & new_n19504_;
  assign new_n19506_ = ~new_n19183_ & ~new_n19186_;
  assign new_n19507_ = ~new_n19505_ & ~new_n19506_;
  assign new_n19508_ = new_n288_ & ~new_n19507_;
  assign new_n19509_ = ~new_n19303_ & new_n19508_;
  assign new_n19510_ = ~new_n19503_ & ~new_n19509_;
  assign new_n19511_ = ~\b[29]  & ~new_n19510_;
  assign new_n19512_ = ~new_n18816_ & ~\quotient[12] ;
  assign new_n19513_ = ~new_n18826_ & new_n19181_;
  assign new_n19514_ = ~new_n19177_ & new_n19513_;
  assign new_n19515_ = ~new_n19178_ & ~new_n19181_;
  assign new_n19516_ = ~new_n19514_ & ~new_n19515_;
  assign new_n19517_ = new_n288_ & ~new_n19516_;
  assign new_n19518_ = ~new_n19303_ & new_n19517_;
  assign new_n19519_ = ~new_n19512_ & ~new_n19518_;
  assign new_n19520_ = ~\b[28]  & ~new_n19519_;
  assign new_n19521_ = ~new_n18825_ & ~\quotient[12] ;
  assign new_n19522_ = ~new_n18835_ & new_n19176_;
  assign new_n19523_ = ~new_n19172_ & new_n19522_;
  assign new_n19524_ = ~new_n19173_ & ~new_n19176_;
  assign new_n19525_ = ~new_n19523_ & ~new_n19524_;
  assign new_n19526_ = new_n288_ & ~new_n19525_;
  assign new_n19527_ = ~new_n19303_ & new_n19526_;
  assign new_n19528_ = ~new_n19521_ & ~new_n19527_;
  assign new_n19529_ = ~\b[27]  & ~new_n19528_;
  assign new_n19530_ = ~new_n18834_ & ~\quotient[12] ;
  assign new_n19531_ = ~new_n18844_ & new_n19171_;
  assign new_n19532_ = ~new_n19167_ & new_n19531_;
  assign new_n19533_ = ~new_n19168_ & ~new_n19171_;
  assign new_n19534_ = ~new_n19532_ & ~new_n19533_;
  assign new_n19535_ = new_n288_ & ~new_n19534_;
  assign new_n19536_ = ~new_n19303_ & new_n19535_;
  assign new_n19537_ = ~new_n19530_ & ~new_n19536_;
  assign new_n19538_ = ~\b[26]  & ~new_n19537_;
  assign new_n19539_ = ~new_n18843_ & ~\quotient[12] ;
  assign new_n19540_ = ~new_n18853_ & new_n19166_;
  assign new_n19541_ = ~new_n19162_ & new_n19540_;
  assign new_n19542_ = ~new_n19163_ & ~new_n19166_;
  assign new_n19543_ = ~new_n19541_ & ~new_n19542_;
  assign new_n19544_ = new_n288_ & ~new_n19543_;
  assign new_n19545_ = ~new_n19303_ & new_n19544_;
  assign new_n19546_ = ~new_n19539_ & ~new_n19545_;
  assign new_n19547_ = ~\b[25]  & ~new_n19546_;
  assign new_n19548_ = ~new_n18852_ & ~\quotient[12] ;
  assign new_n19549_ = ~new_n18862_ & new_n19161_;
  assign new_n19550_ = ~new_n19157_ & new_n19549_;
  assign new_n19551_ = ~new_n19158_ & ~new_n19161_;
  assign new_n19552_ = ~new_n19550_ & ~new_n19551_;
  assign new_n19553_ = new_n288_ & ~new_n19552_;
  assign new_n19554_ = ~new_n19303_ & new_n19553_;
  assign new_n19555_ = ~new_n19548_ & ~new_n19554_;
  assign new_n19556_ = ~\b[24]  & ~new_n19555_;
  assign new_n19557_ = ~new_n18861_ & ~\quotient[12] ;
  assign new_n19558_ = ~new_n18871_ & new_n19156_;
  assign new_n19559_ = ~new_n19152_ & new_n19558_;
  assign new_n19560_ = ~new_n19153_ & ~new_n19156_;
  assign new_n19561_ = ~new_n19559_ & ~new_n19560_;
  assign new_n19562_ = new_n288_ & ~new_n19561_;
  assign new_n19563_ = ~new_n19303_ & new_n19562_;
  assign new_n19564_ = ~new_n19557_ & ~new_n19563_;
  assign new_n19565_ = ~\b[23]  & ~new_n19564_;
  assign new_n19566_ = ~new_n18870_ & ~\quotient[12] ;
  assign new_n19567_ = ~new_n18880_ & new_n19151_;
  assign new_n19568_ = ~new_n19147_ & new_n19567_;
  assign new_n19569_ = ~new_n19148_ & ~new_n19151_;
  assign new_n19570_ = ~new_n19568_ & ~new_n19569_;
  assign new_n19571_ = new_n288_ & ~new_n19570_;
  assign new_n19572_ = ~new_n19303_ & new_n19571_;
  assign new_n19573_ = ~new_n19566_ & ~new_n19572_;
  assign new_n19574_ = ~\b[22]  & ~new_n19573_;
  assign new_n19575_ = ~new_n18879_ & ~\quotient[12] ;
  assign new_n19576_ = ~new_n18889_ & new_n19146_;
  assign new_n19577_ = ~new_n19142_ & new_n19576_;
  assign new_n19578_ = ~new_n19143_ & ~new_n19146_;
  assign new_n19579_ = ~new_n19577_ & ~new_n19578_;
  assign new_n19580_ = new_n288_ & ~new_n19579_;
  assign new_n19581_ = ~new_n19303_ & new_n19580_;
  assign new_n19582_ = ~new_n19575_ & ~new_n19581_;
  assign new_n19583_ = ~\b[21]  & ~new_n19582_;
  assign new_n19584_ = ~new_n18888_ & ~\quotient[12] ;
  assign new_n19585_ = ~new_n18898_ & new_n19141_;
  assign new_n19586_ = ~new_n19137_ & new_n19585_;
  assign new_n19587_ = ~new_n19138_ & ~new_n19141_;
  assign new_n19588_ = ~new_n19586_ & ~new_n19587_;
  assign new_n19589_ = new_n288_ & ~new_n19588_;
  assign new_n19590_ = ~new_n19303_ & new_n19589_;
  assign new_n19591_ = ~new_n19584_ & ~new_n19590_;
  assign new_n19592_ = ~\b[20]  & ~new_n19591_;
  assign new_n19593_ = ~new_n18897_ & ~\quotient[12] ;
  assign new_n19594_ = ~new_n18907_ & new_n19136_;
  assign new_n19595_ = ~new_n19132_ & new_n19594_;
  assign new_n19596_ = ~new_n19133_ & ~new_n19136_;
  assign new_n19597_ = ~new_n19595_ & ~new_n19596_;
  assign new_n19598_ = new_n288_ & ~new_n19597_;
  assign new_n19599_ = ~new_n19303_ & new_n19598_;
  assign new_n19600_ = ~new_n19593_ & ~new_n19599_;
  assign new_n19601_ = ~\b[19]  & ~new_n19600_;
  assign new_n19602_ = ~new_n18906_ & ~\quotient[12] ;
  assign new_n19603_ = ~new_n18916_ & new_n19131_;
  assign new_n19604_ = ~new_n19127_ & new_n19603_;
  assign new_n19605_ = ~new_n19128_ & ~new_n19131_;
  assign new_n19606_ = ~new_n19604_ & ~new_n19605_;
  assign new_n19607_ = new_n288_ & ~new_n19606_;
  assign new_n19608_ = ~new_n19303_ & new_n19607_;
  assign new_n19609_ = ~new_n19602_ & ~new_n19608_;
  assign new_n19610_ = ~\b[18]  & ~new_n19609_;
  assign new_n19611_ = ~new_n18915_ & ~\quotient[12] ;
  assign new_n19612_ = ~new_n18925_ & new_n19126_;
  assign new_n19613_ = ~new_n19122_ & new_n19612_;
  assign new_n19614_ = ~new_n19123_ & ~new_n19126_;
  assign new_n19615_ = ~new_n19613_ & ~new_n19614_;
  assign new_n19616_ = new_n288_ & ~new_n19615_;
  assign new_n19617_ = ~new_n19303_ & new_n19616_;
  assign new_n19618_ = ~new_n19611_ & ~new_n19617_;
  assign new_n19619_ = ~\b[17]  & ~new_n19618_;
  assign new_n19620_ = ~new_n18924_ & ~\quotient[12] ;
  assign new_n19621_ = ~new_n18934_ & new_n19121_;
  assign new_n19622_ = ~new_n19117_ & new_n19621_;
  assign new_n19623_ = ~new_n19118_ & ~new_n19121_;
  assign new_n19624_ = ~new_n19622_ & ~new_n19623_;
  assign new_n19625_ = new_n288_ & ~new_n19624_;
  assign new_n19626_ = ~new_n19303_ & new_n19625_;
  assign new_n19627_ = ~new_n19620_ & ~new_n19626_;
  assign new_n19628_ = ~\b[16]  & ~new_n19627_;
  assign new_n19629_ = ~new_n18933_ & ~\quotient[12] ;
  assign new_n19630_ = ~new_n18943_ & new_n19116_;
  assign new_n19631_ = ~new_n19112_ & new_n19630_;
  assign new_n19632_ = ~new_n19113_ & ~new_n19116_;
  assign new_n19633_ = ~new_n19631_ & ~new_n19632_;
  assign new_n19634_ = new_n288_ & ~new_n19633_;
  assign new_n19635_ = ~new_n19303_ & new_n19634_;
  assign new_n19636_ = ~new_n19629_ & ~new_n19635_;
  assign new_n19637_ = ~\b[15]  & ~new_n19636_;
  assign new_n19638_ = ~new_n18942_ & ~\quotient[12] ;
  assign new_n19639_ = ~new_n18952_ & new_n19111_;
  assign new_n19640_ = ~new_n19107_ & new_n19639_;
  assign new_n19641_ = ~new_n19108_ & ~new_n19111_;
  assign new_n19642_ = ~new_n19640_ & ~new_n19641_;
  assign new_n19643_ = new_n288_ & ~new_n19642_;
  assign new_n19644_ = ~new_n19303_ & new_n19643_;
  assign new_n19645_ = ~new_n19638_ & ~new_n19644_;
  assign new_n19646_ = ~\b[14]  & ~new_n19645_;
  assign new_n19647_ = ~new_n18951_ & ~\quotient[12] ;
  assign new_n19648_ = ~new_n18961_ & new_n19106_;
  assign new_n19649_ = ~new_n19102_ & new_n19648_;
  assign new_n19650_ = ~new_n19103_ & ~new_n19106_;
  assign new_n19651_ = ~new_n19649_ & ~new_n19650_;
  assign new_n19652_ = new_n288_ & ~new_n19651_;
  assign new_n19653_ = ~new_n19303_ & new_n19652_;
  assign new_n19654_ = ~new_n19647_ & ~new_n19653_;
  assign new_n19655_ = ~\b[13]  & ~new_n19654_;
  assign new_n19656_ = ~new_n18960_ & ~\quotient[12] ;
  assign new_n19657_ = ~new_n18970_ & new_n19101_;
  assign new_n19658_ = ~new_n19097_ & new_n19657_;
  assign new_n19659_ = ~new_n19098_ & ~new_n19101_;
  assign new_n19660_ = ~new_n19658_ & ~new_n19659_;
  assign new_n19661_ = new_n288_ & ~new_n19660_;
  assign new_n19662_ = ~new_n19303_ & new_n19661_;
  assign new_n19663_ = ~new_n19656_ & ~new_n19662_;
  assign new_n19664_ = ~\b[12]  & ~new_n19663_;
  assign new_n19665_ = ~new_n18969_ & ~\quotient[12] ;
  assign new_n19666_ = ~new_n18979_ & new_n19096_;
  assign new_n19667_ = ~new_n19092_ & new_n19666_;
  assign new_n19668_ = ~new_n19093_ & ~new_n19096_;
  assign new_n19669_ = ~new_n19667_ & ~new_n19668_;
  assign new_n19670_ = new_n288_ & ~new_n19669_;
  assign new_n19671_ = ~new_n19303_ & new_n19670_;
  assign new_n19672_ = ~new_n19665_ & ~new_n19671_;
  assign new_n19673_ = ~\b[11]  & ~new_n19672_;
  assign new_n19674_ = ~new_n18978_ & ~\quotient[12] ;
  assign new_n19675_ = ~new_n18988_ & new_n19091_;
  assign new_n19676_ = ~new_n19087_ & new_n19675_;
  assign new_n19677_ = ~new_n19088_ & ~new_n19091_;
  assign new_n19678_ = ~new_n19676_ & ~new_n19677_;
  assign new_n19679_ = new_n288_ & ~new_n19678_;
  assign new_n19680_ = ~new_n19303_ & new_n19679_;
  assign new_n19681_ = ~new_n19674_ & ~new_n19680_;
  assign new_n19682_ = ~\b[10]  & ~new_n19681_;
  assign new_n19683_ = ~new_n18987_ & ~\quotient[12] ;
  assign new_n19684_ = ~new_n18997_ & new_n19086_;
  assign new_n19685_ = ~new_n19082_ & new_n19684_;
  assign new_n19686_ = ~new_n19083_ & ~new_n19086_;
  assign new_n19687_ = ~new_n19685_ & ~new_n19686_;
  assign new_n19688_ = new_n288_ & ~new_n19687_;
  assign new_n19689_ = ~new_n19303_ & new_n19688_;
  assign new_n19690_ = ~new_n19683_ & ~new_n19689_;
  assign new_n19691_ = ~\b[9]  & ~new_n19690_;
  assign new_n19692_ = ~new_n18996_ & ~\quotient[12] ;
  assign new_n19693_ = ~new_n19006_ & new_n19081_;
  assign new_n19694_ = ~new_n19077_ & new_n19693_;
  assign new_n19695_ = ~new_n19078_ & ~new_n19081_;
  assign new_n19696_ = ~new_n19694_ & ~new_n19695_;
  assign new_n19697_ = new_n288_ & ~new_n19696_;
  assign new_n19698_ = ~new_n19303_ & new_n19697_;
  assign new_n19699_ = ~new_n19692_ & ~new_n19698_;
  assign new_n19700_ = ~\b[8]  & ~new_n19699_;
  assign new_n19701_ = ~new_n19005_ & ~\quotient[12] ;
  assign new_n19702_ = ~new_n19015_ & new_n19076_;
  assign new_n19703_ = ~new_n19072_ & new_n19702_;
  assign new_n19704_ = ~new_n19073_ & ~new_n19076_;
  assign new_n19705_ = ~new_n19703_ & ~new_n19704_;
  assign new_n19706_ = new_n288_ & ~new_n19705_;
  assign new_n19707_ = ~new_n19303_ & new_n19706_;
  assign new_n19708_ = ~new_n19701_ & ~new_n19707_;
  assign new_n19709_ = ~\b[7]  & ~new_n19708_;
  assign new_n19710_ = ~new_n19014_ & ~\quotient[12] ;
  assign new_n19711_ = ~new_n19024_ & new_n19071_;
  assign new_n19712_ = ~new_n19067_ & new_n19711_;
  assign new_n19713_ = ~new_n19068_ & ~new_n19071_;
  assign new_n19714_ = ~new_n19712_ & ~new_n19713_;
  assign new_n19715_ = new_n288_ & ~new_n19714_;
  assign new_n19716_ = ~new_n19303_ & new_n19715_;
  assign new_n19717_ = ~new_n19710_ & ~new_n19716_;
  assign new_n19718_ = ~\b[6]  & ~new_n19717_;
  assign new_n19719_ = ~new_n19023_ & ~\quotient[12] ;
  assign new_n19720_ = ~new_n19033_ & new_n19066_;
  assign new_n19721_ = ~new_n19062_ & new_n19720_;
  assign new_n19722_ = ~new_n19063_ & ~new_n19066_;
  assign new_n19723_ = ~new_n19721_ & ~new_n19722_;
  assign new_n19724_ = new_n288_ & ~new_n19723_;
  assign new_n19725_ = ~new_n19303_ & new_n19724_;
  assign new_n19726_ = ~new_n19719_ & ~new_n19725_;
  assign new_n19727_ = ~\b[5]  & ~new_n19726_;
  assign new_n19728_ = ~new_n19032_ & ~\quotient[12] ;
  assign new_n19729_ = ~new_n19041_ & new_n19061_;
  assign new_n19730_ = ~new_n19057_ & new_n19729_;
  assign new_n19731_ = ~new_n19058_ & ~new_n19061_;
  assign new_n19732_ = ~new_n19730_ & ~new_n19731_;
  assign new_n19733_ = new_n288_ & ~new_n19732_;
  assign new_n19734_ = ~new_n19303_ & new_n19733_;
  assign new_n19735_ = ~new_n19728_ & ~new_n19734_;
  assign new_n19736_ = ~\b[4]  & ~new_n19735_;
  assign new_n19737_ = ~new_n19040_ & ~\quotient[12] ;
  assign new_n19738_ = ~new_n19052_ & new_n19056_;
  assign new_n19739_ = ~new_n19051_ & new_n19738_;
  assign new_n19740_ = ~new_n19053_ & ~new_n19056_;
  assign new_n19741_ = ~new_n19739_ & ~new_n19740_;
  assign new_n19742_ = new_n288_ & ~new_n19741_;
  assign new_n19743_ = ~new_n19303_ & new_n19742_;
  assign new_n19744_ = ~new_n19737_ & ~new_n19743_;
  assign new_n19745_ = ~\b[3]  & ~new_n19744_;
  assign new_n19746_ = ~new_n19045_ & ~\quotient[12] ;
  assign new_n19747_ = ~new_n19048_ & new_n19050_;
  assign new_n19748_ = ~new_n19046_ & new_n19747_;
  assign new_n19749_ = new_n288_ & ~new_n19748_;
  assign new_n19750_ = ~new_n19051_ & new_n19749_;
  assign new_n19751_ = ~new_n19303_ & new_n19750_;
  assign new_n19752_ = ~new_n19746_ & ~new_n19751_;
  assign new_n19753_ = ~\b[2]  & ~new_n19752_;
  assign new_n19754_ = \b[0]  & ~\b[52] ;
  assign new_n19755_ = new_n397_ & new_n19754_;
  assign new_n19756_ = new_n407_ & new_n19755_;
  assign new_n19757_ = ~new_n19303_ & new_n19756_;
  assign new_n19758_ = \a[12]  & ~new_n19757_;
  assign new_n19759_ = new_n286_ & new_n19050_;
  assign new_n19760_ = new_n337_ & new_n19759_;
  assign new_n19761_ = ~new_n19303_ & new_n19760_;
  assign new_n19762_ = ~new_n19758_ & ~new_n19761_;
  assign new_n19763_ = \b[1]  & ~new_n19762_;
  assign new_n19764_ = ~\b[1]  & ~new_n19761_;
  assign new_n19765_ = ~new_n19758_ & new_n19764_;
  assign new_n19766_ = ~new_n19763_ & ~new_n19765_;
  assign new_n19767_ = ~\a[11]  & \b[0] ;
  assign new_n19768_ = ~new_n19766_ & ~new_n19767_;
  assign new_n19769_ = ~\b[1]  & ~new_n19762_;
  assign new_n19770_ = ~new_n19768_ & ~new_n19769_;
  assign new_n19771_ = \b[2]  & ~new_n19751_;
  assign new_n19772_ = ~new_n19746_ & new_n19771_;
  assign new_n19773_ = ~new_n19753_ & ~new_n19772_;
  assign new_n19774_ = ~new_n19770_ & new_n19773_;
  assign new_n19775_ = ~new_n19753_ & ~new_n19774_;
  assign new_n19776_ = \b[3]  & ~new_n19743_;
  assign new_n19777_ = ~new_n19737_ & new_n19776_;
  assign new_n19778_ = ~new_n19745_ & ~new_n19777_;
  assign new_n19779_ = ~new_n19775_ & new_n19778_;
  assign new_n19780_ = ~new_n19745_ & ~new_n19779_;
  assign new_n19781_ = \b[4]  & ~new_n19734_;
  assign new_n19782_ = ~new_n19728_ & new_n19781_;
  assign new_n19783_ = ~new_n19736_ & ~new_n19782_;
  assign new_n19784_ = ~new_n19780_ & new_n19783_;
  assign new_n19785_ = ~new_n19736_ & ~new_n19784_;
  assign new_n19786_ = \b[5]  & ~new_n19725_;
  assign new_n19787_ = ~new_n19719_ & new_n19786_;
  assign new_n19788_ = ~new_n19727_ & ~new_n19787_;
  assign new_n19789_ = ~new_n19785_ & new_n19788_;
  assign new_n19790_ = ~new_n19727_ & ~new_n19789_;
  assign new_n19791_ = \b[6]  & ~new_n19716_;
  assign new_n19792_ = ~new_n19710_ & new_n19791_;
  assign new_n19793_ = ~new_n19718_ & ~new_n19792_;
  assign new_n19794_ = ~new_n19790_ & new_n19793_;
  assign new_n19795_ = ~new_n19718_ & ~new_n19794_;
  assign new_n19796_ = \b[7]  & ~new_n19707_;
  assign new_n19797_ = ~new_n19701_ & new_n19796_;
  assign new_n19798_ = ~new_n19709_ & ~new_n19797_;
  assign new_n19799_ = ~new_n19795_ & new_n19798_;
  assign new_n19800_ = ~new_n19709_ & ~new_n19799_;
  assign new_n19801_ = \b[8]  & ~new_n19698_;
  assign new_n19802_ = ~new_n19692_ & new_n19801_;
  assign new_n19803_ = ~new_n19700_ & ~new_n19802_;
  assign new_n19804_ = ~new_n19800_ & new_n19803_;
  assign new_n19805_ = ~new_n19700_ & ~new_n19804_;
  assign new_n19806_ = \b[9]  & ~new_n19689_;
  assign new_n19807_ = ~new_n19683_ & new_n19806_;
  assign new_n19808_ = ~new_n19691_ & ~new_n19807_;
  assign new_n19809_ = ~new_n19805_ & new_n19808_;
  assign new_n19810_ = ~new_n19691_ & ~new_n19809_;
  assign new_n19811_ = \b[10]  & ~new_n19680_;
  assign new_n19812_ = ~new_n19674_ & new_n19811_;
  assign new_n19813_ = ~new_n19682_ & ~new_n19812_;
  assign new_n19814_ = ~new_n19810_ & new_n19813_;
  assign new_n19815_ = ~new_n19682_ & ~new_n19814_;
  assign new_n19816_ = \b[11]  & ~new_n19671_;
  assign new_n19817_ = ~new_n19665_ & new_n19816_;
  assign new_n19818_ = ~new_n19673_ & ~new_n19817_;
  assign new_n19819_ = ~new_n19815_ & new_n19818_;
  assign new_n19820_ = ~new_n19673_ & ~new_n19819_;
  assign new_n19821_ = \b[12]  & ~new_n19662_;
  assign new_n19822_ = ~new_n19656_ & new_n19821_;
  assign new_n19823_ = ~new_n19664_ & ~new_n19822_;
  assign new_n19824_ = ~new_n19820_ & new_n19823_;
  assign new_n19825_ = ~new_n19664_ & ~new_n19824_;
  assign new_n19826_ = \b[13]  & ~new_n19653_;
  assign new_n19827_ = ~new_n19647_ & new_n19826_;
  assign new_n19828_ = ~new_n19655_ & ~new_n19827_;
  assign new_n19829_ = ~new_n19825_ & new_n19828_;
  assign new_n19830_ = ~new_n19655_ & ~new_n19829_;
  assign new_n19831_ = \b[14]  & ~new_n19644_;
  assign new_n19832_ = ~new_n19638_ & new_n19831_;
  assign new_n19833_ = ~new_n19646_ & ~new_n19832_;
  assign new_n19834_ = ~new_n19830_ & new_n19833_;
  assign new_n19835_ = ~new_n19646_ & ~new_n19834_;
  assign new_n19836_ = \b[15]  & ~new_n19635_;
  assign new_n19837_ = ~new_n19629_ & new_n19836_;
  assign new_n19838_ = ~new_n19637_ & ~new_n19837_;
  assign new_n19839_ = ~new_n19835_ & new_n19838_;
  assign new_n19840_ = ~new_n19637_ & ~new_n19839_;
  assign new_n19841_ = \b[16]  & ~new_n19626_;
  assign new_n19842_ = ~new_n19620_ & new_n19841_;
  assign new_n19843_ = ~new_n19628_ & ~new_n19842_;
  assign new_n19844_ = ~new_n19840_ & new_n19843_;
  assign new_n19845_ = ~new_n19628_ & ~new_n19844_;
  assign new_n19846_ = \b[17]  & ~new_n19617_;
  assign new_n19847_ = ~new_n19611_ & new_n19846_;
  assign new_n19848_ = ~new_n19619_ & ~new_n19847_;
  assign new_n19849_ = ~new_n19845_ & new_n19848_;
  assign new_n19850_ = ~new_n19619_ & ~new_n19849_;
  assign new_n19851_ = \b[18]  & ~new_n19608_;
  assign new_n19852_ = ~new_n19602_ & new_n19851_;
  assign new_n19853_ = ~new_n19610_ & ~new_n19852_;
  assign new_n19854_ = ~new_n19850_ & new_n19853_;
  assign new_n19855_ = ~new_n19610_ & ~new_n19854_;
  assign new_n19856_ = \b[19]  & ~new_n19599_;
  assign new_n19857_ = ~new_n19593_ & new_n19856_;
  assign new_n19858_ = ~new_n19601_ & ~new_n19857_;
  assign new_n19859_ = ~new_n19855_ & new_n19858_;
  assign new_n19860_ = ~new_n19601_ & ~new_n19859_;
  assign new_n19861_ = \b[20]  & ~new_n19590_;
  assign new_n19862_ = ~new_n19584_ & new_n19861_;
  assign new_n19863_ = ~new_n19592_ & ~new_n19862_;
  assign new_n19864_ = ~new_n19860_ & new_n19863_;
  assign new_n19865_ = ~new_n19592_ & ~new_n19864_;
  assign new_n19866_ = \b[21]  & ~new_n19581_;
  assign new_n19867_ = ~new_n19575_ & new_n19866_;
  assign new_n19868_ = ~new_n19583_ & ~new_n19867_;
  assign new_n19869_ = ~new_n19865_ & new_n19868_;
  assign new_n19870_ = ~new_n19583_ & ~new_n19869_;
  assign new_n19871_ = \b[22]  & ~new_n19572_;
  assign new_n19872_ = ~new_n19566_ & new_n19871_;
  assign new_n19873_ = ~new_n19574_ & ~new_n19872_;
  assign new_n19874_ = ~new_n19870_ & new_n19873_;
  assign new_n19875_ = ~new_n19574_ & ~new_n19874_;
  assign new_n19876_ = \b[23]  & ~new_n19563_;
  assign new_n19877_ = ~new_n19557_ & new_n19876_;
  assign new_n19878_ = ~new_n19565_ & ~new_n19877_;
  assign new_n19879_ = ~new_n19875_ & new_n19878_;
  assign new_n19880_ = ~new_n19565_ & ~new_n19879_;
  assign new_n19881_ = \b[24]  & ~new_n19554_;
  assign new_n19882_ = ~new_n19548_ & new_n19881_;
  assign new_n19883_ = ~new_n19556_ & ~new_n19882_;
  assign new_n19884_ = ~new_n19880_ & new_n19883_;
  assign new_n19885_ = ~new_n19556_ & ~new_n19884_;
  assign new_n19886_ = \b[25]  & ~new_n19545_;
  assign new_n19887_ = ~new_n19539_ & new_n19886_;
  assign new_n19888_ = ~new_n19547_ & ~new_n19887_;
  assign new_n19889_ = ~new_n19885_ & new_n19888_;
  assign new_n19890_ = ~new_n19547_ & ~new_n19889_;
  assign new_n19891_ = \b[26]  & ~new_n19536_;
  assign new_n19892_ = ~new_n19530_ & new_n19891_;
  assign new_n19893_ = ~new_n19538_ & ~new_n19892_;
  assign new_n19894_ = ~new_n19890_ & new_n19893_;
  assign new_n19895_ = ~new_n19538_ & ~new_n19894_;
  assign new_n19896_ = \b[27]  & ~new_n19527_;
  assign new_n19897_ = ~new_n19521_ & new_n19896_;
  assign new_n19898_ = ~new_n19529_ & ~new_n19897_;
  assign new_n19899_ = ~new_n19895_ & new_n19898_;
  assign new_n19900_ = ~new_n19529_ & ~new_n19899_;
  assign new_n19901_ = \b[28]  & ~new_n19518_;
  assign new_n19902_ = ~new_n19512_ & new_n19901_;
  assign new_n19903_ = ~new_n19520_ & ~new_n19902_;
  assign new_n19904_ = ~new_n19900_ & new_n19903_;
  assign new_n19905_ = ~new_n19520_ & ~new_n19904_;
  assign new_n19906_ = \b[29]  & ~new_n19509_;
  assign new_n19907_ = ~new_n19503_ & new_n19906_;
  assign new_n19908_ = ~new_n19511_ & ~new_n19907_;
  assign new_n19909_ = ~new_n19905_ & new_n19908_;
  assign new_n19910_ = ~new_n19511_ & ~new_n19909_;
  assign new_n19911_ = \b[30]  & ~new_n19500_;
  assign new_n19912_ = ~new_n19494_ & new_n19911_;
  assign new_n19913_ = ~new_n19502_ & ~new_n19912_;
  assign new_n19914_ = ~new_n19910_ & new_n19913_;
  assign new_n19915_ = ~new_n19502_ & ~new_n19914_;
  assign new_n19916_ = \b[31]  & ~new_n19491_;
  assign new_n19917_ = ~new_n19485_ & new_n19916_;
  assign new_n19918_ = ~new_n19493_ & ~new_n19917_;
  assign new_n19919_ = ~new_n19915_ & new_n19918_;
  assign new_n19920_ = ~new_n19493_ & ~new_n19919_;
  assign new_n19921_ = \b[32]  & ~new_n19482_;
  assign new_n19922_ = ~new_n19476_ & new_n19921_;
  assign new_n19923_ = ~new_n19484_ & ~new_n19922_;
  assign new_n19924_ = ~new_n19920_ & new_n19923_;
  assign new_n19925_ = ~new_n19484_ & ~new_n19924_;
  assign new_n19926_ = \b[33]  & ~new_n19473_;
  assign new_n19927_ = ~new_n19467_ & new_n19926_;
  assign new_n19928_ = ~new_n19475_ & ~new_n19927_;
  assign new_n19929_ = ~new_n19925_ & new_n19928_;
  assign new_n19930_ = ~new_n19475_ & ~new_n19929_;
  assign new_n19931_ = \b[34]  & ~new_n19464_;
  assign new_n19932_ = ~new_n19458_ & new_n19931_;
  assign new_n19933_ = ~new_n19466_ & ~new_n19932_;
  assign new_n19934_ = ~new_n19930_ & new_n19933_;
  assign new_n19935_ = ~new_n19466_ & ~new_n19934_;
  assign new_n19936_ = \b[35]  & ~new_n19455_;
  assign new_n19937_ = ~new_n19449_ & new_n19936_;
  assign new_n19938_ = ~new_n19457_ & ~new_n19937_;
  assign new_n19939_ = ~new_n19935_ & new_n19938_;
  assign new_n19940_ = ~new_n19457_ & ~new_n19939_;
  assign new_n19941_ = \b[36]  & ~new_n19446_;
  assign new_n19942_ = ~new_n19440_ & new_n19941_;
  assign new_n19943_ = ~new_n19448_ & ~new_n19942_;
  assign new_n19944_ = ~new_n19940_ & new_n19943_;
  assign new_n19945_ = ~new_n19448_ & ~new_n19944_;
  assign new_n19946_ = \b[37]  & ~new_n19437_;
  assign new_n19947_ = ~new_n19431_ & new_n19946_;
  assign new_n19948_ = ~new_n19439_ & ~new_n19947_;
  assign new_n19949_ = ~new_n19945_ & new_n19948_;
  assign new_n19950_ = ~new_n19439_ & ~new_n19949_;
  assign new_n19951_ = \b[38]  & ~new_n19428_;
  assign new_n19952_ = ~new_n19422_ & new_n19951_;
  assign new_n19953_ = ~new_n19430_ & ~new_n19952_;
  assign new_n19954_ = ~new_n19950_ & new_n19953_;
  assign new_n19955_ = ~new_n19430_ & ~new_n19954_;
  assign new_n19956_ = \b[39]  & ~new_n19419_;
  assign new_n19957_ = ~new_n19413_ & new_n19956_;
  assign new_n19958_ = ~new_n19421_ & ~new_n19957_;
  assign new_n19959_ = ~new_n19955_ & new_n19958_;
  assign new_n19960_ = ~new_n19421_ & ~new_n19959_;
  assign new_n19961_ = \b[40]  & ~new_n19410_;
  assign new_n19962_ = ~new_n19404_ & new_n19961_;
  assign new_n19963_ = ~new_n19412_ & ~new_n19962_;
  assign new_n19964_ = ~new_n19960_ & new_n19963_;
  assign new_n19965_ = ~new_n19412_ & ~new_n19964_;
  assign new_n19966_ = \b[41]  & ~new_n19401_;
  assign new_n19967_ = ~new_n19395_ & new_n19966_;
  assign new_n19968_ = ~new_n19403_ & ~new_n19967_;
  assign new_n19969_ = ~new_n19965_ & new_n19968_;
  assign new_n19970_ = ~new_n19403_ & ~new_n19969_;
  assign new_n19971_ = \b[42]  & ~new_n19392_;
  assign new_n19972_ = ~new_n19386_ & new_n19971_;
  assign new_n19973_ = ~new_n19394_ & ~new_n19972_;
  assign new_n19974_ = ~new_n19970_ & new_n19973_;
  assign new_n19975_ = ~new_n19394_ & ~new_n19974_;
  assign new_n19976_ = \b[43]  & ~new_n19383_;
  assign new_n19977_ = ~new_n19377_ & new_n19976_;
  assign new_n19978_ = ~new_n19385_ & ~new_n19977_;
  assign new_n19979_ = ~new_n19975_ & new_n19978_;
  assign new_n19980_ = ~new_n19385_ & ~new_n19979_;
  assign new_n19981_ = \b[44]  & ~new_n19374_;
  assign new_n19982_ = ~new_n19368_ & new_n19981_;
  assign new_n19983_ = ~new_n19376_ & ~new_n19982_;
  assign new_n19984_ = ~new_n19980_ & new_n19983_;
  assign new_n19985_ = ~new_n19376_ & ~new_n19984_;
  assign new_n19986_ = \b[45]  & ~new_n19365_;
  assign new_n19987_ = ~new_n19359_ & new_n19986_;
  assign new_n19988_ = ~new_n19367_ & ~new_n19987_;
  assign new_n19989_ = ~new_n19985_ & new_n19988_;
  assign new_n19990_ = ~new_n19367_ & ~new_n19989_;
  assign new_n19991_ = \b[46]  & ~new_n19356_;
  assign new_n19992_ = ~new_n19350_ & new_n19991_;
  assign new_n19993_ = ~new_n19358_ & ~new_n19992_;
  assign new_n19994_ = ~new_n19990_ & new_n19993_;
  assign new_n19995_ = ~new_n19358_ & ~new_n19994_;
  assign new_n19996_ = \b[47]  & ~new_n19347_;
  assign new_n19997_ = ~new_n19341_ & new_n19996_;
  assign new_n19998_ = ~new_n19349_ & ~new_n19997_;
  assign new_n19999_ = ~new_n19995_ & new_n19998_;
  assign new_n20000_ = ~new_n19349_ & ~new_n19999_;
  assign new_n20001_ = \b[48]  & ~new_n19338_;
  assign new_n20002_ = ~new_n19332_ & new_n20001_;
  assign new_n20003_ = ~new_n19340_ & ~new_n20002_;
  assign new_n20004_ = ~new_n20000_ & new_n20003_;
  assign new_n20005_ = ~new_n19340_ & ~new_n20004_;
  assign new_n20006_ = \b[49]  & ~new_n19329_;
  assign new_n20007_ = ~new_n19323_ & new_n20006_;
  assign new_n20008_ = ~new_n19331_ & ~new_n20007_;
  assign new_n20009_ = ~new_n20005_ & new_n20008_;
  assign new_n20010_ = ~new_n19331_ & ~new_n20009_;
  assign new_n20011_ = \b[50]  & ~new_n19320_;
  assign new_n20012_ = ~new_n19314_ & new_n20011_;
  assign new_n20013_ = ~new_n19322_ & ~new_n20012_;
  assign new_n20014_ = ~new_n20010_ & new_n20013_;
  assign new_n20015_ = ~new_n19322_ & ~new_n20014_;
  assign new_n20016_ = \b[51]  & ~new_n19311_;
  assign new_n20017_ = ~new_n19305_ & new_n20016_;
  assign new_n20018_ = ~new_n19313_ & ~new_n20017_;
  assign new_n20019_ = ~new_n20015_ & new_n20018_;
  assign new_n20020_ = ~new_n19313_ & ~new_n20019_;
  assign new_n20021_ = ~new_n18608_ & ~\quotient[12] ;
  assign new_n20022_ = ~new_n18610_ & new_n19301_;
  assign new_n20023_ = ~new_n19297_ & new_n20022_;
  assign new_n20024_ = ~new_n19298_ & ~new_n19301_;
  assign new_n20025_ = ~new_n20023_ & ~new_n20024_;
  assign new_n20026_ = \quotient[12]  & ~new_n20025_;
  assign new_n20027_ = ~new_n20021_ & ~new_n20026_;
  assign new_n20028_ = ~\b[52]  & ~new_n20027_;
  assign new_n20029_ = \b[52]  & ~new_n20021_;
  assign new_n20030_ = ~new_n20026_ & new_n20029_;
  assign new_n20031_ = new_n595_ & ~new_n20030_;
  assign new_n20032_ = ~new_n20028_ & new_n20031_;
  assign new_n20033_ = ~new_n20020_ & new_n20032_;
  assign new_n20034_ = new_n288_ & ~new_n20027_;
  assign \quotient[11]  = new_n20033_ | new_n20034_;
  assign new_n20036_ = ~new_n19322_ & new_n20018_;
  assign new_n20037_ = ~new_n20014_ & new_n20036_;
  assign new_n20038_ = ~new_n20015_ & ~new_n20018_;
  assign new_n20039_ = ~new_n20037_ & ~new_n20038_;
  assign new_n20040_ = \quotient[11]  & ~new_n20039_;
  assign new_n20041_ = ~new_n19312_ & ~new_n20034_;
  assign new_n20042_ = ~new_n20033_ & new_n20041_;
  assign new_n20043_ = ~new_n20040_ & ~new_n20042_;
  assign new_n20044_ = ~\b[52]  & ~new_n20043_;
  assign new_n20045_ = ~new_n19331_ & new_n20013_;
  assign new_n20046_ = ~new_n20009_ & new_n20045_;
  assign new_n20047_ = ~new_n20010_ & ~new_n20013_;
  assign new_n20048_ = ~new_n20046_ & ~new_n20047_;
  assign new_n20049_ = \quotient[11]  & ~new_n20048_;
  assign new_n20050_ = ~new_n19321_ & ~new_n20034_;
  assign new_n20051_ = ~new_n20033_ & new_n20050_;
  assign new_n20052_ = ~new_n20049_ & ~new_n20051_;
  assign new_n20053_ = ~\b[51]  & ~new_n20052_;
  assign new_n20054_ = ~new_n19340_ & new_n20008_;
  assign new_n20055_ = ~new_n20004_ & new_n20054_;
  assign new_n20056_ = ~new_n20005_ & ~new_n20008_;
  assign new_n20057_ = ~new_n20055_ & ~new_n20056_;
  assign new_n20058_ = \quotient[11]  & ~new_n20057_;
  assign new_n20059_ = ~new_n19330_ & ~new_n20034_;
  assign new_n20060_ = ~new_n20033_ & new_n20059_;
  assign new_n20061_ = ~new_n20058_ & ~new_n20060_;
  assign new_n20062_ = ~\b[50]  & ~new_n20061_;
  assign new_n20063_ = ~new_n19349_ & new_n20003_;
  assign new_n20064_ = ~new_n19999_ & new_n20063_;
  assign new_n20065_ = ~new_n20000_ & ~new_n20003_;
  assign new_n20066_ = ~new_n20064_ & ~new_n20065_;
  assign new_n20067_ = \quotient[11]  & ~new_n20066_;
  assign new_n20068_ = ~new_n19339_ & ~new_n20034_;
  assign new_n20069_ = ~new_n20033_ & new_n20068_;
  assign new_n20070_ = ~new_n20067_ & ~new_n20069_;
  assign new_n20071_ = ~\b[49]  & ~new_n20070_;
  assign new_n20072_ = ~new_n19358_ & new_n19998_;
  assign new_n20073_ = ~new_n19994_ & new_n20072_;
  assign new_n20074_ = ~new_n19995_ & ~new_n19998_;
  assign new_n20075_ = ~new_n20073_ & ~new_n20074_;
  assign new_n20076_ = \quotient[11]  & ~new_n20075_;
  assign new_n20077_ = ~new_n19348_ & ~new_n20034_;
  assign new_n20078_ = ~new_n20033_ & new_n20077_;
  assign new_n20079_ = ~new_n20076_ & ~new_n20078_;
  assign new_n20080_ = ~\b[48]  & ~new_n20079_;
  assign new_n20081_ = ~new_n19367_ & new_n19993_;
  assign new_n20082_ = ~new_n19989_ & new_n20081_;
  assign new_n20083_ = ~new_n19990_ & ~new_n19993_;
  assign new_n20084_ = ~new_n20082_ & ~new_n20083_;
  assign new_n20085_ = \quotient[11]  & ~new_n20084_;
  assign new_n20086_ = ~new_n19357_ & ~new_n20034_;
  assign new_n20087_ = ~new_n20033_ & new_n20086_;
  assign new_n20088_ = ~new_n20085_ & ~new_n20087_;
  assign new_n20089_ = ~\b[47]  & ~new_n20088_;
  assign new_n20090_ = ~new_n19376_ & new_n19988_;
  assign new_n20091_ = ~new_n19984_ & new_n20090_;
  assign new_n20092_ = ~new_n19985_ & ~new_n19988_;
  assign new_n20093_ = ~new_n20091_ & ~new_n20092_;
  assign new_n20094_ = \quotient[11]  & ~new_n20093_;
  assign new_n20095_ = ~new_n19366_ & ~new_n20034_;
  assign new_n20096_ = ~new_n20033_ & new_n20095_;
  assign new_n20097_ = ~new_n20094_ & ~new_n20096_;
  assign new_n20098_ = ~\b[46]  & ~new_n20097_;
  assign new_n20099_ = ~new_n19385_ & new_n19983_;
  assign new_n20100_ = ~new_n19979_ & new_n20099_;
  assign new_n20101_ = ~new_n19980_ & ~new_n19983_;
  assign new_n20102_ = ~new_n20100_ & ~new_n20101_;
  assign new_n20103_ = \quotient[11]  & ~new_n20102_;
  assign new_n20104_ = ~new_n19375_ & ~new_n20034_;
  assign new_n20105_ = ~new_n20033_ & new_n20104_;
  assign new_n20106_ = ~new_n20103_ & ~new_n20105_;
  assign new_n20107_ = ~\b[45]  & ~new_n20106_;
  assign new_n20108_ = ~new_n19394_ & new_n19978_;
  assign new_n20109_ = ~new_n19974_ & new_n20108_;
  assign new_n20110_ = ~new_n19975_ & ~new_n19978_;
  assign new_n20111_ = ~new_n20109_ & ~new_n20110_;
  assign new_n20112_ = \quotient[11]  & ~new_n20111_;
  assign new_n20113_ = ~new_n19384_ & ~new_n20034_;
  assign new_n20114_ = ~new_n20033_ & new_n20113_;
  assign new_n20115_ = ~new_n20112_ & ~new_n20114_;
  assign new_n20116_ = ~\b[44]  & ~new_n20115_;
  assign new_n20117_ = ~new_n19403_ & new_n19973_;
  assign new_n20118_ = ~new_n19969_ & new_n20117_;
  assign new_n20119_ = ~new_n19970_ & ~new_n19973_;
  assign new_n20120_ = ~new_n20118_ & ~new_n20119_;
  assign new_n20121_ = \quotient[11]  & ~new_n20120_;
  assign new_n20122_ = ~new_n19393_ & ~new_n20034_;
  assign new_n20123_ = ~new_n20033_ & new_n20122_;
  assign new_n20124_ = ~new_n20121_ & ~new_n20123_;
  assign new_n20125_ = ~\b[43]  & ~new_n20124_;
  assign new_n20126_ = ~new_n19412_ & new_n19968_;
  assign new_n20127_ = ~new_n19964_ & new_n20126_;
  assign new_n20128_ = ~new_n19965_ & ~new_n19968_;
  assign new_n20129_ = ~new_n20127_ & ~new_n20128_;
  assign new_n20130_ = \quotient[11]  & ~new_n20129_;
  assign new_n20131_ = ~new_n19402_ & ~new_n20034_;
  assign new_n20132_ = ~new_n20033_ & new_n20131_;
  assign new_n20133_ = ~new_n20130_ & ~new_n20132_;
  assign new_n20134_ = ~\b[42]  & ~new_n20133_;
  assign new_n20135_ = ~new_n19421_ & new_n19963_;
  assign new_n20136_ = ~new_n19959_ & new_n20135_;
  assign new_n20137_ = ~new_n19960_ & ~new_n19963_;
  assign new_n20138_ = ~new_n20136_ & ~new_n20137_;
  assign new_n20139_ = \quotient[11]  & ~new_n20138_;
  assign new_n20140_ = ~new_n19411_ & ~new_n20034_;
  assign new_n20141_ = ~new_n20033_ & new_n20140_;
  assign new_n20142_ = ~new_n20139_ & ~new_n20141_;
  assign new_n20143_ = ~\b[41]  & ~new_n20142_;
  assign new_n20144_ = ~new_n19430_ & new_n19958_;
  assign new_n20145_ = ~new_n19954_ & new_n20144_;
  assign new_n20146_ = ~new_n19955_ & ~new_n19958_;
  assign new_n20147_ = ~new_n20145_ & ~new_n20146_;
  assign new_n20148_ = \quotient[11]  & ~new_n20147_;
  assign new_n20149_ = ~new_n19420_ & ~new_n20034_;
  assign new_n20150_ = ~new_n20033_ & new_n20149_;
  assign new_n20151_ = ~new_n20148_ & ~new_n20150_;
  assign new_n20152_ = ~\b[40]  & ~new_n20151_;
  assign new_n20153_ = ~new_n19439_ & new_n19953_;
  assign new_n20154_ = ~new_n19949_ & new_n20153_;
  assign new_n20155_ = ~new_n19950_ & ~new_n19953_;
  assign new_n20156_ = ~new_n20154_ & ~new_n20155_;
  assign new_n20157_ = \quotient[11]  & ~new_n20156_;
  assign new_n20158_ = ~new_n19429_ & ~new_n20034_;
  assign new_n20159_ = ~new_n20033_ & new_n20158_;
  assign new_n20160_ = ~new_n20157_ & ~new_n20159_;
  assign new_n20161_ = ~\b[39]  & ~new_n20160_;
  assign new_n20162_ = ~new_n19448_ & new_n19948_;
  assign new_n20163_ = ~new_n19944_ & new_n20162_;
  assign new_n20164_ = ~new_n19945_ & ~new_n19948_;
  assign new_n20165_ = ~new_n20163_ & ~new_n20164_;
  assign new_n20166_ = \quotient[11]  & ~new_n20165_;
  assign new_n20167_ = ~new_n19438_ & ~new_n20034_;
  assign new_n20168_ = ~new_n20033_ & new_n20167_;
  assign new_n20169_ = ~new_n20166_ & ~new_n20168_;
  assign new_n20170_ = ~\b[38]  & ~new_n20169_;
  assign new_n20171_ = ~new_n19457_ & new_n19943_;
  assign new_n20172_ = ~new_n19939_ & new_n20171_;
  assign new_n20173_ = ~new_n19940_ & ~new_n19943_;
  assign new_n20174_ = ~new_n20172_ & ~new_n20173_;
  assign new_n20175_ = \quotient[11]  & ~new_n20174_;
  assign new_n20176_ = ~new_n19447_ & ~new_n20034_;
  assign new_n20177_ = ~new_n20033_ & new_n20176_;
  assign new_n20178_ = ~new_n20175_ & ~new_n20177_;
  assign new_n20179_ = ~\b[37]  & ~new_n20178_;
  assign new_n20180_ = ~new_n19466_ & new_n19938_;
  assign new_n20181_ = ~new_n19934_ & new_n20180_;
  assign new_n20182_ = ~new_n19935_ & ~new_n19938_;
  assign new_n20183_ = ~new_n20181_ & ~new_n20182_;
  assign new_n20184_ = \quotient[11]  & ~new_n20183_;
  assign new_n20185_ = ~new_n19456_ & ~new_n20034_;
  assign new_n20186_ = ~new_n20033_ & new_n20185_;
  assign new_n20187_ = ~new_n20184_ & ~new_n20186_;
  assign new_n20188_ = ~\b[36]  & ~new_n20187_;
  assign new_n20189_ = ~new_n19475_ & new_n19933_;
  assign new_n20190_ = ~new_n19929_ & new_n20189_;
  assign new_n20191_ = ~new_n19930_ & ~new_n19933_;
  assign new_n20192_ = ~new_n20190_ & ~new_n20191_;
  assign new_n20193_ = \quotient[11]  & ~new_n20192_;
  assign new_n20194_ = ~new_n19465_ & ~new_n20034_;
  assign new_n20195_ = ~new_n20033_ & new_n20194_;
  assign new_n20196_ = ~new_n20193_ & ~new_n20195_;
  assign new_n20197_ = ~\b[35]  & ~new_n20196_;
  assign new_n20198_ = ~new_n19484_ & new_n19928_;
  assign new_n20199_ = ~new_n19924_ & new_n20198_;
  assign new_n20200_ = ~new_n19925_ & ~new_n19928_;
  assign new_n20201_ = ~new_n20199_ & ~new_n20200_;
  assign new_n20202_ = \quotient[11]  & ~new_n20201_;
  assign new_n20203_ = ~new_n19474_ & ~new_n20034_;
  assign new_n20204_ = ~new_n20033_ & new_n20203_;
  assign new_n20205_ = ~new_n20202_ & ~new_n20204_;
  assign new_n20206_ = ~\b[34]  & ~new_n20205_;
  assign new_n20207_ = ~new_n19493_ & new_n19923_;
  assign new_n20208_ = ~new_n19919_ & new_n20207_;
  assign new_n20209_ = ~new_n19920_ & ~new_n19923_;
  assign new_n20210_ = ~new_n20208_ & ~new_n20209_;
  assign new_n20211_ = \quotient[11]  & ~new_n20210_;
  assign new_n20212_ = ~new_n19483_ & ~new_n20034_;
  assign new_n20213_ = ~new_n20033_ & new_n20212_;
  assign new_n20214_ = ~new_n20211_ & ~new_n20213_;
  assign new_n20215_ = ~\b[33]  & ~new_n20214_;
  assign new_n20216_ = ~new_n19502_ & new_n19918_;
  assign new_n20217_ = ~new_n19914_ & new_n20216_;
  assign new_n20218_ = ~new_n19915_ & ~new_n19918_;
  assign new_n20219_ = ~new_n20217_ & ~new_n20218_;
  assign new_n20220_ = \quotient[11]  & ~new_n20219_;
  assign new_n20221_ = ~new_n19492_ & ~new_n20034_;
  assign new_n20222_ = ~new_n20033_ & new_n20221_;
  assign new_n20223_ = ~new_n20220_ & ~new_n20222_;
  assign new_n20224_ = ~\b[32]  & ~new_n20223_;
  assign new_n20225_ = ~new_n19511_ & new_n19913_;
  assign new_n20226_ = ~new_n19909_ & new_n20225_;
  assign new_n20227_ = ~new_n19910_ & ~new_n19913_;
  assign new_n20228_ = ~new_n20226_ & ~new_n20227_;
  assign new_n20229_ = \quotient[11]  & ~new_n20228_;
  assign new_n20230_ = ~new_n19501_ & ~new_n20034_;
  assign new_n20231_ = ~new_n20033_ & new_n20230_;
  assign new_n20232_ = ~new_n20229_ & ~new_n20231_;
  assign new_n20233_ = ~\b[31]  & ~new_n20232_;
  assign new_n20234_ = ~new_n19520_ & new_n19908_;
  assign new_n20235_ = ~new_n19904_ & new_n20234_;
  assign new_n20236_ = ~new_n19905_ & ~new_n19908_;
  assign new_n20237_ = ~new_n20235_ & ~new_n20236_;
  assign new_n20238_ = \quotient[11]  & ~new_n20237_;
  assign new_n20239_ = ~new_n19510_ & ~new_n20034_;
  assign new_n20240_ = ~new_n20033_ & new_n20239_;
  assign new_n20241_ = ~new_n20238_ & ~new_n20240_;
  assign new_n20242_ = ~\b[30]  & ~new_n20241_;
  assign new_n20243_ = ~new_n19529_ & new_n19903_;
  assign new_n20244_ = ~new_n19899_ & new_n20243_;
  assign new_n20245_ = ~new_n19900_ & ~new_n19903_;
  assign new_n20246_ = ~new_n20244_ & ~new_n20245_;
  assign new_n20247_ = \quotient[11]  & ~new_n20246_;
  assign new_n20248_ = ~new_n19519_ & ~new_n20034_;
  assign new_n20249_ = ~new_n20033_ & new_n20248_;
  assign new_n20250_ = ~new_n20247_ & ~new_n20249_;
  assign new_n20251_ = ~\b[29]  & ~new_n20250_;
  assign new_n20252_ = ~new_n19538_ & new_n19898_;
  assign new_n20253_ = ~new_n19894_ & new_n20252_;
  assign new_n20254_ = ~new_n19895_ & ~new_n19898_;
  assign new_n20255_ = ~new_n20253_ & ~new_n20254_;
  assign new_n20256_ = \quotient[11]  & ~new_n20255_;
  assign new_n20257_ = ~new_n19528_ & ~new_n20034_;
  assign new_n20258_ = ~new_n20033_ & new_n20257_;
  assign new_n20259_ = ~new_n20256_ & ~new_n20258_;
  assign new_n20260_ = ~\b[28]  & ~new_n20259_;
  assign new_n20261_ = ~new_n19547_ & new_n19893_;
  assign new_n20262_ = ~new_n19889_ & new_n20261_;
  assign new_n20263_ = ~new_n19890_ & ~new_n19893_;
  assign new_n20264_ = ~new_n20262_ & ~new_n20263_;
  assign new_n20265_ = \quotient[11]  & ~new_n20264_;
  assign new_n20266_ = ~new_n19537_ & ~new_n20034_;
  assign new_n20267_ = ~new_n20033_ & new_n20266_;
  assign new_n20268_ = ~new_n20265_ & ~new_n20267_;
  assign new_n20269_ = ~\b[27]  & ~new_n20268_;
  assign new_n20270_ = ~new_n19556_ & new_n19888_;
  assign new_n20271_ = ~new_n19884_ & new_n20270_;
  assign new_n20272_ = ~new_n19885_ & ~new_n19888_;
  assign new_n20273_ = ~new_n20271_ & ~new_n20272_;
  assign new_n20274_ = \quotient[11]  & ~new_n20273_;
  assign new_n20275_ = ~new_n19546_ & ~new_n20034_;
  assign new_n20276_ = ~new_n20033_ & new_n20275_;
  assign new_n20277_ = ~new_n20274_ & ~new_n20276_;
  assign new_n20278_ = ~\b[26]  & ~new_n20277_;
  assign new_n20279_ = ~new_n19565_ & new_n19883_;
  assign new_n20280_ = ~new_n19879_ & new_n20279_;
  assign new_n20281_ = ~new_n19880_ & ~new_n19883_;
  assign new_n20282_ = ~new_n20280_ & ~new_n20281_;
  assign new_n20283_ = \quotient[11]  & ~new_n20282_;
  assign new_n20284_ = ~new_n19555_ & ~new_n20034_;
  assign new_n20285_ = ~new_n20033_ & new_n20284_;
  assign new_n20286_ = ~new_n20283_ & ~new_n20285_;
  assign new_n20287_ = ~\b[25]  & ~new_n20286_;
  assign new_n20288_ = ~new_n19574_ & new_n19878_;
  assign new_n20289_ = ~new_n19874_ & new_n20288_;
  assign new_n20290_ = ~new_n19875_ & ~new_n19878_;
  assign new_n20291_ = ~new_n20289_ & ~new_n20290_;
  assign new_n20292_ = \quotient[11]  & ~new_n20291_;
  assign new_n20293_ = ~new_n19564_ & ~new_n20034_;
  assign new_n20294_ = ~new_n20033_ & new_n20293_;
  assign new_n20295_ = ~new_n20292_ & ~new_n20294_;
  assign new_n20296_ = ~\b[24]  & ~new_n20295_;
  assign new_n20297_ = ~new_n19583_ & new_n19873_;
  assign new_n20298_ = ~new_n19869_ & new_n20297_;
  assign new_n20299_ = ~new_n19870_ & ~new_n19873_;
  assign new_n20300_ = ~new_n20298_ & ~new_n20299_;
  assign new_n20301_ = \quotient[11]  & ~new_n20300_;
  assign new_n20302_ = ~new_n19573_ & ~new_n20034_;
  assign new_n20303_ = ~new_n20033_ & new_n20302_;
  assign new_n20304_ = ~new_n20301_ & ~new_n20303_;
  assign new_n20305_ = ~\b[23]  & ~new_n20304_;
  assign new_n20306_ = ~new_n19592_ & new_n19868_;
  assign new_n20307_ = ~new_n19864_ & new_n20306_;
  assign new_n20308_ = ~new_n19865_ & ~new_n19868_;
  assign new_n20309_ = ~new_n20307_ & ~new_n20308_;
  assign new_n20310_ = \quotient[11]  & ~new_n20309_;
  assign new_n20311_ = ~new_n19582_ & ~new_n20034_;
  assign new_n20312_ = ~new_n20033_ & new_n20311_;
  assign new_n20313_ = ~new_n20310_ & ~new_n20312_;
  assign new_n20314_ = ~\b[22]  & ~new_n20313_;
  assign new_n20315_ = ~new_n19601_ & new_n19863_;
  assign new_n20316_ = ~new_n19859_ & new_n20315_;
  assign new_n20317_ = ~new_n19860_ & ~new_n19863_;
  assign new_n20318_ = ~new_n20316_ & ~new_n20317_;
  assign new_n20319_ = \quotient[11]  & ~new_n20318_;
  assign new_n20320_ = ~new_n19591_ & ~new_n20034_;
  assign new_n20321_ = ~new_n20033_ & new_n20320_;
  assign new_n20322_ = ~new_n20319_ & ~new_n20321_;
  assign new_n20323_ = ~\b[21]  & ~new_n20322_;
  assign new_n20324_ = ~new_n19610_ & new_n19858_;
  assign new_n20325_ = ~new_n19854_ & new_n20324_;
  assign new_n20326_ = ~new_n19855_ & ~new_n19858_;
  assign new_n20327_ = ~new_n20325_ & ~new_n20326_;
  assign new_n20328_ = \quotient[11]  & ~new_n20327_;
  assign new_n20329_ = ~new_n19600_ & ~new_n20034_;
  assign new_n20330_ = ~new_n20033_ & new_n20329_;
  assign new_n20331_ = ~new_n20328_ & ~new_n20330_;
  assign new_n20332_ = ~\b[20]  & ~new_n20331_;
  assign new_n20333_ = ~new_n19619_ & new_n19853_;
  assign new_n20334_ = ~new_n19849_ & new_n20333_;
  assign new_n20335_ = ~new_n19850_ & ~new_n19853_;
  assign new_n20336_ = ~new_n20334_ & ~new_n20335_;
  assign new_n20337_ = \quotient[11]  & ~new_n20336_;
  assign new_n20338_ = ~new_n19609_ & ~new_n20034_;
  assign new_n20339_ = ~new_n20033_ & new_n20338_;
  assign new_n20340_ = ~new_n20337_ & ~new_n20339_;
  assign new_n20341_ = ~\b[19]  & ~new_n20340_;
  assign new_n20342_ = ~new_n19628_ & new_n19848_;
  assign new_n20343_ = ~new_n19844_ & new_n20342_;
  assign new_n20344_ = ~new_n19845_ & ~new_n19848_;
  assign new_n20345_ = ~new_n20343_ & ~new_n20344_;
  assign new_n20346_ = \quotient[11]  & ~new_n20345_;
  assign new_n20347_ = ~new_n19618_ & ~new_n20034_;
  assign new_n20348_ = ~new_n20033_ & new_n20347_;
  assign new_n20349_ = ~new_n20346_ & ~new_n20348_;
  assign new_n20350_ = ~\b[18]  & ~new_n20349_;
  assign new_n20351_ = ~new_n19637_ & new_n19843_;
  assign new_n20352_ = ~new_n19839_ & new_n20351_;
  assign new_n20353_ = ~new_n19840_ & ~new_n19843_;
  assign new_n20354_ = ~new_n20352_ & ~new_n20353_;
  assign new_n20355_ = \quotient[11]  & ~new_n20354_;
  assign new_n20356_ = ~new_n19627_ & ~new_n20034_;
  assign new_n20357_ = ~new_n20033_ & new_n20356_;
  assign new_n20358_ = ~new_n20355_ & ~new_n20357_;
  assign new_n20359_ = ~\b[17]  & ~new_n20358_;
  assign new_n20360_ = ~new_n19646_ & new_n19838_;
  assign new_n20361_ = ~new_n19834_ & new_n20360_;
  assign new_n20362_ = ~new_n19835_ & ~new_n19838_;
  assign new_n20363_ = ~new_n20361_ & ~new_n20362_;
  assign new_n20364_ = \quotient[11]  & ~new_n20363_;
  assign new_n20365_ = ~new_n19636_ & ~new_n20034_;
  assign new_n20366_ = ~new_n20033_ & new_n20365_;
  assign new_n20367_ = ~new_n20364_ & ~new_n20366_;
  assign new_n20368_ = ~\b[16]  & ~new_n20367_;
  assign new_n20369_ = ~new_n19655_ & new_n19833_;
  assign new_n20370_ = ~new_n19829_ & new_n20369_;
  assign new_n20371_ = ~new_n19830_ & ~new_n19833_;
  assign new_n20372_ = ~new_n20370_ & ~new_n20371_;
  assign new_n20373_ = \quotient[11]  & ~new_n20372_;
  assign new_n20374_ = ~new_n19645_ & ~new_n20034_;
  assign new_n20375_ = ~new_n20033_ & new_n20374_;
  assign new_n20376_ = ~new_n20373_ & ~new_n20375_;
  assign new_n20377_ = ~\b[15]  & ~new_n20376_;
  assign new_n20378_ = ~new_n19664_ & new_n19828_;
  assign new_n20379_ = ~new_n19824_ & new_n20378_;
  assign new_n20380_ = ~new_n19825_ & ~new_n19828_;
  assign new_n20381_ = ~new_n20379_ & ~new_n20380_;
  assign new_n20382_ = \quotient[11]  & ~new_n20381_;
  assign new_n20383_ = ~new_n19654_ & ~new_n20034_;
  assign new_n20384_ = ~new_n20033_ & new_n20383_;
  assign new_n20385_ = ~new_n20382_ & ~new_n20384_;
  assign new_n20386_ = ~\b[14]  & ~new_n20385_;
  assign new_n20387_ = ~new_n19673_ & new_n19823_;
  assign new_n20388_ = ~new_n19819_ & new_n20387_;
  assign new_n20389_ = ~new_n19820_ & ~new_n19823_;
  assign new_n20390_ = ~new_n20388_ & ~new_n20389_;
  assign new_n20391_ = \quotient[11]  & ~new_n20390_;
  assign new_n20392_ = ~new_n19663_ & ~new_n20034_;
  assign new_n20393_ = ~new_n20033_ & new_n20392_;
  assign new_n20394_ = ~new_n20391_ & ~new_n20393_;
  assign new_n20395_ = ~\b[13]  & ~new_n20394_;
  assign new_n20396_ = ~new_n19682_ & new_n19818_;
  assign new_n20397_ = ~new_n19814_ & new_n20396_;
  assign new_n20398_ = ~new_n19815_ & ~new_n19818_;
  assign new_n20399_ = ~new_n20397_ & ~new_n20398_;
  assign new_n20400_ = \quotient[11]  & ~new_n20399_;
  assign new_n20401_ = ~new_n19672_ & ~new_n20034_;
  assign new_n20402_ = ~new_n20033_ & new_n20401_;
  assign new_n20403_ = ~new_n20400_ & ~new_n20402_;
  assign new_n20404_ = ~\b[12]  & ~new_n20403_;
  assign new_n20405_ = ~new_n19691_ & new_n19813_;
  assign new_n20406_ = ~new_n19809_ & new_n20405_;
  assign new_n20407_ = ~new_n19810_ & ~new_n19813_;
  assign new_n20408_ = ~new_n20406_ & ~new_n20407_;
  assign new_n20409_ = \quotient[11]  & ~new_n20408_;
  assign new_n20410_ = ~new_n19681_ & ~new_n20034_;
  assign new_n20411_ = ~new_n20033_ & new_n20410_;
  assign new_n20412_ = ~new_n20409_ & ~new_n20411_;
  assign new_n20413_ = ~\b[11]  & ~new_n20412_;
  assign new_n20414_ = ~new_n19700_ & new_n19808_;
  assign new_n20415_ = ~new_n19804_ & new_n20414_;
  assign new_n20416_ = ~new_n19805_ & ~new_n19808_;
  assign new_n20417_ = ~new_n20415_ & ~new_n20416_;
  assign new_n20418_ = \quotient[11]  & ~new_n20417_;
  assign new_n20419_ = ~new_n19690_ & ~new_n20034_;
  assign new_n20420_ = ~new_n20033_ & new_n20419_;
  assign new_n20421_ = ~new_n20418_ & ~new_n20420_;
  assign new_n20422_ = ~\b[10]  & ~new_n20421_;
  assign new_n20423_ = ~new_n19709_ & new_n19803_;
  assign new_n20424_ = ~new_n19799_ & new_n20423_;
  assign new_n20425_ = ~new_n19800_ & ~new_n19803_;
  assign new_n20426_ = ~new_n20424_ & ~new_n20425_;
  assign new_n20427_ = \quotient[11]  & ~new_n20426_;
  assign new_n20428_ = ~new_n19699_ & ~new_n20034_;
  assign new_n20429_ = ~new_n20033_ & new_n20428_;
  assign new_n20430_ = ~new_n20427_ & ~new_n20429_;
  assign new_n20431_ = ~\b[9]  & ~new_n20430_;
  assign new_n20432_ = ~new_n19718_ & new_n19798_;
  assign new_n20433_ = ~new_n19794_ & new_n20432_;
  assign new_n20434_ = ~new_n19795_ & ~new_n19798_;
  assign new_n20435_ = ~new_n20433_ & ~new_n20434_;
  assign new_n20436_ = \quotient[11]  & ~new_n20435_;
  assign new_n20437_ = ~new_n19708_ & ~new_n20034_;
  assign new_n20438_ = ~new_n20033_ & new_n20437_;
  assign new_n20439_ = ~new_n20436_ & ~new_n20438_;
  assign new_n20440_ = ~\b[8]  & ~new_n20439_;
  assign new_n20441_ = ~new_n19727_ & new_n19793_;
  assign new_n20442_ = ~new_n19789_ & new_n20441_;
  assign new_n20443_ = ~new_n19790_ & ~new_n19793_;
  assign new_n20444_ = ~new_n20442_ & ~new_n20443_;
  assign new_n20445_ = \quotient[11]  & ~new_n20444_;
  assign new_n20446_ = ~new_n19717_ & ~new_n20034_;
  assign new_n20447_ = ~new_n20033_ & new_n20446_;
  assign new_n20448_ = ~new_n20445_ & ~new_n20447_;
  assign new_n20449_ = ~\b[7]  & ~new_n20448_;
  assign new_n20450_ = ~new_n19736_ & new_n19788_;
  assign new_n20451_ = ~new_n19784_ & new_n20450_;
  assign new_n20452_ = ~new_n19785_ & ~new_n19788_;
  assign new_n20453_ = ~new_n20451_ & ~new_n20452_;
  assign new_n20454_ = \quotient[11]  & ~new_n20453_;
  assign new_n20455_ = ~new_n19726_ & ~new_n20034_;
  assign new_n20456_ = ~new_n20033_ & new_n20455_;
  assign new_n20457_ = ~new_n20454_ & ~new_n20456_;
  assign new_n20458_ = ~\b[6]  & ~new_n20457_;
  assign new_n20459_ = ~new_n19745_ & new_n19783_;
  assign new_n20460_ = ~new_n19779_ & new_n20459_;
  assign new_n20461_ = ~new_n19780_ & ~new_n19783_;
  assign new_n20462_ = ~new_n20460_ & ~new_n20461_;
  assign new_n20463_ = \quotient[11]  & ~new_n20462_;
  assign new_n20464_ = ~new_n19735_ & ~new_n20034_;
  assign new_n20465_ = ~new_n20033_ & new_n20464_;
  assign new_n20466_ = ~new_n20463_ & ~new_n20465_;
  assign new_n20467_ = ~\b[5]  & ~new_n20466_;
  assign new_n20468_ = ~new_n19753_ & new_n19778_;
  assign new_n20469_ = ~new_n19774_ & new_n20468_;
  assign new_n20470_ = ~new_n19775_ & ~new_n19778_;
  assign new_n20471_ = ~new_n20469_ & ~new_n20470_;
  assign new_n20472_ = \quotient[11]  & ~new_n20471_;
  assign new_n20473_ = ~new_n19744_ & ~new_n20034_;
  assign new_n20474_ = ~new_n20033_ & new_n20473_;
  assign new_n20475_ = ~new_n20472_ & ~new_n20474_;
  assign new_n20476_ = ~\b[4]  & ~new_n20475_;
  assign new_n20477_ = ~new_n19769_ & new_n19773_;
  assign new_n20478_ = ~new_n19768_ & new_n20477_;
  assign new_n20479_ = ~new_n19770_ & ~new_n19773_;
  assign new_n20480_ = ~new_n20478_ & ~new_n20479_;
  assign new_n20481_ = \quotient[11]  & ~new_n20480_;
  assign new_n20482_ = ~new_n19752_ & ~new_n20034_;
  assign new_n20483_ = ~new_n20033_ & new_n20482_;
  assign new_n20484_ = ~new_n20481_ & ~new_n20483_;
  assign new_n20485_ = ~\b[3]  & ~new_n20484_;
  assign new_n20486_ = ~new_n19765_ & new_n19767_;
  assign new_n20487_ = ~new_n19763_ & new_n20486_;
  assign new_n20488_ = ~new_n19768_ & ~new_n20487_;
  assign new_n20489_ = \quotient[11]  & new_n20488_;
  assign new_n20490_ = ~new_n19762_ & ~new_n20034_;
  assign new_n20491_ = ~new_n20033_ & new_n20490_;
  assign new_n20492_ = ~new_n20489_ & ~new_n20491_;
  assign new_n20493_ = ~\b[2]  & ~new_n20492_;
  assign new_n20494_ = \b[0]  & \quotient[11] ;
  assign new_n20495_ = \a[11]  & ~new_n20494_;
  assign new_n20496_ = new_n19767_ & \quotient[11] ;
  assign new_n20497_ = ~new_n20495_ & ~new_n20496_;
  assign new_n20498_ = \b[1]  & ~new_n20497_;
  assign new_n20499_ = ~\b[1]  & ~new_n20496_;
  assign new_n20500_ = ~new_n20495_ & new_n20499_;
  assign new_n20501_ = ~new_n20498_ & ~new_n20500_;
  assign new_n20502_ = ~\a[10]  & \b[0] ;
  assign new_n20503_ = ~new_n20501_ & ~new_n20502_;
  assign new_n20504_ = ~\b[1]  & ~new_n20497_;
  assign new_n20505_ = ~new_n20503_ & ~new_n20504_;
  assign new_n20506_ = \b[2]  & ~new_n20491_;
  assign new_n20507_ = ~new_n20489_ & new_n20506_;
  assign new_n20508_ = ~new_n20493_ & ~new_n20507_;
  assign new_n20509_ = ~new_n20505_ & new_n20508_;
  assign new_n20510_ = ~new_n20493_ & ~new_n20509_;
  assign new_n20511_ = \b[3]  & ~new_n20483_;
  assign new_n20512_ = ~new_n20481_ & new_n20511_;
  assign new_n20513_ = ~new_n20485_ & ~new_n20512_;
  assign new_n20514_ = ~new_n20510_ & new_n20513_;
  assign new_n20515_ = ~new_n20485_ & ~new_n20514_;
  assign new_n20516_ = \b[4]  & ~new_n20474_;
  assign new_n20517_ = ~new_n20472_ & new_n20516_;
  assign new_n20518_ = ~new_n20476_ & ~new_n20517_;
  assign new_n20519_ = ~new_n20515_ & new_n20518_;
  assign new_n20520_ = ~new_n20476_ & ~new_n20519_;
  assign new_n20521_ = \b[5]  & ~new_n20465_;
  assign new_n20522_ = ~new_n20463_ & new_n20521_;
  assign new_n20523_ = ~new_n20467_ & ~new_n20522_;
  assign new_n20524_ = ~new_n20520_ & new_n20523_;
  assign new_n20525_ = ~new_n20467_ & ~new_n20524_;
  assign new_n20526_ = \b[6]  & ~new_n20456_;
  assign new_n20527_ = ~new_n20454_ & new_n20526_;
  assign new_n20528_ = ~new_n20458_ & ~new_n20527_;
  assign new_n20529_ = ~new_n20525_ & new_n20528_;
  assign new_n20530_ = ~new_n20458_ & ~new_n20529_;
  assign new_n20531_ = \b[7]  & ~new_n20447_;
  assign new_n20532_ = ~new_n20445_ & new_n20531_;
  assign new_n20533_ = ~new_n20449_ & ~new_n20532_;
  assign new_n20534_ = ~new_n20530_ & new_n20533_;
  assign new_n20535_ = ~new_n20449_ & ~new_n20534_;
  assign new_n20536_ = \b[8]  & ~new_n20438_;
  assign new_n20537_ = ~new_n20436_ & new_n20536_;
  assign new_n20538_ = ~new_n20440_ & ~new_n20537_;
  assign new_n20539_ = ~new_n20535_ & new_n20538_;
  assign new_n20540_ = ~new_n20440_ & ~new_n20539_;
  assign new_n20541_ = \b[9]  & ~new_n20429_;
  assign new_n20542_ = ~new_n20427_ & new_n20541_;
  assign new_n20543_ = ~new_n20431_ & ~new_n20542_;
  assign new_n20544_ = ~new_n20540_ & new_n20543_;
  assign new_n20545_ = ~new_n20431_ & ~new_n20544_;
  assign new_n20546_ = \b[10]  & ~new_n20420_;
  assign new_n20547_ = ~new_n20418_ & new_n20546_;
  assign new_n20548_ = ~new_n20422_ & ~new_n20547_;
  assign new_n20549_ = ~new_n20545_ & new_n20548_;
  assign new_n20550_ = ~new_n20422_ & ~new_n20549_;
  assign new_n20551_ = \b[11]  & ~new_n20411_;
  assign new_n20552_ = ~new_n20409_ & new_n20551_;
  assign new_n20553_ = ~new_n20413_ & ~new_n20552_;
  assign new_n20554_ = ~new_n20550_ & new_n20553_;
  assign new_n20555_ = ~new_n20413_ & ~new_n20554_;
  assign new_n20556_ = \b[12]  & ~new_n20402_;
  assign new_n20557_ = ~new_n20400_ & new_n20556_;
  assign new_n20558_ = ~new_n20404_ & ~new_n20557_;
  assign new_n20559_ = ~new_n20555_ & new_n20558_;
  assign new_n20560_ = ~new_n20404_ & ~new_n20559_;
  assign new_n20561_ = \b[13]  & ~new_n20393_;
  assign new_n20562_ = ~new_n20391_ & new_n20561_;
  assign new_n20563_ = ~new_n20395_ & ~new_n20562_;
  assign new_n20564_ = ~new_n20560_ & new_n20563_;
  assign new_n20565_ = ~new_n20395_ & ~new_n20564_;
  assign new_n20566_ = \b[14]  & ~new_n20384_;
  assign new_n20567_ = ~new_n20382_ & new_n20566_;
  assign new_n20568_ = ~new_n20386_ & ~new_n20567_;
  assign new_n20569_ = ~new_n20565_ & new_n20568_;
  assign new_n20570_ = ~new_n20386_ & ~new_n20569_;
  assign new_n20571_ = \b[15]  & ~new_n20375_;
  assign new_n20572_ = ~new_n20373_ & new_n20571_;
  assign new_n20573_ = ~new_n20377_ & ~new_n20572_;
  assign new_n20574_ = ~new_n20570_ & new_n20573_;
  assign new_n20575_ = ~new_n20377_ & ~new_n20574_;
  assign new_n20576_ = \b[16]  & ~new_n20366_;
  assign new_n20577_ = ~new_n20364_ & new_n20576_;
  assign new_n20578_ = ~new_n20368_ & ~new_n20577_;
  assign new_n20579_ = ~new_n20575_ & new_n20578_;
  assign new_n20580_ = ~new_n20368_ & ~new_n20579_;
  assign new_n20581_ = \b[17]  & ~new_n20357_;
  assign new_n20582_ = ~new_n20355_ & new_n20581_;
  assign new_n20583_ = ~new_n20359_ & ~new_n20582_;
  assign new_n20584_ = ~new_n20580_ & new_n20583_;
  assign new_n20585_ = ~new_n20359_ & ~new_n20584_;
  assign new_n20586_ = \b[18]  & ~new_n20348_;
  assign new_n20587_ = ~new_n20346_ & new_n20586_;
  assign new_n20588_ = ~new_n20350_ & ~new_n20587_;
  assign new_n20589_ = ~new_n20585_ & new_n20588_;
  assign new_n20590_ = ~new_n20350_ & ~new_n20589_;
  assign new_n20591_ = \b[19]  & ~new_n20339_;
  assign new_n20592_ = ~new_n20337_ & new_n20591_;
  assign new_n20593_ = ~new_n20341_ & ~new_n20592_;
  assign new_n20594_ = ~new_n20590_ & new_n20593_;
  assign new_n20595_ = ~new_n20341_ & ~new_n20594_;
  assign new_n20596_ = \b[20]  & ~new_n20330_;
  assign new_n20597_ = ~new_n20328_ & new_n20596_;
  assign new_n20598_ = ~new_n20332_ & ~new_n20597_;
  assign new_n20599_ = ~new_n20595_ & new_n20598_;
  assign new_n20600_ = ~new_n20332_ & ~new_n20599_;
  assign new_n20601_ = \b[21]  & ~new_n20321_;
  assign new_n20602_ = ~new_n20319_ & new_n20601_;
  assign new_n20603_ = ~new_n20323_ & ~new_n20602_;
  assign new_n20604_ = ~new_n20600_ & new_n20603_;
  assign new_n20605_ = ~new_n20323_ & ~new_n20604_;
  assign new_n20606_ = \b[22]  & ~new_n20312_;
  assign new_n20607_ = ~new_n20310_ & new_n20606_;
  assign new_n20608_ = ~new_n20314_ & ~new_n20607_;
  assign new_n20609_ = ~new_n20605_ & new_n20608_;
  assign new_n20610_ = ~new_n20314_ & ~new_n20609_;
  assign new_n20611_ = \b[23]  & ~new_n20303_;
  assign new_n20612_ = ~new_n20301_ & new_n20611_;
  assign new_n20613_ = ~new_n20305_ & ~new_n20612_;
  assign new_n20614_ = ~new_n20610_ & new_n20613_;
  assign new_n20615_ = ~new_n20305_ & ~new_n20614_;
  assign new_n20616_ = \b[24]  & ~new_n20294_;
  assign new_n20617_ = ~new_n20292_ & new_n20616_;
  assign new_n20618_ = ~new_n20296_ & ~new_n20617_;
  assign new_n20619_ = ~new_n20615_ & new_n20618_;
  assign new_n20620_ = ~new_n20296_ & ~new_n20619_;
  assign new_n20621_ = \b[25]  & ~new_n20285_;
  assign new_n20622_ = ~new_n20283_ & new_n20621_;
  assign new_n20623_ = ~new_n20287_ & ~new_n20622_;
  assign new_n20624_ = ~new_n20620_ & new_n20623_;
  assign new_n20625_ = ~new_n20287_ & ~new_n20624_;
  assign new_n20626_ = \b[26]  & ~new_n20276_;
  assign new_n20627_ = ~new_n20274_ & new_n20626_;
  assign new_n20628_ = ~new_n20278_ & ~new_n20627_;
  assign new_n20629_ = ~new_n20625_ & new_n20628_;
  assign new_n20630_ = ~new_n20278_ & ~new_n20629_;
  assign new_n20631_ = \b[27]  & ~new_n20267_;
  assign new_n20632_ = ~new_n20265_ & new_n20631_;
  assign new_n20633_ = ~new_n20269_ & ~new_n20632_;
  assign new_n20634_ = ~new_n20630_ & new_n20633_;
  assign new_n20635_ = ~new_n20269_ & ~new_n20634_;
  assign new_n20636_ = \b[28]  & ~new_n20258_;
  assign new_n20637_ = ~new_n20256_ & new_n20636_;
  assign new_n20638_ = ~new_n20260_ & ~new_n20637_;
  assign new_n20639_ = ~new_n20635_ & new_n20638_;
  assign new_n20640_ = ~new_n20260_ & ~new_n20639_;
  assign new_n20641_ = \b[29]  & ~new_n20249_;
  assign new_n20642_ = ~new_n20247_ & new_n20641_;
  assign new_n20643_ = ~new_n20251_ & ~new_n20642_;
  assign new_n20644_ = ~new_n20640_ & new_n20643_;
  assign new_n20645_ = ~new_n20251_ & ~new_n20644_;
  assign new_n20646_ = \b[30]  & ~new_n20240_;
  assign new_n20647_ = ~new_n20238_ & new_n20646_;
  assign new_n20648_ = ~new_n20242_ & ~new_n20647_;
  assign new_n20649_ = ~new_n20645_ & new_n20648_;
  assign new_n20650_ = ~new_n20242_ & ~new_n20649_;
  assign new_n20651_ = \b[31]  & ~new_n20231_;
  assign new_n20652_ = ~new_n20229_ & new_n20651_;
  assign new_n20653_ = ~new_n20233_ & ~new_n20652_;
  assign new_n20654_ = ~new_n20650_ & new_n20653_;
  assign new_n20655_ = ~new_n20233_ & ~new_n20654_;
  assign new_n20656_ = \b[32]  & ~new_n20222_;
  assign new_n20657_ = ~new_n20220_ & new_n20656_;
  assign new_n20658_ = ~new_n20224_ & ~new_n20657_;
  assign new_n20659_ = ~new_n20655_ & new_n20658_;
  assign new_n20660_ = ~new_n20224_ & ~new_n20659_;
  assign new_n20661_ = \b[33]  & ~new_n20213_;
  assign new_n20662_ = ~new_n20211_ & new_n20661_;
  assign new_n20663_ = ~new_n20215_ & ~new_n20662_;
  assign new_n20664_ = ~new_n20660_ & new_n20663_;
  assign new_n20665_ = ~new_n20215_ & ~new_n20664_;
  assign new_n20666_ = \b[34]  & ~new_n20204_;
  assign new_n20667_ = ~new_n20202_ & new_n20666_;
  assign new_n20668_ = ~new_n20206_ & ~new_n20667_;
  assign new_n20669_ = ~new_n20665_ & new_n20668_;
  assign new_n20670_ = ~new_n20206_ & ~new_n20669_;
  assign new_n20671_ = \b[35]  & ~new_n20195_;
  assign new_n20672_ = ~new_n20193_ & new_n20671_;
  assign new_n20673_ = ~new_n20197_ & ~new_n20672_;
  assign new_n20674_ = ~new_n20670_ & new_n20673_;
  assign new_n20675_ = ~new_n20197_ & ~new_n20674_;
  assign new_n20676_ = \b[36]  & ~new_n20186_;
  assign new_n20677_ = ~new_n20184_ & new_n20676_;
  assign new_n20678_ = ~new_n20188_ & ~new_n20677_;
  assign new_n20679_ = ~new_n20675_ & new_n20678_;
  assign new_n20680_ = ~new_n20188_ & ~new_n20679_;
  assign new_n20681_ = \b[37]  & ~new_n20177_;
  assign new_n20682_ = ~new_n20175_ & new_n20681_;
  assign new_n20683_ = ~new_n20179_ & ~new_n20682_;
  assign new_n20684_ = ~new_n20680_ & new_n20683_;
  assign new_n20685_ = ~new_n20179_ & ~new_n20684_;
  assign new_n20686_ = \b[38]  & ~new_n20168_;
  assign new_n20687_ = ~new_n20166_ & new_n20686_;
  assign new_n20688_ = ~new_n20170_ & ~new_n20687_;
  assign new_n20689_ = ~new_n20685_ & new_n20688_;
  assign new_n20690_ = ~new_n20170_ & ~new_n20689_;
  assign new_n20691_ = \b[39]  & ~new_n20159_;
  assign new_n20692_ = ~new_n20157_ & new_n20691_;
  assign new_n20693_ = ~new_n20161_ & ~new_n20692_;
  assign new_n20694_ = ~new_n20690_ & new_n20693_;
  assign new_n20695_ = ~new_n20161_ & ~new_n20694_;
  assign new_n20696_ = \b[40]  & ~new_n20150_;
  assign new_n20697_ = ~new_n20148_ & new_n20696_;
  assign new_n20698_ = ~new_n20152_ & ~new_n20697_;
  assign new_n20699_ = ~new_n20695_ & new_n20698_;
  assign new_n20700_ = ~new_n20152_ & ~new_n20699_;
  assign new_n20701_ = \b[41]  & ~new_n20141_;
  assign new_n20702_ = ~new_n20139_ & new_n20701_;
  assign new_n20703_ = ~new_n20143_ & ~new_n20702_;
  assign new_n20704_ = ~new_n20700_ & new_n20703_;
  assign new_n20705_ = ~new_n20143_ & ~new_n20704_;
  assign new_n20706_ = \b[42]  & ~new_n20132_;
  assign new_n20707_ = ~new_n20130_ & new_n20706_;
  assign new_n20708_ = ~new_n20134_ & ~new_n20707_;
  assign new_n20709_ = ~new_n20705_ & new_n20708_;
  assign new_n20710_ = ~new_n20134_ & ~new_n20709_;
  assign new_n20711_ = \b[43]  & ~new_n20123_;
  assign new_n20712_ = ~new_n20121_ & new_n20711_;
  assign new_n20713_ = ~new_n20125_ & ~new_n20712_;
  assign new_n20714_ = ~new_n20710_ & new_n20713_;
  assign new_n20715_ = ~new_n20125_ & ~new_n20714_;
  assign new_n20716_ = \b[44]  & ~new_n20114_;
  assign new_n20717_ = ~new_n20112_ & new_n20716_;
  assign new_n20718_ = ~new_n20116_ & ~new_n20717_;
  assign new_n20719_ = ~new_n20715_ & new_n20718_;
  assign new_n20720_ = ~new_n20116_ & ~new_n20719_;
  assign new_n20721_ = \b[45]  & ~new_n20105_;
  assign new_n20722_ = ~new_n20103_ & new_n20721_;
  assign new_n20723_ = ~new_n20107_ & ~new_n20722_;
  assign new_n20724_ = ~new_n20720_ & new_n20723_;
  assign new_n20725_ = ~new_n20107_ & ~new_n20724_;
  assign new_n20726_ = \b[46]  & ~new_n20096_;
  assign new_n20727_ = ~new_n20094_ & new_n20726_;
  assign new_n20728_ = ~new_n20098_ & ~new_n20727_;
  assign new_n20729_ = ~new_n20725_ & new_n20728_;
  assign new_n20730_ = ~new_n20098_ & ~new_n20729_;
  assign new_n20731_ = \b[47]  & ~new_n20087_;
  assign new_n20732_ = ~new_n20085_ & new_n20731_;
  assign new_n20733_ = ~new_n20089_ & ~new_n20732_;
  assign new_n20734_ = ~new_n20730_ & new_n20733_;
  assign new_n20735_ = ~new_n20089_ & ~new_n20734_;
  assign new_n20736_ = \b[48]  & ~new_n20078_;
  assign new_n20737_ = ~new_n20076_ & new_n20736_;
  assign new_n20738_ = ~new_n20080_ & ~new_n20737_;
  assign new_n20739_ = ~new_n20735_ & new_n20738_;
  assign new_n20740_ = ~new_n20080_ & ~new_n20739_;
  assign new_n20741_ = \b[49]  & ~new_n20069_;
  assign new_n20742_ = ~new_n20067_ & new_n20741_;
  assign new_n20743_ = ~new_n20071_ & ~new_n20742_;
  assign new_n20744_ = ~new_n20740_ & new_n20743_;
  assign new_n20745_ = ~new_n20071_ & ~new_n20744_;
  assign new_n20746_ = \b[50]  & ~new_n20060_;
  assign new_n20747_ = ~new_n20058_ & new_n20746_;
  assign new_n20748_ = ~new_n20062_ & ~new_n20747_;
  assign new_n20749_ = ~new_n20745_ & new_n20748_;
  assign new_n20750_ = ~new_n20062_ & ~new_n20749_;
  assign new_n20751_ = \b[51]  & ~new_n20051_;
  assign new_n20752_ = ~new_n20049_ & new_n20751_;
  assign new_n20753_ = ~new_n20053_ & ~new_n20752_;
  assign new_n20754_ = ~new_n20750_ & new_n20753_;
  assign new_n20755_ = ~new_n20053_ & ~new_n20754_;
  assign new_n20756_ = \b[52]  & ~new_n20042_;
  assign new_n20757_ = ~new_n20040_ & new_n20756_;
  assign new_n20758_ = ~new_n20044_ & ~new_n20757_;
  assign new_n20759_ = ~new_n20755_ & new_n20758_;
  assign new_n20760_ = ~new_n20044_ & ~new_n20759_;
  assign new_n20761_ = ~new_n19313_ & ~new_n20030_;
  assign new_n20762_ = ~new_n20028_ & new_n20761_;
  assign new_n20763_ = ~new_n20019_ & new_n20762_;
  assign new_n20764_ = ~new_n20028_ & ~new_n20030_;
  assign new_n20765_ = ~new_n20020_ & ~new_n20764_;
  assign new_n20766_ = ~new_n20763_ & ~new_n20765_;
  assign new_n20767_ = \quotient[11]  & ~new_n20766_;
  assign new_n20768_ = ~new_n20027_ & ~new_n20034_;
  assign new_n20769_ = ~new_n20033_ & new_n20768_;
  assign new_n20770_ = ~new_n20767_ & ~new_n20769_;
  assign new_n20771_ = ~\b[53]  & ~new_n20770_;
  assign new_n20772_ = \b[53]  & ~new_n20769_;
  assign new_n20773_ = ~new_n20767_ & new_n20772_;
  assign new_n20774_ = new_n283_ & new_n285_;
  assign new_n20775_ = new_n280_ & new_n20774_;
  assign new_n20776_ = ~new_n20773_ & new_n20775_;
  assign new_n20777_ = ~new_n20771_ & new_n20776_;
  assign new_n20778_ = ~new_n20760_ & new_n20777_;
  assign new_n20779_ = new_n595_ & ~new_n20770_;
  assign \quotient[10]  = new_n20778_ | new_n20779_;
  assign new_n20781_ = ~new_n20053_ & new_n20758_;
  assign new_n20782_ = ~new_n20754_ & new_n20781_;
  assign new_n20783_ = ~new_n20755_ & ~new_n20758_;
  assign new_n20784_ = ~new_n20782_ & ~new_n20783_;
  assign new_n20785_ = \quotient[10]  & ~new_n20784_;
  assign new_n20786_ = ~new_n20043_ & ~new_n20779_;
  assign new_n20787_ = ~new_n20778_ & new_n20786_;
  assign new_n20788_ = ~new_n20785_ & ~new_n20787_;
  assign new_n20789_ = ~new_n20044_ & ~new_n20773_;
  assign new_n20790_ = ~new_n20771_ & new_n20789_;
  assign new_n20791_ = ~new_n20759_ & new_n20790_;
  assign new_n20792_ = ~new_n20771_ & ~new_n20773_;
  assign new_n20793_ = ~new_n20760_ & ~new_n20792_;
  assign new_n20794_ = ~new_n20791_ & ~new_n20793_;
  assign new_n20795_ = \quotient[10]  & ~new_n20794_;
  assign new_n20796_ = ~new_n20770_ & ~new_n20779_;
  assign new_n20797_ = ~new_n20778_ & new_n20796_;
  assign new_n20798_ = ~new_n20795_ & ~new_n20797_;
  assign new_n20799_ = ~\b[54]  & ~new_n20798_;
  assign new_n20800_ = ~\b[53]  & ~new_n20788_;
  assign new_n20801_ = ~new_n20062_ & new_n20753_;
  assign new_n20802_ = ~new_n20749_ & new_n20801_;
  assign new_n20803_ = ~new_n20750_ & ~new_n20753_;
  assign new_n20804_ = ~new_n20802_ & ~new_n20803_;
  assign new_n20805_ = \quotient[10]  & ~new_n20804_;
  assign new_n20806_ = ~new_n20052_ & ~new_n20779_;
  assign new_n20807_ = ~new_n20778_ & new_n20806_;
  assign new_n20808_ = ~new_n20805_ & ~new_n20807_;
  assign new_n20809_ = ~\b[52]  & ~new_n20808_;
  assign new_n20810_ = ~new_n20071_ & new_n20748_;
  assign new_n20811_ = ~new_n20744_ & new_n20810_;
  assign new_n20812_ = ~new_n20745_ & ~new_n20748_;
  assign new_n20813_ = ~new_n20811_ & ~new_n20812_;
  assign new_n20814_ = \quotient[10]  & ~new_n20813_;
  assign new_n20815_ = ~new_n20061_ & ~new_n20779_;
  assign new_n20816_ = ~new_n20778_ & new_n20815_;
  assign new_n20817_ = ~new_n20814_ & ~new_n20816_;
  assign new_n20818_ = ~\b[51]  & ~new_n20817_;
  assign new_n20819_ = ~new_n20080_ & new_n20743_;
  assign new_n20820_ = ~new_n20739_ & new_n20819_;
  assign new_n20821_ = ~new_n20740_ & ~new_n20743_;
  assign new_n20822_ = ~new_n20820_ & ~new_n20821_;
  assign new_n20823_ = \quotient[10]  & ~new_n20822_;
  assign new_n20824_ = ~new_n20070_ & ~new_n20779_;
  assign new_n20825_ = ~new_n20778_ & new_n20824_;
  assign new_n20826_ = ~new_n20823_ & ~new_n20825_;
  assign new_n20827_ = ~\b[50]  & ~new_n20826_;
  assign new_n20828_ = ~new_n20089_ & new_n20738_;
  assign new_n20829_ = ~new_n20734_ & new_n20828_;
  assign new_n20830_ = ~new_n20735_ & ~new_n20738_;
  assign new_n20831_ = ~new_n20829_ & ~new_n20830_;
  assign new_n20832_ = \quotient[10]  & ~new_n20831_;
  assign new_n20833_ = ~new_n20079_ & ~new_n20779_;
  assign new_n20834_ = ~new_n20778_ & new_n20833_;
  assign new_n20835_ = ~new_n20832_ & ~new_n20834_;
  assign new_n20836_ = ~\b[49]  & ~new_n20835_;
  assign new_n20837_ = ~new_n20098_ & new_n20733_;
  assign new_n20838_ = ~new_n20729_ & new_n20837_;
  assign new_n20839_ = ~new_n20730_ & ~new_n20733_;
  assign new_n20840_ = ~new_n20838_ & ~new_n20839_;
  assign new_n20841_ = \quotient[10]  & ~new_n20840_;
  assign new_n20842_ = ~new_n20088_ & ~new_n20779_;
  assign new_n20843_ = ~new_n20778_ & new_n20842_;
  assign new_n20844_ = ~new_n20841_ & ~new_n20843_;
  assign new_n20845_ = ~\b[48]  & ~new_n20844_;
  assign new_n20846_ = ~new_n20107_ & new_n20728_;
  assign new_n20847_ = ~new_n20724_ & new_n20846_;
  assign new_n20848_ = ~new_n20725_ & ~new_n20728_;
  assign new_n20849_ = ~new_n20847_ & ~new_n20848_;
  assign new_n20850_ = \quotient[10]  & ~new_n20849_;
  assign new_n20851_ = ~new_n20097_ & ~new_n20779_;
  assign new_n20852_ = ~new_n20778_ & new_n20851_;
  assign new_n20853_ = ~new_n20850_ & ~new_n20852_;
  assign new_n20854_ = ~\b[47]  & ~new_n20853_;
  assign new_n20855_ = ~new_n20116_ & new_n20723_;
  assign new_n20856_ = ~new_n20719_ & new_n20855_;
  assign new_n20857_ = ~new_n20720_ & ~new_n20723_;
  assign new_n20858_ = ~new_n20856_ & ~new_n20857_;
  assign new_n20859_ = \quotient[10]  & ~new_n20858_;
  assign new_n20860_ = ~new_n20106_ & ~new_n20779_;
  assign new_n20861_ = ~new_n20778_ & new_n20860_;
  assign new_n20862_ = ~new_n20859_ & ~new_n20861_;
  assign new_n20863_ = ~\b[46]  & ~new_n20862_;
  assign new_n20864_ = ~new_n20125_ & new_n20718_;
  assign new_n20865_ = ~new_n20714_ & new_n20864_;
  assign new_n20866_ = ~new_n20715_ & ~new_n20718_;
  assign new_n20867_ = ~new_n20865_ & ~new_n20866_;
  assign new_n20868_ = \quotient[10]  & ~new_n20867_;
  assign new_n20869_ = ~new_n20115_ & ~new_n20779_;
  assign new_n20870_ = ~new_n20778_ & new_n20869_;
  assign new_n20871_ = ~new_n20868_ & ~new_n20870_;
  assign new_n20872_ = ~\b[45]  & ~new_n20871_;
  assign new_n20873_ = ~new_n20134_ & new_n20713_;
  assign new_n20874_ = ~new_n20709_ & new_n20873_;
  assign new_n20875_ = ~new_n20710_ & ~new_n20713_;
  assign new_n20876_ = ~new_n20874_ & ~new_n20875_;
  assign new_n20877_ = \quotient[10]  & ~new_n20876_;
  assign new_n20878_ = ~new_n20124_ & ~new_n20779_;
  assign new_n20879_ = ~new_n20778_ & new_n20878_;
  assign new_n20880_ = ~new_n20877_ & ~new_n20879_;
  assign new_n20881_ = ~\b[44]  & ~new_n20880_;
  assign new_n20882_ = ~new_n20143_ & new_n20708_;
  assign new_n20883_ = ~new_n20704_ & new_n20882_;
  assign new_n20884_ = ~new_n20705_ & ~new_n20708_;
  assign new_n20885_ = ~new_n20883_ & ~new_n20884_;
  assign new_n20886_ = \quotient[10]  & ~new_n20885_;
  assign new_n20887_ = ~new_n20133_ & ~new_n20779_;
  assign new_n20888_ = ~new_n20778_ & new_n20887_;
  assign new_n20889_ = ~new_n20886_ & ~new_n20888_;
  assign new_n20890_ = ~\b[43]  & ~new_n20889_;
  assign new_n20891_ = ~new_n20152_ & new_n20703_;
  assign new_n20892_ = ~new_n20699_ & new_n20891_;
  assign new_n20893_ = ~new_n20700_ & ~new_n20703_;
  assign new_n20894_ = ~new_n20892_ & ~new_n20893_;
  assign new_n20895_ = \quotient[10]  & ~new_n20894_;
  assign new_n20896_ = ~new_n20142_ & ~new_n20779_;
  assign new_n20897_ = ~new_n20778_ & new_n20896_;
  assign new_n20898_ = ~new_n20895_ & ~new_n20897_;
  assign new_n20899_ = ~\b[42]  & ~new_n20898_;
  assign new_n20900_ = ~new_n20161_ & new_n20698_;
  assign new_n20901_ = ~new_n20694_ & new_n20900_;
  assign new_n20902_ = ~new_n20695_ & ~new_n20698_;
  assign new_n20903_ = ~new_n20901_ & ~new_n20902_;
  assign new_n20904_ = \quotient[10]  & ~new_n20903_;
  assign new_n20905_ = ~new_n20151_ & ~new_n20779_;
  assign new_n20906_ = ~new_n20778_ & new_n20905_;
  assign new_n20907_ = ~new_n20904_ & ~new_n20906_;
  assign new_n20908_ = ~\b[41]  & ~new_n20907_;
  assign new_n20909_ = ~new_n20170_ & new_n20693_;
  assign new_n20910_ = ~new_n20689_ & new_n20909_;
  assign new_n20911_ = ~new_n20690_ & ~new_n20693_;
  assign new_n20912_ = ~new_n20910_ & ~new_n20911_;
  assign new_n20913_ = \quotient[10]  & ~new_n20912_;
  assign new_n20914_ = ~new_n20160_ & ~new_n20779_;
  assign new_n20915_ = ~new_n20778_ & new_n20914_;
  assign new_n20916_ = ~new_n20913_ & ~new_n20915_;
  assign new_n20917_ = ~\b[40]  & ~new_n20916_;
  assign new_n20918_ = ~new_n20179_ & new_n20688_;
  assign new_n20919_ = ~new_n20684_ & new_n20918_;
  assign new_n20920_ = ~new_n20685_ & ~new_n20688_;
  assign new_n20921_ = ~new_n20919_ & ~new_n20920_;
  assign new_n20922_ = \quotient[10]  & ~new_n20921_;
  assign new_n20923_ = ~new_n20169_ & ~new_n20779_;
  assign new_n20924_ = ~new_n20778_ & new_n20923_;
  assign new_n20925_ = ~new_n20922_ & ~new_n20924_;
  assign new_n20926_ = ~\b[39]  & ~new_n20925_;
  assign new_n20927_ = ~new_n20188_ & new_n20683_;
  assign new_n20928_ = ~new_n20679_ & new_n20927_;
  assign new_n20929_ = ~new_n20680_ & ~new_n20683_;
  assign new_n20930_ = ~new_n20928_ & ~new_n20929_;
  assign new_n20931_ = \quotient[10]  & ~new_n20930_;
  assign new_n20932_ = ~new_n20178_ & ~new_n20779_;
  assign new_n20933_ = ~new_n20778_ & new_n20932_;
  assign new_n20934_ = ~new_n20931_ & ~new_n20933_;
  assign new_n20935_ = ~\b[38]  & ~new_n20934_;
  assign new_n20936_ = ~new_n20197_ & new_n20678_;
  assign new_n20937_ = ~new_n20674_ & new_n20936_;
  assign new_n20938_ = ~new_n20675_ & ~new_n20678_;
  assign new_n20939_ = ~new_n20937_ & ~new_n20938_;
  assign new_n20940_ = \quotient[10]  & ~new_n20939_;
  assign new_n20941_ = ~new_n20187_ & ~new_n20779_;
  assign new_n20942_ = ~new_n20778_ & new_n20941_;
  assign new_n20943_ = ~new_n20940_ & ~new_n20942_;
  assign new_n20944_ = ~\b[37]  & ~new_n20943_;
  assign new_n20945_ = ~new_n20206_ & new_n20673_;
  assign new_n20946_ = ~new_n20669_ & new_n20945_;
  assign new_n20947_ = ~new_n20670_ & ~new_n20673_;
  assign new_n20948_ = ~new_n20946_ & ~new_n20947_;
  assign new_n20949_ = \quotient[10]  & ~new_n20948_;
  assign new_n20950_ = ~new_n20196_ & ~new_n20779_;
  assign new_n20951_ = ~new_n20778_ & new_n20950_;
  assign new_n20952_ = ~new_n20949_ & ~new_n20951_;
  assign new_n20953_ = ~\b[36]  & ~new_n20952_;
  assign new_n20954_ = ~new_n20215_ & new_n20668_;
  assign new_n20955_ = ~new_n20664_ & new_n20954_;
  assign new_n20956_ = ~new_n20665_ & ~new_n20668_;
  assign new_n20957_ = ~new_n20955_ & ~new_n20956_;
  assign new_n20958_ = \quotient[10]  & ~new_n20957_;
  assign new_n20959_ = ~new_n20205_ & ~new_n20779_;
  assign new_n20960_ = ~new_n20778_ & new_n20959_;
  assign new_n20961_ = ~new_n20958_ & ~new_n20960_;
  assign new_n20962_ = ~\b[35]  & ~new_n20961_;
  assign new_n20963_ = ~new_n20224_ & new_n20663_;
  assign new_n20964_ = ~new_n20659_ & new_n20963_;
  assign new_n20965_ = ~new_n20660_ & ~new_n20663_;
  assign new_n20966_ = ~new_n20964_ & ~new_n20965_;
  assign new_n20967_ = \quotient[10]  & ~new_n20966_;
  assign new_n20968_ = ~new_n20214_ & ~new_n20779_;
  assign new_n20969_ = ~new_n20778_ & new_n20968_;
  assign new_n20970_ = ~new_n20967_ & ~new_n20969_;
  assign new_n20971_ = ~\b[34]  & ~new_n20970_;
  assign new_n20972_ = ~new_n20233_ & new_n20658_;
  assign new_n20973_ = ~new_n20654_ & new_n20972_;
  assign new_n20974_ = ~new_n20655_ & ~new_n20658_;
  assign new_n20975_ = ~new_n20973_ & ~new_n20974_;
  assign new_n20976_ = \quotient[10]  & ~new_n20975_;
  assign new_n20977_ = ~new_n20223_ & ~new_n20779_;
  assign new_n20978_ = ~new_n20778_ & new_n20977_;
  assign new_n20979_ = ~new_n20976_ & ~new_n20978_;
  assign new_n20980_ = ~\b[33]  & ~new_n20979_;
  assign new_n20981_ = ~new_n20242_ & new_n20653_;
  assign new_n20982_ = ~new_n20649_ & new_n20981_;
  assign new_n20983_ = ~new_n20650_ & ~new_n20653_;
  assign new_n20984_ = ~new_n20982_ & ~new_n20983_;
  assign new_n20985_ = \quotient[10]  & ~new_n20984_;
  assign new_n20986_ = ~new_n20232_ & ~new_n20779_;
  assign new_n20987_ = ~new_n20778_ & new_n20986_;
  assign new_n20988_ = ~new_n20985_ & ~new_n20987_;
  assign new_n20989_ = ~\b[32]  & ~new_n20988_;
  assign new_n20990_ = ~new_n20251_ & new_n20648_;
  assign new_n20991_ = ~new_n20644_ & new_n20990_;
  assign new_n20992_ = ~new_n20645_ & ~new_n20648_;
  assign new_n20993_ = ~new_n20991_ & ~new_n20992_;
  assign new_n20994_ = \quotient[10]  & ~new_n20993_;
  assign new_n20995_ = ~new_n20241_ & ~new_n20779_;
  assign new_n20996_ = ~new_n20778_ & new_n20995_;
  assign new_n20997_ = ~new_n20994_ & ~new_n20996_;
  assign new_n20998_ = ~\b[31]  & ~new_n20997_;
  assign new_n20999_ = ~new_n20260_ & new_n20643_;
  assign new_n21000_ = ~new_n20639_ & new_n20999_;
  assign new_n21001_ = ~new_n20640_ & ~new_n20643_;
  assign new_n21002_ = ~new_n21000_ & ~new_n21001_;
  assign new_n21003_ = \quotient[10]  & ~new_n21002_;
  assign new_n21004_ = ~new_n20250_ & ~new_n20779_;
  assign new_n21005_ = ~new_n20778_ & new_n21004_;
  assign new_n21006_ = ~new_n21003_ & ~new_n21005_;
  assign new_n21007_ = ~\b[30]  & ~new_n21006_;
  assign new_n21008_ = ~new_n20269_ & new_n20638_;
  assign new_n21009_ = ~new_n20634_ & new_n21008_;
  assign new_n21010_ = ~new_n20635_ & ~new_n20638_;
  assign new_n21011_ = ~new_n21009_ & ~new_n21010_;
  assign new_n21012_ = \quotient[10]  & ~new_n21011_;
  assign new_n21013_ = ~new_n20259_ & ~new_n20779_;
  assign new_n21014_ = ~new_n20778_ & new_n21013_;
  assign new_n21015_ = ~new_n21012_ & ~new_n21014_;
  assign new_n21016_ = ~\b[29]  & ~new_n21015_;
  assign new_n21017_ = ~new_n20278_ & new_n20633_;
  assign new_n21018_ = ~new_n20629_ & new_n21017_;
  assign new_n21019_ = ~new_n20630_ & ~new_n20633_;
  assign new_n21020_ = ~new_n21018_ & ~new_n21019_;
  assign new_n21021_ = \quotient[10]  & ~new_n21020_;
  assign new_n21022_ = ~new_n20268_ & ~new_n20779_;
  assign new_n21023_ = ~new_n20778_ & new_n21022_;
  assign new_n21024_ = ~new_n21021_ & ~new_n21023_;
  assign new_n21025_ = ~\b[28]  & ~new_n21024_;
  assign new_n21026_ = ~new_n20287_ & new_n20628_;
  assign new_n21027_ = ~new_n20624_ & new_n21026_;
  assign new_n21028_ = ~new_n20625_ & ~new_n20628_;
  assign new_n21029_ = ~new_n21027_ & ~new_n21028_;
  assign new_n21030_ = \quotient[10]  & ~new_n21029_;
  assign new_n21031_ = ~new_n20277_ & ~new_n20779_;
  assign new_n21032_ = ~new_n20778_ & new_n21031_;
  assign new_n21033_ = ~new_n21030_ & ~new_n21032_;
  assign new_n21034_ = ~\b[27]  & ~new_n21033_;
  assign new_n21035_ = ~new_n20296_ & new_n20623_;
  assign new_n21036_ = ~new_n20619_ & new_n21035_;
  assign new_n21037_ = ~new_n20620_ & ~new_n20623_;
  assign new_n21038_ = ~new_n21036_ & ~new_n21037_;
  assign new_n21039_ = \quotient[10]  & ~new_n21038_;
  assign new_n21040_ = ~new_n20286_ & ~new_n20779_;
  assign new_n21041_ = ~new_n20778_ & new_n21040_;
  assign new_n21042_ = ~new_n21039_ & ~new_n21041_;
  assign new_n21043_ = ~\b[26]  & ~new_n21042_;
  assign new_n21044_ = ~new_n20305_ & new_n20618_;
  assign new_n21045_ = ~new_n20614_ & new_n21044_;
  assign new_n21046_ = ~new_n20615_ & ~new_n20618_;
  assign new_n21047_ = ~new_n21045_ & ~new_n21046_;
  assign new_n21048_ = \quotient[10]  & ~new_n21047_;
  assign new_n21049_ = ~new_n20295_ & ~new_n20779_;
  assign new_n21050_ = ~new_n20778_ & new_n21049_;
  assign new_n21051_ = ~new_n21048_ & ~new_n21050_;
  assign new_n21052_ = ~\b[25]  & ~new_n21051_;
  assign new_n21053_ = ~new_n20314_ & new_n20613_;
  assign new_n21054_ = ~new_n20609_ & new_n21053_;
  assign new_n21055_ = ~new_n20610_ & ~new_n20613_;
  assign new_n21056_ = ~new_n21054_ & ~new_n21055_;
  assign new_n21057_ = \quotient[10]  & ~new_n21056_;
  assign new_n21058_ = ~new_n20304_ & ~new_n20779_;
  assign new_n21059_ = ~new_n20778_ & new_n21058_;
  assign new_n21060_ = ~new_n21057_ & ~new_n21059_;
  assign new_n21061_ = ~\b[24]  & ~new_n21060_;
  assign new_n21062_ = ~new_n20323_ & new_n20608_;
  assign new_n21063_ = ~new_n20604_ & new_n21062_;
  assign new_n21064_ = ~new_n20605_ & ~new_n20608_;
  assign new_n21065_ = ~new_n21063_ & ~new_n21064_;
  assign new_n21066_ = \quotient[10]  & ~new_n21065_;
  assign new_n21067_ = ~new_n20313_ & ~new_n20779_;
  assign new_n21068_ = ~new_n20778_ & new_n21067_;
  assign new_n21069_ = ~new_n21066_ & ~new_n21068_;
  assign new_n21070_ = ~\b[23]  & ~new_n21069_;
  assign new_n21071_ = ~new_n20332_ & new_n20603_;
  assign new_n21072_ = ~new_n20599_ & new_n21071_;
  assign new_n21073_ = ~new_n20600_ & ~new_n20603_;
  assign new_n21074_ = ~new_n21072_ & ~new_n21073_;
  assign new_n21075_ = \quotient[10]  & ~new_n21074_;
  assign new_n21076_ = ~new_n20322_ & ~new_n20779_;
  assign new_n21077_ = ~new_n20778_ & new_n21076_;
  assign new_n21078_ = ~new_n21075_ & ~new_n21077_;
  assign new_n21079_ = ~\b[22]  & ~new_n21078_;
  assign new_n21080_ = ~new_n20341_ & new_n20598_;
  assign new_n21081_ = ~new_n20594_ & new_n21080_;
  assign new_n21082_ = ~new_n20595_ & ~new_n20598_;
  assign new_n21083_ = ~new_n21081_ & ~new_n21082_;
  assign new_n21084_ = \quotient[10]  & ~new_n21083_;
  assign new_n21085_ = ~new_n20331_ & ~new_n20779_;
  assign new_n21086_ = ~new_n20778_ & new_n21085_;
  assign new_n21087_ = ~new_n21084_ & ~new_n21086_;
  assign new_n21088_ = ~\b[21]  & ~new_n21087_;
  assign new_n21089_ = ~new_n20350_ & new_n20593_;
  assign new_n21090_ = ~new_n20589_ & new_n21089_;
  assign new_n21091_ = ~new_n20590_ & ~new_n20593_;
  assign new_n21092_ = ~new_n21090_ & ~new_n21091_;
  assign new_n21093_ = \quotient[10]  & ~new_n21092_;
  assign new_n21094_ = ~new_n20340_ & ~new_n20779_;
  assign new_n21095_ = ~new_n20778_ & new_n21094_;
  assign new_n21096_ = ~new_n21093_ & ~new_n21095_;
  assign new_n21097_ = ~\b[20]  & ~new_n21096_;
  assign new_n21098_ = ~new_n20359_ & new_n20588_;
  assign new_n21099_ = ~new_n20584_ & new_n21098_;
  assign new_n21100_ = ~new_n20585_ & ~new_n20588_;
  assign new_n21101_ = ~new_n21099_ & ~new_n21100_;
  assign new_n21102_ = \quotient[10]  & ~new_n21101_;
  assign new_n21103_ = ~new_n20349_ & ~new_n20779_;
  assign new_n21104_ = ~new_n20778_ & new_n21103_;
  assign new_n21105_ = ~new_n21102_ & ~new_n21104_;
  assign new_n21106_ = ~\b[19]  & ~new_n21105_;
  assign new_n21107_ = ~new_n20368_ & new_n20583_;
  assign new_n21108_ = ~new_n20579_ & new_n21107_;
  assign new_n21109_ = ~new_n20580_ & ~new_n20583_;
  assign new_n21110_ = ~new_n21108_ & ~new_n21109_;
  assign new_n21111_ = \quotient[10]  & ~new_n21110_;
  assign new_n21112_ = ~new_n20358_ & ~new_n20779_;
  assign new_n21113_ = ~new_n20778_ & new_n21112_;
  assign new_n21114_ = ~new_n21111_ & ~new_n21113_;
  assign new_n21115_ = ~\b[18]  & ~new_n21114_;
  assign new_n21116_ = ~new_n20377_ & new_n20578_;
  assign new_n21117_ = ~new_n20574_ & new_n21116_;
  assign new_n21118_ = ~new_n20575_ & ~new_n20578_;
  assign new_n21119_ = ~new_n21117_ & ~new_n21118_;
  assign new_n21120_ = \quotient[10]  & ~new_n21119_;
  assign new_n21121_ = ~new_n20367_ & ~new_n20779_;
  assign new_n21122_ = ~new_n20778_ & new_n21121_;
  assign new_n21123_ = ~new_n21120_ & ~new_n21122_;
  assign new_n21124_ = ~\b[17]  & ~new_n21123_;
  assign new_n21125_ = ~new_n20386_ & new_n20573_;
  assign new_n21126_ = ~new_n20569_ & new_n21125_;
  assign new_n21127_ = ~new_n20570_ & ~new_n20573_;
  assign new_n21128_ = ~new_n21126_ & ~new_n21127_;
  assign new_n21129_ = \quotient[10]  & ~new_n21128_;
  assign new_n21130_ = ~new_n20376_ & ~new_n20779_;
  assign new_n21131_ = ~new_n20778_ & new_n21130_;
  assign new_n21132_ = ~new_n21129_ & ~new_n21131_;
  assign new_n21133_ = ~\b[16]  & ~new_n21132_;
  assign new_n21134_ = ~new_n20395_ & new_n20568_;
  assign new_n21135_ = ~new_n20564_ & new_n21134_;
  assign new_n21136_ = ~new_n20565_ & ~new_n20568_;
  assign new_n21137_ = ~new_n21135_ & ~new_n21136_;
  assign new_n21138_ = \quotient[10]  & ~new_n21137_;
  assign new_n21139_ = ~new_n20385_ & ~new_n20779_;
  assign new_n21140_ = ~new_n20778_ & new_n21139_;
  assign new_n21141_ = ~new_n21138_ & ~new_n21140_;
  assign new_n21142_ = ~\b[15]  & ~new_n21141_;
  assign new_n21143_ = ~new_n20404_ & new_n20563_;
  assign new_n21144_ = ~new_n20559_ & new_n21143_;
  assign new_n21145_ = ~new_n20560_ & ~new_n20563_;
  assign new_n21146_ = ~new_n21144_ & ~new_n21145_;
  assign new_n21147_ = \quotient[10]  & ~new_n21146_;
  assign new_n21148_ = ~new_n20394_ & ~new_n20779_;
  assign new_n21149_ = ~new_n20778_ & new_n21148_;
  assign new_n21150_ = ~new_n21147_ & ~new_n21149_;
  assign new_n21151_ = ~\b[14]  & ~new_n21150_;
  assign new_n21152_ = ~new_n20413_ & new_n20558_;
  assign new_n21153_ = ~new_n20554_ & new_n21152_;
  assign new_n21154_ = ~new_n20555_ & ~new_n20558_;
  assign new_n21155_ = ~new_n21153_ & ~new_n21154_;
  assign new_n21156_ = \quotient[10]  & ~new_n21155_;
  assign new_n21157_ = ~new_n20403_ & ~new_n20779_;
  assign new_n21158_ = ~new_n20778_ & new_n21157_;
  assign new_n21159_ = ~new_n21156_ & ~new_n21158_;
  assign new_n21160_ = ~\b[13]  & ~new_n21159_;
  assign new_n21161_ = ~new_n20422_ & new_n20553_;
  assign new_n21162_ = ~new_n20549_ & new_n21161_;
  assign new_n21163_ = ~new_n20550_ & ~new_n20553_;
  assign new_n21164_ = ~new_n21162_ & ~new_n21163_;
  assign new_n21165_ = \quotient[10]  & ~new_n21164_;
  assign new_n21166_ = ~new_n20412_ & ~new_n20779_;
  assign new_n21167_ = ~new_n20778_ & new_n21166_;
  assign new_n21168_ = ~new_n21165_ & ~new_n21167_;
  assign new_n21169_ = ~\b[12]  & ~new_n21168_;
  assign new_n21170_ = ~new_n20431_ & new_n20548_;
  assign new_n21171_ = ~new_n20544_ & new_n21170_;
  assign new_n21172_ = ~new_n20545_ & ~new_n20548_;
  assign new_n21173_ = ~new_n21171_ & ~new_n21172_;
  assign new_n21174_ = \quotient[10]  & ~new_n21173_;
  assign new_n21175_ = ~new_n20421_ & ~new_n20779_;
  assign new_n21176_ = ~new_n20778_ & new_n21175_;
  assign new_n21177_ = ~new_n21174_ & ~new_n21176_;
  assign new_n21178_ = ~\b[11]  & ~new_n21177_;
  assign new_n21179_ = ~new_n20440_ & new_n20543_;
  assign new_n21180_ = ~new_n20539_ & new_n21179_;
  assign new_n21181_ = ~new_n20540_ & ~new_n20543_;
  assign new_n21182_ = ~new_n21180_ & ~new_n21181_;
  assign new_n21183_ = \quotient[10]  & ~new_n21182_;
  assign new_n21184_ = ~new_n20430_ & ~new_n20779_;
  assign new_n21185_ = ~new_n20778_ & new_n21184_;
  assign new_n21186_ = ~new_n21183_ & ~new_n21185_;
  assign new_n21187_ = ~\b[10]  & ~new_n21186_;
  assign new_n21188_ = ~new_n20449_ & new_n20538_;
  assign new_n21189_ = ~new_n20534_ & new_n21188_;
  assign new_n21190_ = ~new_n20535_ & ~new_n20538_;
  assign new_n21191_ = ~new_n21189_ & ~new_n21190_;
  assign new_n21192_ = \quotient[10]  & ~new_n21191_;
  assign new_n21193_ = ~new_n20439_ & ~new_n20779_;
  assign new_n21194_ = ~new_n20778_ & new_n21193_;
  assign new_n21195_ = ~new_n21192_ & ~new_n21194_;
  assign new_n21196_ = ~\b[9]  & ~new_n21195_;
  assign new_n21197_ = ~new_n20458_ & new_n20533_;
  assign new_n21198_ = ~new_n20529_ & new_n21197_;
  assign new_n21199_ = ~new_n20530_ & ~new_n20533_;
  assign new_n21200_ = ~new_n21198_ & ~new_n21199_;
  assign new_n21201_ = \quotient[10]  & ~new_n21200_;
  assign new_n21202_ = ~new_n20448_ & ~new_n20779_;
  assign new_n21203_ = ~new_n20778_ & new_n21202_;
  assign new_n21204_ = ~new_n21201_ & ~new_n21203_;
  assign new_n21205_ = ~\b[8]  & ~new_n21204_;
  assign new_n21206_ = ~new_n20467_ & new_n20528_;
  assign new_n21207_ = ~new_n20524_ & new_n21206_;
  assign new_n21208_ = ~new_n20525_ & ~new_n20528_;
  assign new_n21209_ = ~new_n21207_ & ~new_n21208_;
  assign new_n21210_ = \quotient[10]  & ~new_n21209_;
  assign new_n21211_ = ~new_n20457_ & ~new_n20779_;
  assign new_n21212_ = ~new_n20778_ & new_n21211_;
  assign new_n21213_ = ~new_n21210_ & ~new_n21212_;
  assign new_n21214_ = ~\b[7]  & ~new_n21213_;
  assign new_n21215_ = ~new_n20476_ & new_n20523_;
  assign new_n21216_ = ~new_n20519_ & new_n21215_;
  assign new_n21217_ = ~new_n20520_ & ~new_n20523_;
  assign new_n21218_ = ~new_n21216_ & ~new_n21217_;
  assign new_n21219_ = \quotient[10]  & ~new_n21218_;
  assign new_n21220_ = ~new_n20466_ & ~new_n20779_;
  assign new_n21221_ = ~new_n20778_ & new_n21220_;
  assign new_n21222_ = ~new_n21219_ & ~new_n21221_;
  assign new_n21223_ = ~\b[6]  & ~new_n21222_;
  assign new_n21224_ = ~new_n20485_ & new_n20518_;
  assign new_n21225_ = ~new_n20514_ & new_n21224_;
  assign new_n21226_ = ~new_n20515_ & ~new_n20518_;
  assign new_n21227_ = ~new_n21225_ & ~new_n21226_;
  assign new_n21228_ = \quotient[10]  & ~new_n21227_;
  assign new_n21229_ = ~new_n20475_ & ~new_n20779_;
  assign new_n21230_ = ~new_n20778_ & new_n21229_;
  assign new_n21231_ = ~new_n21228_ & ~new_n21230_;
  assign new_n21232_ = ~\b[5]  & ~new_n21231_;
  assign new_n21233_ = ~new_n20493_ & new_n20513_;
  assign new_n21234_ = ~new_n20509_ & new_n21233_;
  assign new_n21235_ = ~new_n20510_ & ~new_n20513_;
  assign new_n21236_ = ~new_n21234_ & ~new_n21235_;
  assign new_n21237_ = \quotient[10]  & ~new_n21236_;
  assign new_n21238_ = ~new_n20484_ & ~new_n20779_;
  assign new_n21239_ = ~new_n20778_ & new_n21238_;
  assign new_n21240_ = ~new_n21237_ & ~new_n21239_;
  assign new_n21241_ = ~\b[4]  & ~new_n21240_;
  assign new_n21242_ = ~new_n20504_ & new_n20508_;
  assign new_n21243_ = ~new_n20503_ & new_n21242_;
  assign new_n21244_ = ~new_n20505_ & ~new_n20508_;
  assign new_n21245_ = ~new_n21243_ & ~new_n21244_;
  assign new_n21246_ = \quotient[10]  & ~new_n21245_;
  assign new_n21247_ = ~new_n20492_ & ~new_n20779_;
  assign new_n21248_ = ~new_n20778_ & new_n21247_;
  assign new_n21249_ = ~new_n21246_ & ~new_n21248_;
  assign new_n21250_ = ~\b[3]  & ~new_n21249_;
  assign new_n21251_ = ~new_n20500_ & new_n20502_;
  assign new_n21252_ = ~new_n20498_ & new_n21251_;
  assign new_n21253_ = ~new_n20503_ & ~new_n21252_;
  assign new_n21254_ = \quotient[10]  & new_n21253_;
  assign new_n21255_ = ~new_n20497_ & ~new_n20779_;
  assign new_n21256_ = ~new_n20778_ & new_n21255_;
  assign new_n21257_ = ~new_n21254_ & ~new_n21256_;
  assign new_n21258_ = ~\b[2]  & ~new_n21257_;
  assign new_n21259_ = \b[0]  & \quotient[10] ;
  assign new_n21260_ = \a[10]  & ~new_n21259_;
  assign new_n21261_ = new_n20502_ & \quotient[10] ;
  assign new_n21262_ = ~new_n21260_ & ~new_n21261_;
  assign new_n21263_ = \b[1]  & ~new_n21262_;
  assign new_n21264_ = ~\b[1]  & ~new_n21261_;
  assign new_n21265_ = ~new_n21260_ & new_n21264_;
  assign new_n21266_ = ~new_n21263_ & ~new_n21265_;
  assign new_n21267_ = ~\a[9]  & \b[0] ;
  assign new_n21268_ = ~new_n21266_ & ~new_n21267_;
  assign new_n21269_ = ~\b[1]  & ~new_n21262_;
  assign new_n21270_ = ~new_n21268_ & ~new_n21269_;
  assign new_n21271_ = \b[2]  & ~new_n21256_;
  assign new_n21272_ = ~new_n21254_ & new_n21271_;
  assign new_n21273_ = ~new_n21258_ & ~new_n21272_;
  assign new_n21274_ = ~new_n21270_ & new_n21273_;
  assign new_n21275_ = ~new_n21258_ & ~new_n21274_;
  assign new_n21276_ = \b[3]  & ~new_n21248_;
  assign new_n21277_ = ~new_n21246_ & new_n21276_;
  assign new_n21278_ = ~new_n21250_ & ~new_n21277_;
  assign new_n21279_ = ~new_n21275_ & new_n21278_;
  assign new_n21280_ = ~new_n21250_ & ~new_n21279_;
  assign new_n21281_ = \b[4]  & ~new_n21239_;
  assign new_n21282_ = ~new_n21237_ & new_n21281_;
  assign new_n21283_ = ~new_n21241_ & ~new_n21282_;
  assign new_n21284_ = ~new_n21280_ & new_n21283_;
  assign new_n21285_ = ~new_n21241_ & ~new_n21284_;
  assign new_n21286_ = \b[5]  & ~new_n21230_;
  assign new_n21287_ = ~new_n21228_ & new_n21286_;
  assign new_n21288_ = ~new_n21232_ & ~new_n21287_;
  assign new_n21289_ = ~new_n21285_ & new_n21288_;
  assign new_n21290_ = ~new_n21232_ & ~new_n21289_;
  assign new_n21291_ = \b[6]  & ~new_n21221_;
  assign new_n21292_ = ~new_n21219_ & new_n21291_;
  assign new_n21293_ = ~new_n21223_ & ~new_n21292_;
  assign new_n21294_ = ~new_n21290_ & new_n21293_;
  assign new_n21295_ = ~new_n21223_ & ~new_n21294_;
  assign new_n21296_ = \b[7]  & ~new_n21212_;
  assign new_n21297_ = ~new_n21210_ & new_n21296_;
  assign new_n21298_ = ~new_n21214_ & ~new_n21297_;
  assign new_n21299_ = ~new_n21295_ & new_n21298_;
  assign new_n21300_ = ~new_n21214_ & ~new_n21299_;
  assign new_n21301_ = \b[8]  & ~new_n21203_;
  assign new_n21302_ = ~new_n21201_ & new_n21301_;
  assign new_n21303_ = ~new_n21205_ & ~new_n21302_;
  assign new_n21304_ = ~new_n21300_ & new_n21303_;
  assign new_n21305_ = ~new_n21205_ & ~new_n21304_;
  assign new_n21306_ = \b[9]  & ~new_n21194_;
  assign new_n21307_ = ~new_n21192_ & new_n21306_;
  assign new_n21308_ = ~new_n21196_ & ~new_n21307_;
  assign new_n21309_ = ~new_n21305_ & new_n21308_;
  assign new_n21310_ = ~new_n21196_ & ~new_n21309_;
  assign new_n21311_ = \b[10]  & ~new_n21185_;
  assign new_n21312_ = ~new_n21183_ & new_n21311_;
  assign new_n21313_ = ~new_n21187_ & ~new_n21312_;
  assign new_n21314_ = ~new_n21310_ & new_n21313_;
  assign new_n21315_ = ~new_n21187_ & ~new_n21314_;
  assign new_n21316_ = \b[11]  & ~new_n21176_;
  assign new_n21317_ = ~new_n21174_ & new_n21316_;
  assign new_n21318_ = ~new_n21178_ & ~new_n21317_;
  assign new_n21319_ = ~new_n21315_ & new_n21318_;
  assign new_n21320_ = ~new_n21178_ & ~new_n21319_;
  assign new_n21321_ = \b[12]  & ~new_n21167_;
  assign new_n21322_ = ~new_n21165_ & new_n21321_;
  assign new_n21323_ = ~new_n21169_ & ~new_n21322_;
  assign new_n21324_ = ~new_n21320_ & new_n21323_;
  assign new_n21325_ = ~new_n21169_ & ~new_n21324_;
  assign new_n21326_ = \b[13]  & ~new_n21158_;
  assign new_n21327_ = ~new_n21156_ & new_n21326_;
  assign new_n21328_ = ~new_n21160_ & ~new_n21327_;
  assign new_n21329_ = ~new_n21325_ & new_n21328_;
  assign new_n21330_ = ~new_n21160_ & ~new_n21329_;
  assign new_n21331_ = \b[14]  & ~new_n21149_;
  assign new_n21332_ = ~new_n21147_ & new_n21331_;
  assign new_n21333_ = ~new_n21151_ & ~new_n21332_;
  assign new_n21334_ = ~new_n21330_ & new_n21333_;
  assign new_n21335_ = ~new_n21151_ & ~new_n21334_;
  assign new_n21336_ = \b[15]  & ~new_n21140_;
  assign new_n21337_ = ~new_n21138_ & new_n21336_;
  assign new_n21338_ = ~new_n21142_ & ~new_n21337_;
  assign new_n21339_ = ~new_n21335_ & new_n21338_;
  assign new_n21340_ = ~new_n21142_ & ~new_n21339_;
  assign new_n21341_ = \b[16]  & ~new_n21131_;
  assign new_n21342_ = ~new_n21129_ & new_n21341_;
  assign new_n21343_ = ~new_n21133_ & ~new_n21342_;
  assign new_n21344_ = ~new_n21340_ & new_n21343_;
  assign new_n21345_ = ~new_n21133_ & ~new_n21344_;
  assign new_n21346_ = \b[17]  & ~new_n21122_;
  assign new_n21347_ = ~new_n21120_ & new_n21346_;
  assign new_n21348_ = ~new_n21124_ & ~new_n21347_;
  assign new_n21349_ = ~new_n21345_ & new_n21348_;
  assign new_n21350_ = ~new_n21124_ & ~new_n21349_;
  assign new_n21351_ = \b[18]  & ~new_n21113_;
  assign new_n21352_ = ~new_n21111_ & new_n21351_;
  assign new_n21353_ = ~new_n21115_ & ~new_n21352_;
  assign new_n21354_ = ~new_n21350_ & new_n21353_;
  assign new_n21355_ = ~new_n21115_ & ~new_n21354_;
  assign new_n21356_ = \b[19]  & ~new_n21104_;
  assign new_n21357_ = ~new_n21102_ & new_n21356_;
  assign new_n21358_ = ~new_n21106_ & ~new_n21357_;
  assign new_n21359_ = ~new_n21355_ & new_n21358_;
  assign new_n21360_ = ~new_n21106_ & ~new_n21359_;
  assign new_n21361_ = \b[20]  & ~new_n21095_;
  assign new_n21362_ = ~new_n21093_ & new_n21361_;
  assign new_n21363_ = ~new_n21097_ & ~new_n21362_;
  assign new_n21364_ = ~new_n21360_ & new_n21363_;
  assign new_n21365_ = ~new_n21097_ & ~new_n21364_;
  assign new_n21366_ = \b[21]  & ~new_n21086_;
  assign new_n21367_ = ~new_n21084_ & new_n21366_;
  assign new_n21368_ = ~new_n21088_ & ~new_n21367_;
  assign new_n21369_ = ~new_n21365_ & new_n21368_;
  assign new_n21370_ = ~new_n21088_ & ~new_n21369_;
  assign new_n21371_ = \b[22]  & ~new_n21077_;
  assign new_n21372_ = ~new_n21075_ & new_n21371_;
  assign new_n21373_ = ~new_n21079_ & ~new_n21372_;
  assign new_n21374_ = ~new_n21370_ & new_n21373_;
  assign new_n21375_ = ~new_n21079_ & ~new_n21374_;
  assign new_n21376_ = \b[23]  & ~new_n21068_;
  assign new_n21377_ = ~new_n21066_ & new_n21376_;
  assign new_n21378_ = ~new_n21070_ & ~new_n21377_;
  assign new_n21379_ = ~new_n21375_ & new_n21378_;
  assign new_n21380_ = ~new_n21070_ & ~new_n21379_;
  assign new_n21381_ = \b[24]  & ~new_n21059_;
  assign new_n21382_ = ~new_n21057_ & new_n21381_;
  assign new_n21383_ = ~new_n21061_ & ~new_n21382_;
  assign new_n21384_ = ~new_n21380_ & new_n21383_;
  assign new_n21385_ = ~new_n21061_ & ~new_n21384_;
  assign new_n21386_ = \b[25]  & ~new_n21050_;
  assign new_n21387_ = ~new_n21048_ & new_n21386_;
  assign new_n21388_ = ~new_n21052_ & ~new_n21387_;
  assign new_n21389_ = ~new_n21385_ & new_n21388_;
  assign new_n21390_ = ~new_n21052_ & ~new_n21389_;
  assign new_n21391_ = \b[26]  & ~new_n21041_;
  assign new_n21392_ = ~new_n21039_ & new_n21391_;
  assign new_n21393_ = ~new_n21043_ & ~new_n21392_;
  assign new_n21394_ = ~new_n21390_ & new_n21393_;
  assign new_n21395_ = ~new_n21043_ & ~new_n21394_;
  assign new_n21396_ = \b[27]  & ~new_n21032_;
  assign new_n21397_ = ~new_n21030_ & new_n21396_;
  assign new_n21398_ = ~new_n21034_ & ~new_n21397_;
  assign new_n21399_ = ~new_n21395_ & new_n21398_;
  assign new_n21400_ = ~new_n21034_ & ~new_n21399_;
  assign new_n21401_ = \b[28]  & ~new_n21023_;
  assign new_n21402_ = ~new_n21021_ & new_n21401_;
  assign new_n21403_ = ~new_n21025_ & ~new_n21402_;
  assign new_n21404_ = ~new_n21400_ & new_n21403_;
  assign new_n21405_ = ~new_n21025_ & ~new_n21404_;
  assign new_n21406_ = \b[29]  & ~new_n21014_;
  assign new_n21407_ = ~new_n21012_ & new_n21406_;
  assign new_n21408_ = ~new_n21016_ & ~new_n21407_;
  assign new_n21409_ = ~new_n21405_ & new_n21408_;
  assign new_n21410_ = ~new_n21016_ & ~new_n21409_;
  assign new_n21411_ = \b[30]  & ~new_n21005_;
  assign new_n21412_ = ~new_n21003_ & new_n21411_;
  assign new_n21413_ = ~new_n21007_ & ~new_n21412_;
  assign new_n21414_ = ~new_n21410_ & new_n21413_;
  assign new_n21415_ = ~new_n21007_ & ~new_n21414_;
  assign new_n21416_ = \b[31]  & ~new_n20996_;
  assign new_n21417_ = ~new_n20994_ & new_n21416_;
  assign new_n21418_ = ~new_n20998_ & ~new_n21417_;
  assign new_n21419_ = ~new_n21415_ & new_n21418_;
  assign new_n21420_ = ~new_n20998_ & ~new_n21419_;
  assign new_n21421_ = \b[32]  & ~new_n20987_;
  assign new_n21422_ = ~new_n20985_ & new_n21421_;
  assign new_n21423_ = ~new_n20989_ & ~new_n21422_;
  assign new_n21424_ = ~new_n21420_ & new_n21423_;
  assign new_n21425_ = ~new_n20989_ & ~new_n21424_;
  assign new_n21426_ = \b[33]  & ~new_n20978_;
  assign new_n21427_ = ~new_n20976_ & new_n21426_;
  assign new_n21428_ = ~new_n20980_ & ~new_n21427_;
  assign new_n21429_ = ~new_n21425_ & new_n21428_;
  assign new_n21430_ = ~new_n20980_ & ~new_n21429_;
  assign new_n21431_ = \b[34]  & ~new_n20969_;
  assign new_n21432_ = ~new_n20967_ & new_n21431_;
  assign new_n21433_ = ~new_n20971_ & ~new_n21432_;
  assign new_n21434_ = ~new_n21430_ & new_n21433_;
  assign new_n21435_ = ~new_n20971_ & ~new_n21434_;
  assign new_n21436_ = \b[35]  & ~new_n20960_;
  assign new_n21437_ = ~new_n20958_ & new_n21436_;
  assign new_n21438_ = ~new_n20962_ & ~new_n21437_;
  assign new_n21439_ = ~new_n21435_ & new_n21438_;
  assign new_n21440_ = ~new_n20962_ & ~new_n21439_;
  assign new_n21441_ = \b[36]  & ~new_n20951_;
  assign new_n21442_ = ~new_n20949_ & new_n21441_;
  assign new_n21443_ = ~new_n20953_ & ~new_n21442_;
  assign new_n21444_ = ~new_n21440_ & new_n21443_;
  assign new_n21445_ = ~new_n20953_ & ~new_n21444_;
  assign new_n21446_ = \b[37]  & ~new_n20942_;
  assign new_n21447_ = ~new_n20940_ & new_n21446_;
  assign new_n21448_ = ~new_n20944_ & ~new_n21447_;
  assign new_n21449_ = ~new_n21445_ & new_n21448_;
  assign new_n21450_ = ~new_n20944_ & ~new_n21449_;
  assign new_n21451_ = \b[38]  & ~new_n20933_;
  assign new_n21452_ = ~new_n20931_ & new_n21451_;
  assign new_n21453_ = ~new_n20935_ & ~new_n21452_;
  assign new_n21454_ = ~new_n21450_ & new_n21453_;
  assign new_n21455_ = ~new_n20935_ & ~new_n21454_;
  assign new_n21456_ = \b[39]  & ~new_n20924_;
  assign new_n21457_ = ~new_n20922_ & new_n21456_;
  assign new_n21458_ = ~new_n20926_ & ~new_n21457_;
  assign new_n21459_ = ~new_n21455_ & new_n21458_;
  assign new_n21460_ = ~new_n20926_ & ~new_n21459_;
  assign new_n21461_ = \b[40]  & ~new_n20915_;
  assign new_n21462_ = ~new_n20913_ & new_n21461_;
  assign new_n21463_ = ~new_n20917_ & ~new_n21462_;
  assign new_n21464_ = ~new_n21460_ & new_n21463_;
  assign new_n21465_ = ~new_n20917_ & ~new_n21464_;
  assign new_n21466_ = \b[41]  & ~new_n20906_;
  assign new_n21467_ = ~new_n20904_ & new_n21466_;
  assign new_n21468_ = ~new_n20908_ & ~new_n21467_;
  assign new_n21469_ = ~new_n21465_ & new_n21468_;
  assign new_n21470_ = ~new_n20908_ & ~new_n21469_;
  assign new_n21471_ = \b[42]  & ~new_n20897_;
  assign new_n21472_ = ~new_n20895_ & new_n21471_;
  assign new_n21473_ = ~new_n20899_ & ~new_n21472_;
  assign new_n21474_ = ~new_n21470_ & new_n21473_;
  assign new_n21475_ = ~new_n20899_ & ~new_n21474_;
  assign new_n21476_ = \b[43]  & ~new_n20888_;
  assign new_n21477_ = ~new_n20886_ & new_n21476_;
  assign new_n21478_ = ~new_n20890_ & ~new_n21477_;
  assign new_n21479_ = ~new_n21475_ & new_n21478_;
  assign new_n21480_ = ~new_n20890_ & ~new_n21479_;
  assign new_n21481_ = \b[44]  & ~new_n20879_;
  assign new_n21482_ = ~new_n20877_ & new_n21481_;
  assign new_n21483_ = ~new_n20881_ & ~new_n21482_;
  assign new_n21484_ = ~new_n21480_ & new_n21483_;
  assign new_n21485_ = ~new_n20881_ & ~new_n21484_;
  assign new_n21486_ = \b[45]  & ~new_n20870_;
  assign new_n21487_ = ~new_n20868_ & new_n21486_;
  assign new_n21488_ = ~new_n20872_ & ~new_n21487_;
  assign new_n21489_ = ~new_n21485_ & new_n21488_;
  assign new_n21490_ = ~new_n20872_ & ~new_n21489_;
  assign new_n21491_ = \b[46]  & ~new_n20861_;
  assign new_n21492_ = ~new_n20859_ & new_n21491_;
  assign new_n21493_ = ~new_n20863_ & ~new_n21492_;
  assign new_n21494_ = ~new_n21490_ & new_n21493_;
  assign new_n21495_ = ~new_n20863_ & ~new_n21494_;
  assign new_n21496_ = \b[47]  & ~new_n20852_;
  assign new_n21497_ = ~new_n20850_ & new_n21496_;
  assign new_n21498_ = ~new_n20854_ & ~new_n21497_;
  assign new_n21499_ = ~new_n21495_ & new_n21498_;
  assign new_n21500_ = ~new_n20854_ & ~new_n21499_;
  assign new_n21501_ = \b[48]  & ~new_n20843_;
  assign new_n21502_ = ~new_n20841_ & new_n21501_;
  assign new_n21503_ = ~new_n20845_ & ~new_n21502_;
  assign new_n21504_ = ~new_n21500_ & new_n21503_;
  assign new_n21505_ = ~new_n20845_ & ~new_n21504_;
  assign new_n21506_ = \b[49]  & ~new_n20834_;
  assign new_n21507_ = ~new_n20832_ & new_n21506_;
  assign new_n21508_ = ~new_n20836_ & ~new_n21507_;
  assign new_n21509_ = ~new_n21505_ & new_n21508_;
  assign new_n21510_ = ~new_n20836_ & ~new_n21509_;
  assign new_n21511_ = \b[50]  & ~new_n20825_;
  assign new_n21512_ = ~new_n20823_ & new_n21511_;
  assign new_n21513_ = ~new_n20827_ & ~new_n21512_;
  assign new_n21514_ = ~new_n21510_ & new_n21513_;
  assign new_n21515_ = ~new_n20827_ & ~new_n21514_;
  assign new_n21516_ = \b[51]  & ~new_n20816_;
  assign new_n21517_ = ~new_n20814_ & new_n21516_;
  assign new_n21518_ = ~new_n20818_ & ~new_n21517_;
  assign new_n21519_ = ~new_n21515_ & new_n21518_;
  assign new_n21520_ = ~new_n20818_ & ~new_n21519_;
  assign new_n21521_ = \b[52]  & ~new_n20807_;
  assign new_n21522_ = ~new_n20805_ & new_n21521_;
  assign new_n21523_ = ~new_n20809_ & ~new_n21522_;
  assign new_n21524_ = ~new_n21520_ & new_n21523_;
  assign new_n21525_ = ~new_n20809_ & ~new_n21524_;
  assign new_n21526_ = \b[53]  & ~new_n20787_;
  assign new_n21527_ = ~new_n20785_ & new_n21526_;
  assign new_n21528_ = ~new_n20800_ & ~new_n21527_;
  assign new_n21529_ = ~new_n21525_ & new_n21528_;
  assign new_n21530_ = ~new_n20800_ & ~new_n21529_;
  assign new_n21531_ = \b[54]  & ~new_n20797_;
  assign new_n21532_ = ~new_n20795_ & new_n21531_;
  assign new_n21533_ = ~new_n20799_ & ~new_n21532_;
  assign new_n21534_ = ~new_n21530_ & new_n21533_;
  assign new_n21535_ = ~new_n20799_ & ~new_n21534_;
  assign new_n21536_ = new_n396_ & new_n406_;
  assign new_n21537_ = new_n403_ & new_n21536_;
  assign \quotient[9]  = ~new_n21535_ & new_n21537_;
  assign new_n21539_ = ~new_n20788_ & ~\quotient[9] ;
  assign new_n21540_ = ~new_n20809_ & new_n21528_;
  assign new_n21541_ = ~new_n21524_ & new_n21540_;
  assign new_n21542_ = ~new_n21525_ & ~new_n21528_;
  assign new_n21543_ = ~new_n21541_ & ~new_n21542_;
  assign new_n21544_ = new_n21537_ & ~new_n21543_;
  assign new_n21545_ = ~new_n21535_ & new_n21544_;
  assign new_n21546_ = ~new_n21539_ & ~new_n21545_;
  assign new_n21547_ = ~\b[54]  & ~new_n21546_;
  assign new_n21548_ = ~new_n20808_ & ~\quotient[9] ;
  assign new_n21549_ = ~new_n20818_ & new_n21523_;
  assign new_n21550_ = ~new_n21519_ & new_n21549_;
  assign new_n21551_ = ~new_n21520_ & ~new_n21523_;
  assign new_n21552_ = ~new_n21550_ & ~new_n21551_;
  assign new_n21553_ = new_n21537_ & ~new_n21552_;
  assign new_n21554_ = ~new_n21535_ & new_n21553_;
  assign new_n21555_ = ~new_n21548_ & ~new_n21554_;
  assign new_n21556_ = ~\b[53]  & ~new_n21555_;
  assign new_n21557_ = ~new_n20817_ & ~\quotient[9] ;
  assign new_n21558_ = ~new_n20827_ & new_n21518_;
  assign new_n21559_ = ~new_n21514_ & new_n21558_;
  assign new_n21560_ = ~new_n21515_ & ~new_n21518_;
  assign new_n21561_ = ~new_n21559_ & ~new_n21560_;
  assign new_n21562_ = new_n21537_ & ~new_n21561_;
  assign new_n21563_ = ~new_n21535_ & new_n21562_;
  assign new_n21564_ = ~new_n21557_ & ~new_n21563_;
  assign new_n21565_ = ~\b[52]  & ~new_n21564_;
  assign new_n21566_ = ~new_n20826_ & ~\quotient[9] ;
  assign new_n21567_ = ~new_n20836_ & new_n21513_;
  assign new_n21568_ = ~new_n21509_ & new_n21567_;
  assign new_n21569_ = ~new_n21510_ & ~new_n21513_;
  assign new_n21570_ = ~new_n21568_ & ~new_n21569_;
  assign new_n21571_ = new_n21537_ & ~new_n21570_;
  assign new_n21572_ = ~new_n21535_ & new_n21571_;
  assign new_n21573_ = ~new_n21566_ & ~new_n21572_;
  assign new_n21574_ = ~\b[51]  & ~new_n21573_;
  assign new_n21575_ = ~new_n20835_ & ~\quotient[9] ;
  assign new_n21576_ = ~new_n20845_ & new_n21508_;
  assign new_n21577_ = ~new_n21504_ & new_n21576_;
  assign new_n21578_ = ~new_n21505_ & ~new_n21508_;
  assign new_n21579_ = ~new_n21577_ & ~new_n21578_;
  assign new_n21580_ = new_n21537_ & ~new_n21579_;
  assign new_n21581_ = ~new_n21535_ & new_n21580_;
  assign new_n21582_ = ~new_n21575_ & ~new_n21581_;
  assign new_n21583_ = ~\b[50]  & ~new_n21582_;
  assign new_n21584_ = ~new_n20844_ & ~\quotient[9] ;
  assign new_n21585_ = ~new_n20854_ & new_n21503_;
  assign new_n21586_ = ~new_n21499_ & new_n21585_;
  assign new_n21587_ = ~new_n21500_ & ~new_n21503_;
  assign new_n21588_ = ~new_n21586_ & ~new_n21587_;
  assign new_n21589_ = new_n21537_ & ~new_n21588_;
  assign new_n21590_ = ~new_n21535_ & new_n21589_;
  assign new_n21591_ = ~new_n21584_ & ~new_n21590_;
  assign new_n21592_ = ~\b[49]  & ~new_n21591_;
  assign new_n21593_ = ~new_n20853_ & ~\quotient[9] ;
  assign new_n21594_ = ~new_n20863_ & new_n21498_;
  assign new_n21595_ = ~new_n21494_ & new_n21594_;
  assign new_n21596_ = ~new_n21495_ & ~new_n21498_;
  assign new_n21597_ = ~new_n21595_ & ~new_n21596_;
  assign new_n21598_ = new_n21537_ & ~new_n21597_;
  assign new_n21599_ = ~new_n21535_ & new_n21598_;
  assign new_n21600_ = ~new_n21593_ & ~new_n21599_;
  assign new_n21601_ = ~\b[48]  & ~new_n21600_;
  assign new_n21602_ = ~new_n20862_ & ~\quotient[9] ;
  assign new_n21603_ = ~new_n20872_ & new_n21493_;
  assign new_n21604_ = ~new_n21489_ & new_n21603_;
  assign new_n21605_ = ~new_n21490_ & ~new_n21493_;
  assign new_n21606_ = ~new_n21604_ & ~new_n21605_;
  assign new_n21607_ = new_n21537_ & ~new_n21606_;
  assign new_n21608_ = ~new_n21535_ & new_n21607_;
  assign new_n21609_ = ~new_n21602_ & ~new_n21608_;
  assign new_n21610_ = ~\b[47]  & ~new_n21609_;
  assign new_n21611_ = ~new_n20871_ & ~\quotient[9] ;
  assign new_n21612_ = ~new_n20881_ & new_n21488_;
  assign new_n21613_ = ~new_n21484_ & new_n21612_;
  assign new_n21614_ = ~new_n21485_ & ~new_n21488_;
  assign new_n21615_ = ~new_n21613_ & ~new_n21614_;
  assign new_n21616_ = new_n21537_ & ~new_n21615_;
  assign new_n21617_ = ~new_n21535_ & new_n21616_;
  assign new_n21618_ = ~new_n21611_ & ~new_n21617_;
  assign new_n21619_ = ~\b[46]  & ~new_n21618_;
  assign new_n21620_ = ~new_n20880_ & ~\quotient[9] ;
  assign new_n21621_ = ~new_n20890_ & new_n21483_;
  assign new_n21622_ = ~new_n21479_ & new_n21621_;
  assign new_n21623_ = ~new_n21480_ & ~new_n21483_;
  assign new_n21624_ = ~new_n21622_ & ~new_n21623_;
  assign new_n21625_ = new_n21537_ & ~new_n21624_;
  assign new_n21626_ = ~new_n21535_ & new_n21625_;
  assign new_n21627_ = ~new_n21620_ & ~new_n21626_;
  assign new_n21628_ = ~\b[45]  & ~new_n21627_;
  assign new_n21629_ = ~new_n20889_ & ~\quotient[9] ;
  assign new_n21630_ = ~new_n20899_ & new_n21478_;
  assign new_n21631_ = ~new_n21474_ & new_n21630_;
  assign new_n21632_ = ~new_n21475_ & ~new_n21478_;
  assign new_n21633_ = ~new_n21631_ & ~new_n21632_;
  assign new_n21634_ = new_n21537_ & ~new_n21633_;
  assign new_n21635_ = ~new_n21535_ & new_n21634_;
  assign new_n21636_ = ~new_n21629_ & ~new_n21635_;
  assign new_n21637_ = ~\b[44]  & ~new_n21636_;
  assign new_n21638_ = ~new_n20898_ & ~\quotient[9] ;
  assign new_n21639_ = ~new_n20908_ & new_n21473_;
  assign new_n21640_ = ~new_n21469_ & new_n21639_;
  assign new_n21641_ = ~new_n21470_ & ~new_n21473_;
  assign new_n21642_ = ~new_n21640_ & ~new_n21641_;
  assign new_n21643_ = new_n21537_ & ~new_n21642_;
  assign new_n21644_ = ~new_n21535_ & new_n21643_;
  assign new_n21645_ = ~new_n21638_ & ~new_n21644_;
  assign new_n21646_ = ~\b[43]  & ~new_n21645_;
  assign new_n21647_ = ~new_n20907_ & ~\quotient[9] ;
  assign new_n21648_ = ~new_n20917_ & new_n21468_;
  assign new_n21649_ = ~new_n21464_ & new_n21648_;
  assign new_n21650_ = ~new_n21465_ & ~new_n21468_;
  assign new_n21651_ = ~new_n21649_ & ~new_n21650_;
  assign new_n21652_ = new_n21537_ & ~new_n21651_;
  assign new_n21653_ = ~new_n21535_ & new_n21652_;
  assign new_n21654_ = ~new_n21647_ & ~new_n21653_;
  assign new_n21655_ = ~\b[42]  & ~new_n21654_;
  assign new_n21656_ = ~new_n20916_ & ~\quotient[9] ;
  assign new_n21657_ = ~new_n20926_ & new_n21463_;
  assign new_n21658_ = ~new_n21459_ & new_n21657_;
  assign new_n21659_ = ~new_n21460_ & ~new_n21463_;
  assign new_n21660_ = ~new_n21658_ & ~new_n21659_;
  assign new_n21661_ = new_n21537_ & ~new_n21660_;
  assign new_n21662_ = ~new_n21535_ & new_n21661_;
  assign new_n21663_ = ~new_n21656_ & ~new_n21662_;
  assign new_n21664_ = ~\b[41]  & ~new_n21663_;
  assign new_n21665_ = ~new_n20925_ & ~\quotient[9] ;
  assign new_n21666_ = ~new_n20935_ & new_n21458_;
  assign new_n21667_ = ~new_n21454_ & new_n21666_;
  assign new_n21668_ = ~new_n21455_ & ~new_n21458_;
  assign new_n21669_ = ~new_n21667_ & ~new_n21668_;
  assign new_n21670_ = new_n21537_ & ~new_n21669_;
  assign new_n21671_ = ~new_n21535_ & new_n21670_;
  assign new_n21672_ = ~new_n21665_ & ~new_n21671_;
  assign new_n21673_ = ~\b[40]  & ~new_n21672_;
  assign new_n21674_ = ~new_n20934_ & ~\quotient[9] ;
  assign new_n21675_ = ~new_n20944_ & new_n21453_;
  assign new_n21676_ = ~new_n21449_ & new_n21675_;
  assign new_n21677_ = ~new_n21450_ & ~new_n21453_;
  assign new_n21678_ = ~new_n21676_ & ~new_n21677_;
  assign new_n21679_ = new_n21537_ & ~new_n21678_;
  assign new_n21680_ = ~new_n21535_ & new_n21679_;
  assign new_n21681_ = ~new_n21674_ & ~new_n21680_;
  assign new_n21682_ = ~\b[39]  & ~new_n21681_;
  assign new_n21683_ = ~new_n20943_ & ~\quotient[9] ;
  assign new_n21684_ = ~new_n20953_ & new_n21448_;
  assign new_n21685_ = ~new_n21444_ & new_n21684_;
  assign new_n21686_ = ~new_n21445_ & ~new_n21448_;
  assign new_n21687_ = ~new_n21685_ & ~new_n21686_;
  assign new_n21688_ = new_n21537_ & ~new_n21687_;
  assign new_n21689_ = ~new_n21535_ & new_n21688_;
  assign new_n21690_ = ~new_n21683_ & ~new_n21689_;
  assign new_n21691_ = ~\b[38]  & ~new_n21690_;
  assign new_n21692_ = ~new_n20952_ & ~\quotient[9] ;
  assign new_n21693_ = ~new_n20962_ & new_n21443_;
  assign new_n21694_ = ~new_n21439_ & new_n21693_;
  assign new_n21695_ = ~new_n21440_ & ~new_n21443_;
  assign new_n21696_ = ~new_n21694_ & ~new_n21695_;
  assign new_n21697_ = new_n21537_ & ~new_n21696_;
  assign new_n21698_ = ~new_n21535_ & new_n21697_;
  assign new_n21699_ = ~new_n21692_ & ~new_n21698_;
  assign new_n21700_ = ~\b[37]  & ~new_n21699_;
  assign new_n21701_ = ~new_n20961_ & ~\quotient[9] ;
  assign new_n21702_ = ~new_n20971_ & new_n21438_;
  assign new_n21703_ = ~new_n21434_ & new_n21702_;
  assign new_n21704_ = ~new_n21435_ & ~new_n21438_;
  assign new_n21705_ = ~new_n21703_ & ~new_n21704_;
  assign new_n21706_ = new_n21537_ & ~new_n21705_;
  assign new_n21707_ = ~new_n21535_ & new_n21706_;
  assign new_n21708_ = ~new_n21701_ & ~new_n21707_;
  assign new_n21709_ = ~\b[36]  & ~new_n21708_;
  assign new_n21710_ = ~new_n20970_ & ~\quotient[9] ;
  assign new_n21711_ = ~new_n20980_ & new_n21433_;
  assign new_n21712_ = ~new_n21429_ & new_n21711_;
  assign new_n21713_ = ~new_n21430_ & ~new_n21433_;
  assign new_n21714_ = ~new_n21712_ & ~new_n21713_;
  assign new_n21715_ = new_n21537_ & ~new_n21714_;
  assign new_n21716_ = ~new_n21535_ & new_n21715_;
  assign new_n21717_ = ~new_n21710_ & ~new_n21716_;
  assign new_n21718_ = ~\b[35]  & ~new_n21717_;
  assign new_n21719_ = ~new_n20979_ & ~\quotient[9] ;
  assign new_n21720_ = ~new_n20989_ & new_n21428_;
  assign new_n21721_ = ~new_n21424_ & new_n21720_;
  assign new_n21722_ = ~new_n21425_ & ~new_n21428_;
  assign new_n21723_ = ~new_n21721_ & ~new_n21722_;
  assign new_n21724_ = new_n21537_ & ~new_n21723_;
  assign new_n21725_ = ~new_n21535_ & new_n21724_;
  assign new_n21726_ = ~new_n21719_ & ~new_n21725_;
  assign new_n21727_ = ~\b[34]  & ~new_n21726_;
  assign new_n21728_ = ~new_n20988_ & ~\quotient[9] ;
  assign new_n21729_ = ~new_n20998_ & new_n21423_;
  assign new_n21730_ = ~new_n21419_ & new_n21729_;
  assign new_n21731_ = ~new_n21420_ & ~new_n21423_;
  assign new_n21732_ = ~new_n21730_ & ~new_n21731_;
  assign new_n21733_ = new_n21537_ & ~new_n21732_;
  assign new_n21734_ = ~new_n21535_ & new_n21733_;
  assign new_n21735_ = ~new_n21728_ & ~new_n21734_;
  assign new_n21736_ = ~\b[33]  & ~new_n21735_;
  assign new_n21737_ = ~new_n20997_ & ~\quotient[9] ;
  assign new_n21738_ = ~new_n21007_ & new_n21418_;
  assign new_n21739_ = ~new_n21414_ & new_n21738_;
  assign new_n21740_ = ~new_n21415_ & ~new_n21418_;
  assign new_n21741_ = ~new_n21739_ & ~new_n21740_;
  assign new_n21742_ = new_n21537_ & ~new_n21741_;
  assign new_n21743_ = ~new_n21535_ & new_n21742_;
  assign new_n21744_ = ~new_n21737_ & ~new_n21743_;
  assign new_n21745_ = ~\b[32]  & ~new_n21744_;
  assign new_n21746_ = ~new_n21006_ & ~\quotient[9] ;
  assign new_n21747_ = ~new_n21016_ & new_n21413_;
  assign new_n21748_ = ~new_n21409_ & new_n21747_;
  assign new_n21749_ = ~new_n21410_ & ~new_n21413_;
  assign new_n21750_ = ~new_n21748_ & ~new_n21749_;
  assign new_n21751_ = new_n21537_ & ~new_n21750_;
  assign new_n21752_ = ~new_n21535_ & new_n21751_;
  assign new_n21753_ = ~new_n21746_ & ~new_n21752_;
  assign new_n21754_ = ~\b[31]  & ~new_n21753_;
  assign new_n21755_ = ~new_n21015_ & ~\quotient[9] ;
  assign new_n21756_ = ~new_n21025_ & new_n21408_;
  assign new_n21757_ = ~new_n21404_ & new_n21756_;
  assign new_n21758_ = ~new_n21405_ & ~new_n21408_;
  assign new_n21759_ = ~new_n21757_ & ~new_n21758_;
  assign new_n21760_ = new_n21537_ & ~new_n21759_;
  assign new_n21761_ = ~new_n21535_ & new_n21760_;
  assign new_n21762_ = ~new_n21755_ & ~new_n21761_;
  assign new_n21763_ = ~\b[30]  & ~new_n21762_;
  assign new_n21764_ = ~new_n21024_ & ~\quotient[9] ;
  assign new_n21765_ = ~new_n21034_ & new_n21403_;
  assign new_n21766_ = ~new_n21399_ & new_n21765_;
  assign new_n21767_ = ~new_n21400_ & ~new_n21403_;
  assign new_n21768_ = ~new_n21766_ & ~new_n21767_;
  assign new_n21769_ = new_n21537_ & ~new_n21768_;
  assign new_n21770_ = ~new_n21535_ & new_n21769_;
  assign new_n21771_ = ~new_n21764_ & ~new_n21770_;
  assign new_n21772_ = ~\b[29]  & ~new_n21771_;
  assign new_n21773_ = ~new_n21033_ & ~\quotient[9] ;
  assign new_n21774_ = ~new_n21043_ & new_n21398_;
  assign new_n21775_ = ~new_n21394_ & new_n21774_;
  assign new_n21776_ = ~new_n21395_ & ~new_n21398_;
  assign new_n21777_ = ~new_n21775_ & ~new_n21776_;
  assign new_n21778_ = new_n21537_ & ~new_n21777_;
  assign new_n21779_ = ~new_n21535_ & new_n21778_;
  assign new_n21780_ = ~new_n21773_ & ~new_n21779_;
  assign new_n21781_ = ~\b[28]  & ~new_n21780_;
  assign new_n21782_ = ~new_n21042_ & ~\quotient[9] ;
  assign new_n21783_ = ~new_n21052_ & new_n21393_;
  assign new_n21784_ = ~new_n21389_ & new_n21783_;
  assign new_n21785_ = ~new_n21390_ & ~new_n21393_;
  assign new_n21786_ = ~new_n21784_ & ~new_n21785_;
  assign new_n21787_ = new_n21537_ & ~new_n21786_;
  assign new_n21788_ = ~new_n21535_ & new_n21787_;
  assign new_n21789_ = ~new_n21782_ & ~new_n21788_;
  assign new_n21790_ = ~\b[27]  & ~new_n21789_;
  assign new_n21791_ = ~new_n21051_ & ~\quotient[9] ;
  assign new_n21792_ = ~new_n21061_ & new_n21388_;
  assign new_n21793_ = ~new_n21384_ & new_n21792_;
  assign new_n21794_ = ~new_n21385_ & ~new_n21388_;
  assign new_n21795_ = ~new_n21793_ & ~new_n21794_;
  assign new_n21796_ = new_n21537_ & ~new_n21795_;
  assign new_n21797_ = ~new_n21535_ & new_n21796_;
  assign new_n21798_ = ~new_n21791_ & ~new_n21797_;
  assign new_n21799_ = ~\b[26]  & ~new_n21798_;
  assign new_n21800_ = ~new_n21060_ & ~\quotient[9] ;
  assign new_n21801_ = ~new_n21070_ & new_n21383_;
  assign new_n21802_ = ~new_n21379_ & new_n21801_;
  assign new_n21803_ = ~new_n21380_ & ~new_n21383_;
  assign new_n21804_ = ~new_n21802_ & ~new_n21803_;
  assign new_n21805_ = new_n21537_ & ~new_n21804_;
  assign new_n21806_ = ~new_n21535_ & new_n21805_;
  assign new_n21807_ = ~new_n21800_ & ~new_n21806_;
  assign new_n21808_ = ~\b[25]  & ~new_n21807_;
  assign new_n21809_ = ~new_n21069_ & ~\quotient[9] ;
  assign new_n21810_ = ~new_n21079_ & new_n21378_;
  assign new_n21811_ = ~new_n21374_ & new_n21810_;
  assign new_n21812_ = ~new_n21375_ & ~new_n21378_;
  assign new_n21813_ = ~new_n21811_ & ~new_n21812_;
  assign new_n21814_ = new_n21537_ & ~new_n21813_;
  assign new_n21815_ = ~new_n21535_ & new_n21814_;
  assign new_n21816_ = ~new_n21809_ & ~new_n21815_;
  assign new_n21817_ = ~\b[24]  & ~new_n21816_;
  assign new_n21818_ = ~new_n21078_ & ~\quotient[9] ;
  assign new_n21819_ = ~new_n21088_ & new_n21373_;
  assign new_n21820_ = ~new_n21369_ & new_n21819_;
  assign new_n21821_ = ~new_n21370_ & ~new_n21373_;
  assign new_n21822_ = ~new_n21820_ & ~new_n21821_;
  assign new_n21823_ = new_n21537_ & ~new_n21822_;
  assign new_n21824_ = ~new_n21535_ & new_n21823_;
  assign new_n21825_ = ~new_n21818_ & ~new_n21824_;
  assign new_n21826_ = ~\b[23]  & ~new_n21825_;
  assign new_n21827_ = ~new_n21087_ & ~\quotient[9] ;
  assign new_n21828_ = ~new_n21097_ & new_n21368_;
  assign new_n21829_ = ~new_n21364_ & new_n21828_;
  assign new_n21830_ = ~new_n21365_ & ~new_n21368_;
  assign new_n21831_ = ~new_n21829_ & ~new_n21830_;
  assign new_n21832_ = new_n21537_ & ~new_n21831_;
  assign new_n21833_ = ~new_n21535_ & new_n21832_;
  assign new_n21834_ = ~new_n21827_ & ~new_n21833_;
  assign new_n21835_ = ~\b[22]  & ~new_n21834_;
  assign new_n21836_ = ~new_n21096_ & ~\quotient[9] ;
  assign new_n21837_ = ~new_n21106_ & new_n21363_;
  assign new_n21838_ = ~new_n21359_ & new_n21837_;
  assign new_n21839_ = ~new_n21360_ & ~new_n21363_;
  assign new_n21840_ = ~new_n21838_ & ~new_n21839_;
  assign new_n21841_ = new_n21537_ & ~new_n21840_;
  assign new_n21842_ = ~new_n21535_ & new_n21841_;
  assign new_n21843_ = ~new_n21836_ & ~new_n21842_;
  assign new_n21844_ = ~\b[21]  & ~new_n21843_;
  assign new_n21845_ = ~new_n21105_ & ~\quotient[9] ;
  assign new_n21846_ = ~new_n21115_ & new_n21358_;
  assign new_n21847_ = ~new_n21354_ & new_n21846_;
  assign new_n21848_ = ~new_n21355_ & ~new_n21358_;
  assign new_n21849_ = ~new_n21847_ & ~new_n21848_;
  assign new_n21850_ = new_n21537_ & ~new_n21849_;
  assign new_n21851_ = ~new_n21535_ & new_n21850_;
  assign new_n21852_ = ~new_n21845_ & ~new_n21851_;
  assign new_n21853_ = ~\b[20]  & ~new_n21852_;
  assign new_n21854_ = ~new_n21114_ & ~\quotient[9] ;
  assign new_n21855_ = ~new_n21124_ & new_n21353_;
  assign new_n21856_ = ~new_n21349_ & new_n21855_;
  assign new_n21857_ = ~new_n21350_ & ~new_n21353_;
  assign new_n21858_ = ~new_n21856_ & ~new_n21857_;
  assign new_n21859_ = new_n21537_ & ~new_n21858_;
  assign new_n21860_ = ~new_n21535_ & new_n21859_;
  assign new_n21861_ = ~new_n21854_ & ~new_n21860_;
  assign new_n21862_ = ~\b[19]  & ~new_n21861_;
  assign new_n21863_ = ~new_n21123_ & ~\quotient[9] ;
  assign new_n21864_ = ~new_n21133_ & new_n21348_;
  assign new_n21865_ = ~new_n21344_ & new_n21864_;
  assign new_n21866_ = ~new_n21345_ & ~new_n21348_;
  assign new_n21867_ = ~new_n21865_ & ~new_n21866_;
  assign new_n21868_ = new_n21537_ & ~new_n21867_;
  assign new_n21869_ = ~new_n21535_ & new_n21868_;
  assign new_n21870_ = ~new_n21863_ & ~new_n21869_;
  assign new_n21871_ = ~\b[18]  & ~new_n21870_;
  assign new_n21872_ = ~new_n21132_ & ~\quotient[9] ;
  assign new_n21873_ = ~new_n21142_ & new_n21343_;
  assign new_n21874_ = ~new_n21339_ & new_n21873_;
  assign new_n21875_ = ~new_n21340_ & ~new_n21343_;
  assign new_n21876_ = ~new_n21874_ & ~new_n21875_;
  assign new_n21877_ = new_n21537_ & ~new_n21876_;
  assign new_n21878_ = ~new_n21535_ & new_n21877_;
  assign new_n21879_ = ~new_n21872_ & ~new_n21878_;
  assign new_n21880_ = ~\b[17]  & ~new_n21879_;
  assign new_n21881_ = ~new_n21141_ & ~\quotient[9] ;
  assign new_n21882_ = ~new_n21151_ & new_n21338_;
  assign new_n21883_ = ~new_n21334_ & new_n21882_;
  assign new_n21884_ = ~new_n21335_ & ~new_n21338_;
  assign new_n21885_ = ~new_n21883_ & ~new_n21884_;
  assign new_n21886_ = new_n21537_ & ~new_n21885_;
  assign new_n21887_ = ~new_n21535_ & new_n21886_;
  assign new_n21888_ = ~new_n21881_ & ~new_n21887_;
  assign new_n21889_ = ~\b[16]  & ~new_n21888_;
  assign new_n21890_ = ~new_n21150_ & ~\quotient[9] ;
  assign new_n21891_ = ~new_n21160_ & new_n21333_;
  assign new_n21892_ = ~new_n21329_ & new_n21891_;
  assign new_n21893_ = ~new_n21330_ & ~new_n21333_;
  assign new_n21894_ = ~new_n21892_ & ~new_n21893_;
  assign new_n21895_ = new_n21537_ & ~new_n21894_;
  assign new_n21896_ = ~new_n21535_ & new_n21895_;
  assign new_n21897_ = ~new_n21890_ & ~new_n21896_;
  assign new_n21898_ = ~\b[15]  & ~new_n21897_;
  assign new_n21899_ = ~new_n21159_ & ~\quotient[9] ;
  assign new_n21900_ = ~new_n21169_ & new_n21328_;
  assign new_n21901_ = ~new_n21324_ & new_n21900_;
  assign new_n21902_ = ~new_n21325_ & ~new_n21328_;
  assign new_n21903_ = ~new_n21901_ & ~new_n21902_;
  assign new_n21904_ = new_n21537_ & ~new_n21903_;
  assign new_n21905_ = ~new_n21535_ & new_n21904_;
  assign new_n21906_ = ~new_n21899_ & ~new_n21905_;
  assign new_n21907_ = ~\b[14]  & ~new_n21906_;
  assign new_n21908_ = ~new_n21168_ & ~\quotient[9] ;
  assign new_n21909_ = ~new_n21178_ & new_n21323_;
  assign new_n21910_ = ~new_n21319_ & new_n21909_;
  assign new_n21911_ = ~new_n21320_ & ~new_n21323_;
  assign new_n21912_ = ~new_n21910_ & ~new_n21911_;
  assign new_n21913_ = new_n21537_ & ~new_n21912_;
  assign new_n21914_ = ~new_n21535_ & new_n21913_;
  assign new_n21915_ = ~new_n21908_ & ~new_n21914_;
  assign new_n21916_ = ~\b[13]  & ~new_n21915_;
  assign new_n21917_ = ~new_n21177_ & ~\quotient[9] ;
  assign new_n21918_ = ~new_n21187_ & new_n21318_;
  assign new_n21919_ = ~new_n21314_ & new_n21918_;
  assign new_n21920_ = ~new_n21315_ & ~new_n21318_;
  assign new_n21921_ = ~new_n21919_ & ~new_n21920_;
  assign new_n21922_ = new_n21537_ & ~new_n21921_;
  assign new_n21923_ = ~new_n21535_ & new_n21922_;
  assign new_n21924_ = ~new_n21917_ & ~new_n21923_;
  assign new_n21925_ = ~\b[12]  & ~new_n21924_;
  assign new_n21926_ = ~new_n21186_ & ~\quotient[9] ;
  assign new_n21927_ = ~new_n21196_ & new_n21313_;
  assign new_n21928_ = ~new_n21309_ & new_n21927_;
  assign new_n21929_ = ~new_n21310_ & ~new_n21313_;
  assign new_n21930_ = ~new_n21928_ & ~new_n21929_;
  assign new_n21931_ = new_n21537_ & ~new_n21930_;
  assign new_n21932_ = ~new_n21535_ & new_n21931_;
  assign new_n21933_ = ~new_n21926_ & ~new_n21932_;
  assign new_n21934_ = ~\b[11]  & ~new_n21933_;
  assign new_n21935_ = ~new_n21195_ & ~\quotient[9] ;
  assign new_n21936_ = ~new_n21205_ & new_n21308_;
  assign new_n21937_ = ~new_n21304_ & new_n21936_;
  assign new_n21938_ = ~new_n21305_ & ~new_n21308_;
  assign new_n21939_ = ~new_n21937_ & ~new_n21938_;
  assign new_n21940_ = new_n21537_ & ~new_n21939_;
  assign new_n21941_ = ~new_n21535_ & new_n21940_;
  assign new_n21942_ = ~new_n21935_ & ~new_n21941_;
  assign new_n21943_ = ~\b[10]  & ~new_n21942_;
  assign new_n21944_ = ~new_n21204_ & ~\quotient[9] ;
  assign new_n21945_ = ~new_n21214_ & new_n21303_;
  assign new_n21946_ = ~new_n21299_ & new_n21945_;
  assign new_n21947_ = ~new_n21300_ & ~new_n21303_;
  assign new_n21948_ = ~new_n21946_ & ~new_n21947_;
  assign new_n21949_ = new_n21537_ & ~new_n21948_;
  assign new_n21950_ = ~new_n21535_ & new_n21949_;
  assign new_n21951_ = ~new_n21944_ & ~new_n21950_;
  assign new_n21952_ = ~\b[9]  & ~new_n21951_;
  assign new_n21953_ = ~new_n21213_ & ~\quotient[9] ;
  assign new_n21954_ = ~new_n21223_ & new_n21298_;
  assign new_n21955_ = ~new_n21294_ & new_n21954_;
  assign new_n21956_ = ~new_n21295_ & ~new_n21298_;
  assign new_n21957_ = ~new_n21955_ & ~new_n21956_;
  assign new_n21958_ = new_n21537_ & ~new_n21957_;
  assign new_n21959_ = ~new_n21535_ & new_n21958_;
  assign new_n21960_ = ~new_n21953_ & ~new_n21959_;
  assign new_n21961_ = ~\b[8]  & ~new_n21960_;
  assign new_n21962_ = ~new_n21222_ & ~\quotient[9] ;
  assign new_n21963_ = ~new_n21232_ & new_n21293_;
  assign new_n21964_ = ~new_n21289_ & new_n21963_;
  assign new_n21965_ = ~new_n21290_ & ~new_n21293_;
  assign new_n21966_ = ~new_n21964_ & ~new_n21965_;
  assign new_n21967_ = new_n21537_ & ~new_n21966_;
  assign new_n21968_ = ~new_n21535_ & new_n21967_;
  assign new_n21969_ = ~new_n21962_ & ~new_n21968_;
  assign new_n21970_ = ~\b[7]  & ~new_n21969_;
  assign new_n21971_ = ~new_n21231_ & ~\quotient[9] ;
  assign new_n21972_ = ~new_n21241_ & new_n21288_;
  assign new_n21973_ = ~new_n21284_ & new_n21972_;
  assign new_n21974_ = ~new_n21285_ & ~new_n21288_;
  assign new_n21975_ = ~new_n21973_ & ~new_n21974_;
  assign new_n21976_ = new_n21537_ & ~new_n21975_;
  assign new_n21977_ = ~new_n21535_ & new_n21976_;
  assign new_n21978_ = ~new_n21971_ & ~new_n21977_;
  assign new_n21979_ = ~\b[6]  & ~new_n21978_;
  assign new_n21980_ = ~new_n21240_ & ~\quotient[9] ;
  assign new_n21981_ = ~new_n21250_ & new_n21283_;
  assign new_n21982_ = ~new_n21279_ & new_n21981_;
  assign new_n21983_ = ~new_n21280_ & ~new_n21283_;
  assign new_n21984_ = ~new_n21982_ & ~new_n21983_;
  assign new_n21985_ = new_n21537_ & ~new_n21984_;
  assign new_n21986_ = ~new_n21535_ & new_n21985_;
  assign new_n21987_ = ~new_n21980_ & ~new_n21986_;
  assign new_n21988_ = ~\b[5]  & ~new_n21987_;
  assign new_n21989_ = ~new_n21249_ & ~\quotient[9] ;
  assign new_n21990_ = ~new_n21258_ & new_n21278_;
  assign new_n21991_ = ~new_n21274_ & new_n21990_;
  assign new_n21992_ = ~new_n21275_ & ~new_n21278_;
  assign new_n21993_ = ~new_n21991_ & ~new_n21992_;
  assign new_n21994_ = new_n21537_ & ~new_n21993_;
  assign new_n21995_ = ~new_n21535_ & new_n21994_;
  assign new_n21996_ = ~new_n21989_ & ~new_n21995_;
  assign new_n21997_ = ~\b[4]  & ~new_n21996_;
  assign new_n21998_ = ~new_n21257_ & ~\quotient[9] ;
  assign new_n21999_ = ~new_n21269_ & new_n21273_;
  assign new_n22000_ = ~new_n21268_ & new_n21999_;
  assign new_n22001_ = ~new_n21270_ & ~new_n21273_;
  assign new_n22002_ = ~new_n22000_ & ~new_n22001_;
  assign new_n22003_ = new_n21537_ & ~new_n22002_;
  assign new_n22004_ = ~new_n21535_ & new_n22003_;
  assign new_n22005_ = ~new_n21998_ & ~new_n22004_;
  assign new_n22006_ = ~\b[3]  & ~new_n22005_;
  assign new_n22007_ = ~new_n21262_ & ~\quotient[9] ;
  assign new_n22008_ = ~new_n21265_ & new_n21267_;
  assign new_n22009_ = ~new_n21263_ & new_n22008_;
  assign new_n22010_ = new_n21537_ & ~new_n22009_;
  assign new_n22011_ = ~new_n21268_ & new_n22010_;
  assign new_n22012_ = ~new_n21535_ & new_n22011_;
  assign new_n22013_ = ~new_n22007_ & ~new_n22012_;
  assign new_n22014_ = ~\b[2]  & ~new_n22013_;
  assign new_n22015_ = \b[0]  & ~\b[55] ;
  assign new_n22016_ = new_n283_ & new_n22015_;
  assign new_n22017_ = new_n280_ & new_n22016_;
  assign new_n22018_ = ~new_n21535_ & new_n22017_;
  assign new_n22019_ = \a[9]  & ~new_n22018_;
  assign new_n22020_ = new_n396_ & new_n21267_;
  assign new_n22021_ = new_n406_ & new_n22020_;
  assign new_n22022_ = new_n403_ & new_n22021_;
  assign new_n22023_ = ~new_n21535_ & new_n22022_;
  assign new_n22024_ = ~new_n22019_ & ~new_n22023_;
  assign new_n22025_ = \b[1]  & ~new_n22024_;
  assign new_n22026_ = ~\b[1]  & ~new_n22023_;
  assign new_n22027_ = ~new_n22019_ & new_n22026_;
  assign new_n22028_ = ~new_n22025_ & ~new_n22027_;
  assign new_n22029_ = ~\a[8]  & \b[0] ;
  assign new_n22030_ = ~new_n22028_ & ~new_n22029_;
  assign new_n22031_ = ~\b[1]  & ~new_n22024_;
  assign new_n22032_ = ~new_n22030_ & ~new_n22031_;
  assign new_n22033_ = \b[2]  & ~new_n22012_;
  assign new_n22034_ = ~new_n22007_ & new_n22033_;
  assign new_n22035_ = ~new_n22014_ & ~new_n22034_;
  assign new_n22036_ = ~new_n22032_ & new_n22035_;
  assign new_n22037_ = ~new_n22014_ & ~new_n22036_;
  assign new_n22038_ = \b[3]  & ~new_n22004_;
  assign new_n22039_ = ~new_n21998_ & new_n22038_;
  assign new_n22040_ = ~new_n22006_ & ~new_n22039_;
  assign new_n22041_ = ~new_n22037_ & new_n22040_;
  assign new_n22042_ = ~new_n22006_ & ~new_n22041_;
  assign new_n22043_ = \b[4]  & ~new_n21995_;
  assign new_n22044_ = ~new_n21989_ & new_n22043_;
  assign new_n22045_ = ~new_n21997_ & ~new_n22044_;
  assign new_n22046_ = ~new_n22042_ & new_n22045_;
  assign new_n22047_ = ~new_n21997_ & ~new_n22046_;
  assign new_n22048_ = \b[5]  & ~new_n21986_;
  assign new_n22049_ = ~new_n21980_ & new_n22048_;
  assign new_n22050_ = ~new_n21988_ & ~new_n22049_;
  assign new_n22051_ = ~new_n22047_ & new_n22050_;
  assign new_n22052_ = ~new_n21988_ & ~new_n22051_;
  assign new_n22053_ = \b[6]  & ~new_n21977_;
  assign new_n22054_ = ~new_n21971_ & new_n22053_;
  assign new_n22055_ = ~new_n21979_ & ~new_n22054_;
  assign new_n22056_ = ~new_n22052_ & new_n22055_;
  assign new_n22057_ = ~new_n21979_ & ~new_n22056_;
  assign new_n22058_ = \b[7]  & ~new_n21968_;
  assign new_n22059_ = ~new_n21962_ & new_n22058_;
  assign new_n22060_ = ~new_n21970_ & ~new_n22059_;
  assign new_n22061_ = ~new_n22057_ & new_n22060_;
  assign new_n22062_ = ~new_n21970_ & ~new_n22061_;
  assign new_n22063_ = \b[8]  & ~new_n21959_;
  assign new_n22064_ = ~new_n21953_ & new_n22063_;
  assign new_n22065_ = ~new_n21961_ & ~new_n22064_;
  assign new_n22066_ = ~new_n22062_ & new_n22065_;
  assign new_n22067_ = ~new_n21961_ & ~new_n22066_;
  assign new_n22068_ = \b[9]  & ~new_n21950_;
  assign new_n22069_ = ~new_n21944_ & new_n22068_;
  assign new_n22070_ = ~new_n21952_ & ~new_n22069_;
  assign new_n22071_ = ~new_n22067_ & new_n22070_;
  assign new_n22072_ = ~new_n21952_ & ~new_n22071_;
  assign new_n22073_ = \b[10]  & ~new_n21941_;
  assign new_n22074_ = ~new_n21935_ & new_n22073_;
  assign new_n22075_ = ~new_n21943_ & ~new_n22074_;
  assign new_n22076_ = ~new_n22072_ & new_n22075_;
  assign new_n22077_ = ~new_n21943_ & ~new_n22076_;
  assign new_n22078_ = \b[11]  & ~new_n21932_;
  assign new_n22079_ = ~new_n21926_ & new_n22078_;
  assign new_n22080_ = ~new_n21934_ & ~new_n22079_;
  assign new_n22081_ = ~new_n22077_ & new_n22080_;
  assign new_n22082_ = ~new_n21934_ & ~new_n22081_;
  assign new_n22083_ = \b[12]  & ~new_n21923_;
  assign new_n22084_ = ~new_n21917_ & new_n22083_;
  assign new_n22085_ = ~new_n21925_ & ~new_n22084_;
  assign new_n22086_ = ~new_n22082_ & new_n22085_;
  assign new_n22087_ = ~new_n21925_ & ~new_n22086_;
  assign new_n22088_ = \b[13]  & ~new_n21914_;
  assign new_n22089_ = ~new_n21908_ & new_n22088_;
  assign new_n22090_ = ~new_n21916_ & ~new_n22089_;
  assign new_n22091_ = ~new_n22087_ & new_n22090_;
  assign new_n22092_ = ~new_n21916_ & ~new_n22091_;
  assign new_n22093_ = \b[14]  & ~new_n21905_;
  assign new_n22094_ = ~new_n21899_ & new_n22093_;
  assign new_n22095_ = ~new_n21907_ & ~new_n22094_;
  assign new_n22096_ = ~new_n22092_ & new_n22095_;
  assign new_n22097_ = ~new_n21907_ & ~new_n22096_;
  assign new_n22098_ = \b[15]  & ~new_n21896_;
  assign new_n22099_ = ~new_n21890_ & new_n22098_;
  assign new_n22100_ = ~new_n21898_ & ~new_n22099_;
  assign new_n22101_ = ~new_n22097_ & new_n22100_;
  assign new_n22102_ = ~new_n21898_ & ~new_n22101_;
  assign new_n22103_ = \b[16]  & ~new_n21887_;
  assign new_n22104_ = ~new_n21881_ & new_n22103_;
  assign new_n22105_ = ~new_n21889_ & ~new_n22104_;
  assign new_n22106_ = ~new_n22102_ & new_n22105_;
  assign new_n22107_ = ~new_n21889_ & ~new_n22106_;
  assign new_n22108_ = \b[17]  & ~new_n21878_;
  assign new_n22109_ = ~new_n21872_ & new_n22108_;
  assign new_n22110_ = ~new_n21880_ & ~new_n22109_;
  assign new_n22111_ = ~new_n22107_ & new_n22110_;
  assign new_n22112_ = ~new_n21880_ & ~new_n22111_;
  assign new_n22113_ = \b[18]  & ~new_n21869_;
  assign new_n22114_ = ~new_n21863_ & new_n22113_;
  assign new_n22115_ = ~new_n21871_ & ~new_n22114_;
  assign new_n22116_ = ~new_n22112_ & new_n22115_;
  assign new_n22117_ = ~new_n21871_ & ~new_n22116_;
  assign new_n22118_ = \b[19]  & ~new_n21860_;
  assign new_n22119_ = ~new_n21854_ & new_n22118_;
  assign new_n22120_ = ~new_n21862_ & ~new_n22119_;
  assign new_n22121_ = ~new_n22117_ & new_n22120_;
  assign new_n22122_ = ~new_n21862_ & ~new_n22121_;
  assign new_n22123_ = \b[20]  & ~new_n21851_;
  assign new_n22124_ = ~new_n21845_ & new_n22123_;
  assign new_n22125_ = ~new_n21853_ & ~new_n22124_;
  assign new_n22126_ = ~new_n22122_ & new_n22125_;
  assign new_n22127_ = ~new_n21853_ & ~new_n22126_;
  assign new_n22128_ = \b[21]  & ~new_n21842_;
  assign new_n22129_ = ~new_n21836_ & new_n22128_;
  assign new_n22130_ = ~new_n21844_ & ~new_n22129_;
  assign new_n22131_ = ~new_n22127_ & new_n22130_;
  assign new_n22132_ = ~new_n21844_ & ~new_n22131_;
  assign new_n22133_ = \b[22]  & ~new_n21833_;
  assign new_n22134_ = ~new_n21827_ & new_n22133_;
  assign new_n22135_ = ~new_n21835_ & ~new_n22134_;
  assign new_n22136_ = ~new_n22132_ & new_n22135_;
  assign new_n22137_ = ~new_n21835_ & ~new_n22136_;
  assign new_n22138_ = \b[23]  & ~new_n21824_;
  assign new_n22139_ = ~new_n21818_ & new_n22138_;
  assign new_n22140_ = ~new_n21826_ & ~new_n22139_;
  assign new_n22141_ = ~new_n22137_ & new_n22140_;
  assign new_n22142_ = ~new_n21826_ & ~new_n22141_;
  assign new_n22143_ = \b[24]  & ~new_n21815_;
  assign new_n22144_ = ~new_n21809_ & new_n22143_;
  assign new_n22145_ = ~new_n21817_ & ~new_n22144_;
  assign new_n22146_ = ~new_n22142_ & new_n22145_;
  assign new_n22147_ = ~new_n21817_ & ~new_n22146_;
  assign new_n22148_ = \b[25]  & ~new_n21806_;
  assign new_n22149_ = ~new_n21800_ & new_n22148_;
  assign new_n22150_ = ~new_n21808_ & ~new_n22149_;
  assign new_n22151_ = ~new_n22147_ & new_n22150_;
  assign new_n22152_ = ~new_n21808_ & ~new_n22151_;
  assign new_n22153_ = \b[26]  & ~new_n21797_;
  assign new_n22154_ = ~new_n21791_ & new_n22153_;
  assign new_n22155_ = ~new_n21799_ & ~new_n22154_;
  assign new_n22156_ = ~new_n22152_ & new_n22155_;
  assign new_n22157_ = ~new_n21799_ & ~new_n22156_;
  assign new_n22158_ = \b[27]  & ~new_n21788_;
  assign new_n22159_ = ~new_n21782_ & new_n22158_;
  assign new_n22160_ = ~new_n21790_ & ~new_n22159_;
  assign new_n22161_ = ~new_n22157_ & new_n22160_;
  assign new_n22162_ = ~new_n21790_ & ~new_n22161_;
  assign new_n22163_ = \b[28]  & ~new_n21779_;
  assign new_n22164_ = ~new_n21773_ & new_n22163_;
  assign new_n22165_ = ~new_n21781_ & ~new_n22164_;
  assign new_n22166_ = ~new_n22162_ & new_n22165_;
  assign new_n22167_ = ~new_n21781_ & ~new_n22166_;
  assign new_n22168_ = \b[29]  & ~new_n21770_;
  assign new_n22169_ = ~new_n21764_ & new_n22168_;
  assign new_n22170_ = ~new_n21772_ & ~new_n22169_;
  assign new_n22171_ = ~new_n22167_ & new_n22170_;
  assign new_n22172_ = ~new_n21772_ & ~new_n22171_;
  assign new_n22173_ = \b[30]  & ~new_n21761_;
  assign new_n22174_ = ~new_n21755_ & new_n22173_;
  assign new_n22175_ = ~new_n21763_ & ~new_n22174_;
  assign new_n22176_ = ~new_n22172_ & new_n22175_;
  assign new_n22177_ = ~new_n21763_ & ~new_n22176_;
  assign new_n22178_ = \b[31]  & ~new_n21752_;
  assign new_n22179_ = ~new_n21746_ & new_n22178_;
  assign new_n22180_ = ~new_n21754_ & ~new_n22179_;
  assign new_n22181_ = ~new_n22177_ & new_n22180_;
  assign new_n22182_ = ~new_n21754_ & ~new_n22181_;
  assign new_n22183_ = \b[32]  & ~new_n21743_;
  assign new_n22184_ = ~new_n21737_ & new_n22183_;
  assign new_n22185_ = ~new_n21745_ & ~new_n22184_;
  assign new_n22186_ = ~new_n22182_ & new_n22185_;
  assign new_n22187_ = ~new_n21745_ & ~new_n22186_;
  assign new_n22188_ = \b[33]  & ~new_n21734_;
  assign new_n22189_ = ~new_n21728_ & new_n22188_;
  assign new_n22190_ = ~new_n21736_ & ~new_n22189_;
  assign new_n22191_ = ~new_n22187_ & new_n22190_;
  assign new_n22192_ = ~new_n21736_ & ~new_n22191_;
  assign new_n22193_ = \b[34]  & ~new_n21725_;
  assign new_n22194_ = ~new_n21719_ & new_n22193_;
  assign new_n22195_ = ~new_n21727_ & ~new_n22194_;
  assign new_n22196_ = ~new_n22192_ & new_n22195_;
  assign new_n22197_ = ~new_n21727_ & ~new_n22196_;
  assign new_n22198_ = \b[35]  & ~new_n21716_;
  assign new_n22199_ = ~new_n21710_ & new_n22198_;
  assign new_n22200_ = ~new_n21718_ & ~new_n22199_;
  assign new_n22201_ = ~new_n22197_ & new_n22200_;
  assign new_n22202_ = ~new_n21718_ & ~new_n22201_;
  assign new_n22203_ = \b[36]  & ~new_n21707_;
  assign new_n22204_ = ~new_n21701_ & new_n22203_;
  assign new_n22205_ = ~new_n21709_ & ~new_n22204_;
  assign new_n22206_ = ~new_n22202_ & new_n22205_;
  assign new_n22207_ = ~new_n21709_ & ~new_n22206_;
  assign new_n22208_ = \b[37]  & ~new_n21698_;
  assign new_n22209_ = ~new_n21692_ & new_n22208_;
  assign new_n22210_ = ~new_n21700_ & ~new_n22209_;
  assign new_n22211_ = ~new_n22207_ & new_n22210_;
  assign new_n22212_ = ~new_n21700_ & ~new_n22211_;
  assign new_n22213_ = \b[38]  & ~new_n21689_;
  assign new_n22214_ = ~new_n21683_ & new_n22213_;
  assign new_n22215_ = ~new_n21691_ & ~new_n22214_;
  assign new_n22216_ = ~new_n22212_ & new_n22215_;
  assign new_n22217_ = ~new_n21691_ & ~new_n22216_;
  assign new_n22218_ = \b[39]  & ~new_n21680_;
  assign new_n22219_ = ~new_n21674_ & new_n22218_;
  assign new_n22220_ = ~new_n21682_ & ~new_n22219_;
  assign new_n22221_ = ~new_n22217_ & new_n22220_;
  assign new_n22222_ = ~new_n21682_ & ~new_n22221_;
  assign new_n22223_ = \b[40]  & ~new_n21671_;
  assign new_n22224_ = ~new_n21665_ & new_n22223_;
  assign new_n22225_ = ~new_n21673_ & ~new_n22224_;
  assign new_n22226_ = ~new_n22222_ & new_n22225_;
  assign new_n22227_ = ~new_n21673_ & ~new_n22226_;
  assign new_n22228_ = \b[41]  & ~new_n21662_;
  assign new_n22229_ = ~new_n21656_ & new_n22228_;
  assign new_n22230_ = ~new_n21664_ & ~new_n22229_;
  assign new_n22231_ = ~new_n22227_ & new_n22230_;
  assign new_n22232_ = ~new_n21664_ & ~new_n22231_;
  assign new_n22233_ = \b[42]  & ~new_n21653_;
  assign new_n22234_ = ~new_n21647_ & new_n22233_;
  assign new_n22235_ = ~new_n21655_ & ~new_n22234_;
  assign new_n22236_ = ~new_n22232_ & new_n22235_;
  assign new_n22237_ = ~new_n21655_ & ~new_n22236_;
  assign new_n22238_ = \b[43]  & ~new_n21644_;
  assign new_n22239_ = ~new_n21638_ & new_n22238_;
  assign new_n22240_ = ~new_n21646_ & ~new_n22239_;
  assign new_n22241_ = ~new_n22237_ & new_n22240_;
  assign new_n22242_ = ~new_n21646_ & ~new_n22241_;
  assign new_n22243_ = \b[44]  & ~new_n21635_;
  assign new_n22244_ = ~new_n21629_ & new_n22243_;
  assign new_n22245_ = ~new_n21637_ & ~new_n22244_;
  assign new_n22246_ = ~new_n22242_ & new_n22245_;
  assign new_n22247_ = ~new_n21637_ & ~new_n22246_;
  assign new_n22248_ = \b[45]  & ~new_n21626_;
  assign new_n22249_ = ~new_n21620_ & new_n22248_;
  assign new_n22250_ = ~new_n21628_ & ~new_n22249_;
  assign new_n22251_ = ~new_n22247_ & new_n22250_;
  assign new_n22252_ = ~new_n21628_ & ~new_n22251_;
  assign new_n22253_ = \b[46]  & ~new_n21617_;
  assign new_n22254_ = ~new_n21611_ & new_n22253_;
  assign new_n22255_ = ~new_n21619_ & ~new_n22254_;
  assign new_n22256_ = ~new_n22252_ & new_n22255_;
  assign new_n22257_ = ~new_n21619_ & ~new_n22256_;
  assign new_n22258_ = \b[47]  & ~new_n21608_;
  assign new_n22259_ = ~new_n21602_ & new_n22258_;
  assign new_n22260_ = ~new_n21610_ & ~new_n22259_;
  assign new_n22261_ = ~new_n22257_ & new_n22260_;
  assign new_n22262_ = ~new_n21610_ & ~new_n22261_;
  assign new_n22263_ = \b[48]  & ~new_n21599_;
  assign new_n22264_ = ~new_n21593_ & new_n22263_;
  assign new_n22265_ = ~new_n21601_ & ~new_n22264_;
  assign new_n22266_ = ~new_n22262_ & new_n22265_;
  assign new_n22267_ = ~new_n21601_ & ~new_n22266_;
  assign new_n22268_ = \b[49]  & ~new_n21590_;
  assign new_n22269_ = ~new_n21584_ & new_n22268_;
  assign new_n22270_ = ~new_n21592_ & ~new_n22269_;
  assign new_n22271_ = ~new_n22267_ & new_n22270_;
  assign new_n22272_ = ~new_n21592_ & ~new_n22271_;
  assign new_n22273_ = \b[50]  & ~new_n21581_;
  assign new_n22274_ = ~new_n21575_ & new_n22273_;
  assign new_n22275_ = ~new_n21583_ & ~new_n22274_;
  assign new_n22276_ = ~new_n22272_ & new_n22275_;
  assign new_n22277_ = ~new_n21583_ & ~new_n22276_;
  assign new_n22278_ = \b[51]  & ~new_n21572_;
  assign new_n22279_ = ~new_n21566_ & new_n22278_;
  assign new_n22280_ = ~new_n21574_ & ~new_n22279_;
  assign new_n22281_ = ~new_n22277_ & new_n22280_;
  assign new_n22282_ = ~new_n21574_ & ~new_n22281_;
  assign new_n22283_ = \b[52]  & ~new_n21563_;
  assign new_n22284_ = ~new_n21557_ & new_n22283_;
  assign new_n22285_ = ~new_n21565_ & ~new_n22284_;
  assign new_n22286_ = ~new_n22282_ & new_n22285_;
  assign new_n22287_ = ~new_n21565_ & ~new_n22286_;
  assign new_n22288_ = \b[53]  & ~new_n21554_;
  assign new_n22289_ = ~new_n21548_ & new_n22288_;
  assign new_n22290_ = ~new_n21556_ & ~new_n22289_;
  assign new_n22291_ = ~new_n22287_ & new_n22290_;
  assign new_n22292_ = ~new_n21556_ & ~new_n22291_;
  assign new_n22293_ = \b[54]  & ~new_n21545_;
  assign new_n22294_ = ~new_n21539_ & new_n22293_;
  assign new_n22295_ = ~new_n21547_ & ~new_n22294_;
  assign new_n22296_ = ~new_n22292_ & new_n22295_;
  assign new_n22297_ = ~new_n21547_ & ~new_n22296_;
  assign new_n22298_ = ~new_n20798_ & ~\quotient[9] ;
  assign new_n22299_ = ~new_n20800_ & new_n21533_;
  assign new_n22300_ = ~new_n21529_ & new_n22299_;
  assign new_n22301_ = ~new_n21530_ & ~new_n21533_;
  assign new_n22302_ = ~new_n22300_ & ~new_n22301_;
  assign new_n22303_ = \quotient[9]  & ~new_n22302_;
  assign new_n22304_ = ~new_n22298_ & ~new_n22303_;
  assign new_n22305_ = ~\b[55]  & ~new_n22304_;
  assign new_n22306_ = \b[55]  & ~new_n22298_;
  assign new_n22307_ = ~new_n22303_ & new_n22306_;
  assign new_n22308_ = new_n337_ & ~new_n22307_;
  assign new_n22309_ = ~new_n22305_ & new_n22308_;
  assign new_n22310_ = ~new_n22297_ & new_n22309_;
  assign new_n22311_ = new_n21537_ & ~new_n22304_;
  assign \quotient[8]  = new_n22310_ | new_n22311_;
  assign new_n22313_ = ~new_n21556_ & new_n22295_;
  assign new_n22314_ = ~new_n22291_ & new_n22313_;
  assign new_n22315_ = ~new_n22292_ & ~new_n22295_;
  assign new_n22316_ = ~new_n22314_ & ~new_n22315_;
  assign new_n22317_ = \quotient[8]  & ~new_n22316_;
  assign new_n22318_ = ~new_n21546_ & ~new_n22311_;
  assign new_n22319_ = ~new_n22310_ & new_n22318_;
  assign new_n22320_ = ~new_n22317_ & ~new_n22319_;
  assign new_n22321_ = ~\b[55]  & ~new_n22320_;
  assign new_n22322_ = ~new_n21565_ & new_n22290_;
  assign new_n22323_ = ~new_n22286_ & new_n22322_;
  assign new_n22324_ = ~new_n22287_ & ~new_n22290_;
  assign new_n22325_ = ~new_n22323_ & ~new_n22324_;
  assign new_n22326_ = \quotient[8]  & ~new_n22325_;
  assign new_n22327_ = ~new_n21555_ & ~new_n22311_;
  assign new_n22328_ = ~new_n22310_ & new_n22327_;
  assign new_n22329_ = ~new_n22326_ & ~new_n22328_;
  assign new_n22330_ = ~\b[54]  & ~new_n22329_;
  assign new_n22331_ = ~new_n21574_ & new_n22285_;
  assign new_n22332_ = ~new_n22281_ & new_n22331_;
  assign new_n22333_ = ~new_n22282_ & ~new_n22285_;
  assign new_n22334_ = ~new_n22332_ & ~new_n22333_;
  assign new_n22335_ = \quotient[8]  & ~new_n22334_;
  assign new_n22336_ = ~new_n21564_ & ~new_n22311_;
  assign new_n22337_ = ~new_n22310_ & new_n22336_;
  assign new_n22338_ = ~new_n22335_ & ~new_n22337_;
  assign new_n22339_ = ~\b[53]  & ~new_n22338_;
  assign new_n22340_ = ~new_n21583_ & new_n22280_;
  assign new_n22341_ = ~new_n22276_ & new_n22340_;
  assign new_n22342_ = ~new_n22277_ & ~new_n22280_;
  assign new_n22343_ = ~new_n22341_ & ~new_n22342_;
  assign new_n22344_ = \quotient[8]  & ~new_n22343_;
  assign new_n22345_ = ~new_n21573_ & ~new_n22311_;
  assign new_n22346_ = ~new_n22310_ & new_n22345_;
  assign new_n22347_ = ~new_n22344_ & ~new_n22346_;
  assign new_n22348_ = ~\b[52]  & ~new_n22347_;
  assign new_n22349_ = ~new_n21592_ & new_n22275_;
  assign new_n22350_ = ~new_n22271_ & new_n22349_;
  assign new_n22351_ = ~new_n22272_ & ~new_n22275_;
  assign new_n22352_ = ~new_n22350_ & ~new_n22351_;
  assign new_n22353_ = \quotient[8]  & ~new_n22352_;
  assign new_n22354_ = ~new_n21582_ & ~new_n22311_;
  assign new_n22355_ = ~new_n22310_ & new_n22354_;
  assign new_n22356_ = ~new_n22353_ & ~new_n22355_;
  assign new_n22357_ = ~\b[51]  & ~new_n22356_;
  assign new_n22358_ = ~new_n21601_ & new_n22270_;
  assign new_n22359_ = ~new_n22266_ & new_n22358_;
  assign new_n22360_ = ~new_n22267_ & ~new_n22270_;
  assign new_n22361_ = ~new_n22359_ & ~new_n22360_;
  assign new_n22362_ = \quotient[8]  & ~new_n22361_;
  assign new_n22363_ = ~new_n21591_ & ~new_n22311_;
  assign new_n22364_ = ~new_n22310_ & new_n22363_;
  assign new_n22365_ = ~new_n22362_ & ~new_n22364_;
  assign new_n22366_ = ~\b[50]  & ~new_n22365_;
  assign new_n22367_ = ~new_n21610_ & new_n22265_;
  assign new_n22368_ = ~new_n22261_ & new_n22367_;
  assign new_n22369_ = ~new_n22262_ & ~new_n22265_;
  assign new_n22370_ = ~new_n22368_ & ~new_n22369_;
  assign new_n22371_ = \quotient[8]  & ~new_n22370_;
  assign new_n22372_ = ~new_n21600_ & ~new_n22311_;
  assign new_n22373_ = ~new_n22310_ & new_n22372_;
  assign new_n22374_ = ~new_n22371_ & ~new_n22373_;
  assign new_n22375_ = ~\b[49]  & ~new_n22374_;
  assign new_n22376_ = ~new_n21619_ & new_n22260_;
  assign new_n22377_ = ~new_n22256_ & new_n22376_;
  assign new_n22378_ = ~new_n22257_ & ~new_n22260_;
  assign new_n22379_ = ~new_n22377_ & ~new_n22378_;
  assign new_n22380_ = \quotient[8]  & ~new_n22379_;
  assign new_n22381_ = ~new_n21609_ & ~new_n22311_;
  assign new_n22382_ = ~new_n22310_ & new_n22381_;
  assign new_n22383_ = ~new_n22380_ & ~new_n22382_;
  assign new_n22384_ = ~\b[48]  & ~new_n22383_;
  assign new_n22385_ = ~new_n21628_ & new_n22255_;
  assign new_n22386_ = ~new_n22251_ & new_n22385_;
  assign new_n22387_ = ~new_n22252_ & ~new_n22255_;
  assign new_n22388_ = ~new_n22386_ & ~new_n22387_;
  assign new_n22389_ = \quotient[8]  & ~new_n22388_;
  assign new_n22390_ = ~new_n21618_ & ~new_n22311_;
  assign new_n22391_ = ~new_n22310_ & new_n22390_;
  assign new_n22392_ = ~new_n22389_ & ~new_n22391_;
  assign new_n22393_ = ~\b[47]  & ~new_n22392_;
  assign new_n22394_ = ~new_n21637_ & new_n22250_;
  assign new_n22395_ = ~new_n22246_ & new_n22394_;
  assign new_n22396_ = ~new_n22247_ & ~new_n22250_;
  assign new_n22397_ = ~new_n22395_ & ~new_n22396_;
  assign new_n22398_ = \quotient[8]  & ~new_n22397_;
  assign new_n22399_ = ~new_n21627_ & ~new_n22311_;
  assign new_n22400_ = ~new_n22310_ & new_n22399_;
  assign new_n22401_ = ~new_n22398_ & ~new_n22400_;
  assign new_n22402_ = ~\b[46]  & ~new_n22401_;
  assign new_n22403_ = ~new_n21646_ & new_n22245_;
  assign new_n22404_ = ~new_n22241_ & new_n22403_;
  assign new_n22405_ = ~new_n22242_ & ~new_n22245_;
  assign new_n22406_ = ~new_n22404_ & ~new_n22405_;
  assign new_n22407_ = \quotient[8]  & ~new_n22406_;
  assign new_n22408_ = ~new_n21636_ & ~new_n22311_;
  assign new_n22409_ = ~new_n22310_ & new_n22408_;
  assign new_n22410_ = ~new_n22407_ & ~new_n22409_;
  assign new_n22411_ = ~\b[45]  & ~new_n22410_;
  assign new_n22412_ = ~new_n21655_ & new_n22240_;
  assign new_n22413_ = ~new_n22236_ & new_n22412_;
  assign new_n22414_ = ~new_n22237_ & ~new_n22240_;
  assign new_n22415_ = ~new_n22413_ & ~new_n22414_;
  assign new_n22416_ = \quotient[8]  & ~new_n22415_;
  assign new_n22417_ = ~new_n21645_ & ~new_n22311_;
  assign new_n22418_ = ~new_n22310_ & new_n22417_;
  assign new_n22419_ = ~new_n22416_ & ~new_n22418_;
  assign new_n22420_ = ~\b[44]  & ~new_n22419_;
  assign new_n22421_ = ~new_n21664_ & new_n22235_;
  assign new_n22422_ = ~new_n22231_ & new_n22421_;
  assign new_n22423_ = ~new_n22232_ & ~new_n22235_;
  assign new_n22424_ = ~new_n22422_ & ~new_n22423_;
  assign new_n22425_ = \quotient[8]  & ~new_n22424_;
  assign new_n22426_ = ~new_n21654_ & ~new_n22311_;
  assign new_n22427_ = ~new_n22310_ & new_n22426_;
  assign new_n22428_ = ~new_n22425_ & ~new_n22427_;
  assign new_n22429_ = ~\b[43]  & ~new_n22428_;
  assign new_n22430_ = ~new_n21673_ & new_n22230_;
  assign new_n22431_ = ~new_n22226_ & new_n22430_;
  assign new_n22432_ = ~new_n22227_ & ~new_n22230_;
  assign new_n22433_ = ~new_n22431_ & ~new_n22432_;
  assign new_n22434_ = \quotient[8]  & ~new_n22433_;
  assign new_n22435_ = ~new_n21663_ & ~new_n22311_;
  assign new_n22436_ = ~new_n22310_ & new_n22435_;
  assign new_n22437_ = ~new_n22434_ & ~new_n22436_;
  assign new_n22438_ = ~\b[42]  & ~new_n22437_;
  assign new_n22439_ = ~new_n21682_ & new_n22225_;
  assign new_n22440_ = ~new_n22221_ & new_n22439_;
  assign new_n22441_ = ~new_n22222_ & ~new_n22225_;
  assign new_n22442_ = ~new_n22440_ & ~new_n22441_;
  assign new_n22443_ = \quotient[8]  & ~new_n22442_;
  assign new_n22444_ = ~new_n21672_ & ~new_n22311_;
  assign new_n22445_ = ~new_n22310_ & new_n22444_;
  assign new_n22446_ = ~new_n22443_ & ~new_n22445_;
  assign new_n22447_ = ~\b[41]  & ~new_n22446_;
  assign new_n22448_ = ~new_n21691_ & new_n22220_;
  assign new_n22449_ = ~new_n22216_ & new_n22448_;
  assign new_n22450_ = ~new_n22217_ & ~new_n22220_;
  assign new_n22451_ = ~new_n22449_ & ~new_n22450_;
  assign new_n22452_ = \quotient[8]  & ~new_n22451_;
  assign new_n22453_ = ~new_n21681_ & ~new_n22311_;
  assign new_n22454_ = ~new_n22310_ & new_n22453_;
  assign new_n22455_ = ~new_n22452_ & ~new_n22454_;
  assign new_n22456_ = ~\b[40]  & ~new_n22455_;
  assign new_n22457_ = ~new_n21700_ & new_n22215_;
  assign new_n22458_ = ~new_n22211_ & new_n22457_;
  assign new_n22459_ = ~new_n22212_ & ~new_n22215_;
  assign new_n22460_ = ~new_n22458_ & ~new_n22459_;
  assign new_n22461_ = \quotient[8]  & ~new_n22460_;
  assign new_n22462_ = ~new_n21690_ & ~new_n22311_;
  assign new_n22463_ = ~new_n22310_ & new_n22462_;
  assign new_n22464_ = ~new_n22461_ & ~new_n22463_;
  assign new_n22465_ = ~\b[39]  & ~new_n22464_;
  assign new_n22466_ = ~new_n21709_ & new_n22210_;
  assign new_n22467_ = ~new_n22206_ & new_n22466_;
  assign new_n22468_ = ~new_n22207_ & ~new_n22210_;
  assign new_n22469_ = ~new_n22467_ & ~new_n22468_;
  assign new_n22470_ = \quotient[8]  & ~new_n22469_;
  assign new_n22471_ = ~new_n21699_ & ~new_n22311_;
  assign new_n22472_ = ~new_n22310_ & new_n22471_;
  assign new_n22473_ = ~new_n22470_ & ~new_n22472_;
  assign new_n22474_ = ~\b[38]  & ~new_n22473_;
  assign new_n22475_ = ~new_n21718_ & new_n22205_;
  assign new_n22476_ = ~new_n22201_ & new_n22475_;
  assign new_n22477_ = ~new_n22202_ & ~new_n22205_;
  assign new_n22478_ = ~new_n22476_ & ~new_n22477_;
  assign new_n22479_ = \quotient[8]  & ~new_n22478_;
  assign new_n22480_ = ~new_n21708_ & ~new_n22311_;
  assign new_n22481_ = ~new_n22310_ & new_n22480_;
  assign new_n22482_ = ~new_n22479_ & ~new_n22481_;
  assign new_n22483_ = ~\b[37]  & ~new_n22482_;
  assign new_n22484_ = ~new_n21727_ & new_n22200_;
  assign new_n22485_ = ~new_n22196_ & new_n22484_;
  assign new_n22486_ = ~new_n22197_ & ~new_n22200_;
  assign new_n22487_ = ~new_n22485_ & ~new_n22486_;
  assign new_n22488_ = \quotient[8]  & ~new_n22487_;
  assign new_n22489_ = ~new_n21717_ & ~new_n22311_;
  assign new_n22490_ = ~new_n22310_ & new_n22489_;
  assign new_n22491_ = ~new_n22488_ & ~new_n22490_;
  assign new_n22492_ = ~\b[36]  & ~new_n22491_;
  assign new_n22493_ = ~new_n21736_ & new_n22195_;
  assign new_n22494_ = ~new_n22191_ & new_n22493_;
  assign new_n22495_ = ~new_n22192_ & ~new_n22195_;
  assign new_n22496_ = ~new_n22494_ & ~new_n22495_;
  assign new_n22497_ = \quotient[8]  & ~new_n22496_;
  assign new_n22498_ = ~new_n21726_ & ~new_n22311_;
  assign new_n22499_ = ~new_n22310_ & new_n22498_;
  assign new_n22500_ = ~new_n22497_ & ~new_n22499_;
  assign new_n22501_ = ~\b[35]  & ~new_n22500_;
  assign new_n22502_ = ~new_n21745_ & new_n22190_;
  assign new_n22503_ = ~new_n22186_ & new_n22502_;
  assign new_n22504_ = ~new_n22187_ & ~new_n22190_;
  assign new_n22505_ = ~new_n22503_ & ~new_n22504_;
  assign new_n22506_ = \quotient[8]  & ~new_n22505_;
  assign new_n22507_ = ~new_n21735_ & ~new_n22311_;
  assign new_n22508_ = ~new_n22310_ & new_n22507_;
  assign new_n22509_ = ~new_n22506_ & ~new_n22508_;
  assign new_n22510_ = ~\b[34]  & ~new_n22509_;
  assign new_n22511_ = ~new_n21754_ & new_n22185_;
  assign new_n22512_ = ~new_n22181_ & new_n22511_;
  assign new_n22513_ = ~new_n22182_ & ~new_n22185_;
  assign new_n22514_ = ~new_n22512_ & ~new_n22513_;
  assign new_n22515_ = \quotient[8]  & ~new_n22514_;
  assign new_n22516_ = ~new_n21744_ & ~new_n22311_;
  assign new_n22517_ = ~new_n22310_ & new_n22516_;
  assign new_n22518_ = ~new_n22515_ & ~new_n22517_;
  assign new_n22519_ = ~\b[33]  & ~new_n22518_;
  assign new_n22520_ = ~new_n21763_ & new_n22180_;
  assign new_n22521_ = ~new_n22176_ & new_n22520_;
  assign new_n22522_ = ~new_n22177_ & ~new_n22180_;
  assign new_n22523_ = ~new_n22521_ & ~new_n22522_;
  assign new_n22524_ = \quotient[8]  & ~new_n22523_;
  assign new_n22525_ = ~new_n21753_ & ~new_n22311_;
  assign new_n22526_ = ~new_n22310_ & new_n22525_;
  assign new_n22527_ = ~new_n22524_ & ~new_n22526_;
  assign new_n22528_ = ~\b[32]  & ~new_n22527_;
  assign new_n22529_ = ~new_n21772_ & new_n22175_;
  assign new_n22530_ = ~new_n22171_ & new_n22529_;
  assign new_n22531_ = ~new_n22172_ & ~new_n22175_;
  assign new_n22532_ = ~new_n22530_ & ~new_n22531_;
  assign new_n22533_ = \quotient[8]  & ~new_n22532_;
  assign new_n22534_ = ~new_n21762_ & ~new_n22311_;
  assign new_n22535_ = ~new_n22310_ & new_n22534_;
  assign new_n22536_ = ~new_n22533_ & ~new_n22535_;
  assign new_n22537_ = ~\b[31]  & ~new_n22536_;
  assign new_n22538_ = ~new_n21781_ & new_n22170_;
  assign new_n22539_ = ~new_n22166_ & new_n22538_;
  assign new_n22540_ = ~new_n22167_ & ~new_n22170_;
  assign new_n22541_ = ~new_n22539_ & ~new_n22540_;
  assign new_n22542_ = \quotient[8]  & ~new_n22541_;
  assign new_n22543_ = ~new_n21771_ & ~new_n22311_;
  assign new_n22544_ = ~new_n22310_ & new_n22543_;
  assign new_n22545_ = ~new_n22542_ & ~new_n22544_;
  assign new_n22546_ = ~\b[30]  & ~new_n22545_;
  assign new_n22547_ = ~new_n21790_ & new_n22165_;
  assign new_n22548_ = ~new_n22161_ & new_n22547_;
  assign new_n22549_ = ~new_n22162_ & ~new_n22165_;
  assign new_n22550_ = ~new_n22548_ & ~new_n22549_;
  assign new_n22551_ = \quotient[8]  & ~new_n22550_;
  assign new_n22552_ = ~new_n21780_ & ~new_n22311_;
  assign new_n22553_ = ~new_n22310_ & new_n22552_;
  assign new_n22554_ = ~new_n22551_ & ~new_n22553_;
  assign new_n22555_ = ~\b[29]  & ~new_n22554_;
  assign new_n22556_ = ~new_n21799_ & new_n22160_;
  assign new_n22557_ = ~new_n22156_ & new_n22556_;
  assign new_n22558_ = ~new_n22157_ & ~new_n22160_;
  assign new_n22559_ = ~new_n22557_ & ~new_n22558_;
  assign new_n22560_ = \quotient[8]  & ~new_n22559_;
  assign new_n22561_ = ~new_n21789_ & ~new_n22311_;
  assign new_n22562_ = ~new_n22310_ & new_n22561_;
  assign new_n22563_ = ~new_n22560_ & ~new_n22562_;
  assign new_n22564_ = ~\b[28]  & ~new_n22563_;
  assign new_n22565_ = ~new_n21808_ & new_n22155_;
  assign new_n22566_ = ~new_n22151_ & new_n22565_;
  assign new_n22567_ = ~new_n22152_ & ~new_n22155_;
  assign new_n22568_ = ~new_n22566_ & ~new_n22567_;
  assign new_n22569_ = \quotient[8]  & ~new_n22568_;
  assign new_n22570_ = ~new_n21798_ & ~new_n22311_;
  assign new_n22571_ = ~new_n22310_ & new_n22570_;
  assign new_n22572_ = ~new_n22569_ & ~new_n22571_;
  assign new_n22573_ = ~\b[27]  & ~new_n22572_;
  assign new_n22574_ = ~new_n21817_ & new_n22150_;
  assign new_n22575_ = ~new_n22146_ & new_n22574_;
  assign new_n22576_ = ~new_n22147_ & ~new_n22150_;
  assign new_n22577_ = ~new_n22575_ & ~new_n22576_;
  assign new_n22578_ = \quotient[8]  & ~new_n22577_;
  assign new_n22579_ = ~new_n21807_ & ~new_n22311_;
  assign new_n22580_ = ~new_n22310_ & new_n22579_;
  assign new_n22581_ = ~new_n22578_ & ~new_n22580_;
  assign new_n22582_ = ~\b[26]  & ~new_n22581_;
  assign new_n22583_ = ~new_n21826_ & new_n22145_;
  assign new_n22584_ = ~new_n22141_ & new_n22583_;
  assign new_n22585_ = ~new_n22142_ & ~new_n22145_;
  assign new_n22586_ = ~new_n22584_ & ~new_n22585_;
  assign new_n22587_ = \quotient[8]  & ~new_n22586_;
  assign new_n22588_ = ~new_n21816_ & ~new_n22311_;
  assign new_n22589_ = ~new_n22310_ & new_n22588_;
  assign new_n22590_ = ~new_n22587_ & ~new_n22589_;
  assign new_n22591_ = ~\b[25]  & ~new_n22590_;
  assign new_n22592_ = ~new_n21835_ & new_n22140_;
  assign new_n22593_ = ~new_n22136_ & new_n22592_;
  assign new_n22594_ = ~new_n22137_ & ~new_n22140_;
  assign new_n22595_ = ~new_n22593_ & ~new_n22594_;
  assign new_n22596_ = \quotient[8]  & ~new_n22595_;
  assign new_n22597_ = ~new_n21825_ & ~new_n22311_;
  assign new_n22598_ = ~new_n22310_ & new_n22597_;
  assign new_n22599_ = ~new_n22596_ & ~new_n22598_;
  assign new_n22600_ = ~\b[24]  & ~new_n22599_;
  assign new_n22601_ = ~new_n21844_ & new_n22135_;
  assign new_n22602_ = ~new_n22131_ & new_n22601_;
  assign new_n22603_ = ~new_n22132_ & ~new_n22135_;
  assign new_n22604_ = ~new_n22602_ & ~new_n22603_;
  assign new_n22605_ = \quotient[8]  & ~new_n22604_;
  assign new_n22606_ = ~new_n21834_ & ~new_n22311_;
  assign new_n22607_ = ~new_n22310_ & new_n22606_;
  assign new_n22608_ = ~new_n22605_ & ~new_n22607_;
  assign new_n22609_ = ~\b[23]  & ~new_n22608_;
  assign new_n22610_ = ~new_n21853_ & new_n22130_;
  assign new_n22611_ = ~new_n22126_ & new_n22610_;
  assign new_n22612_ = ~new_n22127_ & ~new_n22130_;
  assign new_n22613_ = ~new_n22611_ & ~new_n22612_;
  assign new_n22614_ = \quotient[8]  & ~new_n22613_;
  assign new_n22615_ = ~new_n21843_ & ~new_n22311_;
  assign new_n22616_ = ~new_n22310_ & new_n22615_;
  assign new_n22617_ = ~new_n22614_ & ~new_n22616_;
  assign new_n22618_ = ~\b[22]  & ~new_n22617_;
  assign new_n22619_ = ~new_n21862_ & new_n22125_;
  assign new_n22620_ = ~new_n22121_ & new_n22619_;
  assign new_n22621_ = ~new_n22122_ & ~new_n22125_;
  assign new_n22622_ = ~new_n22620_ & ~new_n22621_;
  assign new_n22623_ = \quotient[8]  & ~new_n22622_;
  assign new_n22624_ = ~new_n21852_ & ~new_n22311_;
  assign new_n22625_ = ~new_n22310_ & new_n22624_;
  assign new_n22626_ = ~new_n22623_ & ~new_n22625_;
  assign new_n22627_ = ~\b[21]  & ~new_n22626_;
  assign new_n22628_ = ~new_n21871_ & new_n22120_;
  assign new_n22629_ = ~new_n22116_ & new_n22628_;
  assign new_n22630_ = ~new_n22117_ & ~new_n22120_;
  assign new_n22631_ = ~new_n22629_ & ~new_n22630_;
  assign new_n22632_ = \quotient[8]  & ~new_n22631_;
  assign new_n22633_ = ~new_n21861_ & ~new_n22311_;
  assign new_n22634_ = ~new_n22310_ & new_n22633_;
  assign new_n22635_ = ~new_n22632_ & ~new_n22634_;
  assign new_n22636_ = ~\b[20]  & ~new_n22635_;
  assign new_n22637_ = ~new_n21880_ & new_n22115_;
  assign new_n22638_ = ~new_n22111_ & new_n22637_;
  assign new_n22639_ = ~new_n22112_ & ~new_n22115_;
  assign new_n22640_ = ~new_n22638_ & ~new_n22639_;
  assign new_n22641_ = \quotient[8]  & ~new_n22640_;
  assign new_n22642_ = ~new_n21870_ & ~new_n22311_;
  assign new_n22643_ = ~new_n22310_ & new_n22642_;
  assign new_n22644_ = ~new_n22641_ & ~new_n22643_;
  assign new_n22645_ = ~\b[19]  & ~new_n22644_;
  assign new_n22646_ = ~new_n21889_ & new_n22110_;
  assign new_n22647_ = ~new_n22106_ & new_n22646_;
  assign new_n22648_ = ~new_n22107_ & ~new_n22110_;
  assign new_n22649_ = ~new_n22647_ & ~new_n22648_;
  assign new_n22650_ = \quotient[8]  & ~new_n22649_;
  assign new_n22651_ = ~new_n21879_ & ~new_n22311_;
  assign new_n22652_ = ~new_n22310_ & new_n22651_;
  assign new_n22653_ = ~new_n22650_ & ~new_n22652_;
  assign new_n22654_ = ~\b[18]  & ~new_n22653_;
  assign new_n22655_ = ~new_n21898_ & new_n22105_;
  assign new_n22656_ = ~new_n22101_ & new_n22655_;
  assign new_n22657_ = ~new_n22102_ & ~new_n22105_;
  assign new_n22658_ = ~new_n22656_ & ~new_n22657_;
  assign new_n22659_ = \quotient[8]  & ~new_n22658_;
  assign new_n22660_ = ~new_n21888_ & ~new_n22311_;
  assign new_n22661_ = ~new_n22310_ & new_n22660_;
  assign new_n22662_ = ~new_n22659_ & ~new_n22661_;
  assign new_n22663_ = ~\b[17]  & ~new_n22662_;
  assign new_n22664_ = ~new_n21907_ & new_n22100_;
  assign new_n22665_ = ~new_n22096_ & new_n22664_;
  assign new_n22666_ = ~new_n22097_ & ~new_n22100_;
  assign new_n22667_ = ~new_n22665_ & ~new_n22666_;
  assign new_n22668_ = \quotient[8]  & ~new_n22667_;
  assign new_n22669_ = ~new_n21897_ & ~new_n22311_;
  assign new_n22670_ = ~new_n22310_ & new_n22669_;
  assign new_n22671_ = ~new_n22668_ & ~new_n22670_;
  assign new_n22672_ = ~\b[16]  & ~new_n22671_;
  assign new_n22673_ = ~new_n21916_ & new_n22095_;
  assign new_n22674_ = ~new_n22091_ & new_n22673_;
  assign new_n22675_ = ~new_n22092_ & ~new_n22095_;
  assign new_n22676_ = ~new_n22674_ & ~new_n22675_;
  assign new_n22677_ = \quotient[8]  & ~new_n22676_;
  assign new_n22678_ = ~new_n21906_ & ~new_n22311_;
  assign new_n22679_ = ~new_n22310_ & new_n22678_;
  assign new_n22680_ = ~new_n22677_ & ~new_n22679_;
  assign new_n22681_ = ~\b[15]  & ~new_n22680_;
  assign new_n22682_ = ~new_n21925_ & new_n22090_;
  assign new_n22683_ = ~new_n22086_ & new_n22682_;
  assign new_n22684_ = ~new_n22087_ & ~new_n22090_;
  assign new_n22685_ = ~new_n22683_ & ~new_n22684_;
  assign new_n22686_ = \quotient[8]  & ~new_n22685_;
  assign new_n22687_ = ~new_n21915_ & ~new_n22311_;
  assign new_n22688_ = ~new_n22310_ & new_n22687_;
  assign new_n22689_ = ~new_n22686_ & ~new_n22688_;
  assign new_n22690_ = ~\b[14]  & ~new_n22689_;
  assign new_n22691_ = ~new_n21934_ & new_n22085_;
  assign new_n22692_ = ~new_n22081_ & new_n22691_;
  assign new_n22693_ = ~new_n22082_ & ~new_n22085_;
  assign new_n22694_ = ~new_n22692_ & ~new_n22693_;
  assign new_n22695_ = \quotient[8]  & ~new_n22694_;
  assign new_n22696_ = ~new_n21924_ & ~new_n22311_;
  assign new_n22697_ = ~new_n22310_ & new_n22696_;
  assign new_n22698_ = ~new_n22695_ & ~new_n22697_;
  assign new_n22699_ = ~\b[13]  & ~new_n22698_;
  assign new_n22700_ = ~new_n21943_ & new_n22080_;
  assign new_n22701_ = ~new_n22076_ & new_n22700_;
  assign new_n22702_ = ~new_n22077_ & ~new_n22080_;
  assign new_n22703_ = ~new_n22701_ & ~new_n22702_;
  assign new_n22704_ = \quotient[8]  & ~new_n22703_;
  assign new_n22705_ = ~new_n21933_ & ~new_n22311_;
  assign new_n22706_ = ~new_n22310_ & new_n22705_;
  assign new_n22707_ = ~new_n22704_ & ~new_n22706_;
  assign new_n22708_ = ~\b[12]  & ~new_n22707_;
  assign new_n22709_ = ~new_n21952_ & new_n22075_;
  assign new_n22710_ = ~new_n22071_ & new_n22709_;
  assign new_n22711_ = ~new_n22072_ & ~new_n22075_;
  assign new_n22712_ = ~new_n22710_ & ~new_n22711_;
  assign new_n22713_ = \quotient[8]  & ~new_n22712_;
  assign new_n22714_ = ~new_n21942_ & ~new_n22311_;
  assign new_n22715_ = ~new_n22310_ & new_n22714_;
  assign new_n22716_ = ~new_n22713_ & ~new_n22715_;
  assign new_n22717_ = ~\b[11]  & ~new_n22716_;
  assign new_n22718_ = ~new_n21961_ & new_n22070_;
  assign new_n22719_ = ~new_n22066_ & new_n22718_;
  assign new_n22720_ = ~new_n22067_ & ~new_n22070_;
  assign new_n22721_ = ~new_n22719_ & ~new_n22720_;
  assign new_n22722_ = \quotient[8]  & ~new_n22721_;
  assign new_n22723_ = ~new_n21951_ & ~new_n22311_;
  assign new_n22724_ = ~new_n22310_ & new_n22723_;
  assign new_n22725_ = ~new_n22722_ & ~new_n22724_;
  assign new_n22726_ = ~\b[10]  & ~new_n22725_;
  assign new_n22727_ = ~new_n21970_ & new_n22065_;
  assign new_n22728_ = ~new_n22061_ & new_n22727_;
  assign new_n22729_ = ~new_n22062_ & ~new_n22065_;
  assign new_n22730_ = ~new_n22728_ & ~new_n22729_;
  assign new_n22731_ = \quotient[8]  & ~new_n22730_;
  assign new_n22732_ = ~new_n21960_ & ~new_n22311_;
  assign new_n22733_ = ~new_n22310_ & new_n22732_;
  assign new_n22734_ = ~new_n22731_ & ~new_n22733_;
  assign new_n22735_ = ~\b[9]  & ~new_n22734_;
  assign new_n22736_ = ~new_n21979_ & new_n22060_;
  assign new_n22737_ = ~new_n22056_ & new_n22736_;
  assign new_n22738_ = ~new_n22057_ & ~new_n22060_;
  assign new_n22739_ = ~new_n22737_ & ~new_n22738_;
  assign new_n22740_ = \quotient[8]  & ~new_n22739_;
  assign new_n22741_ = ~new_n21969_ & ~new_n22311_;
  assign new_n22742_ = ~new_n22310_ & new_n22741_;
  assign new_n22743_ = ~new_n22740_ & ~new_n22742_;
  assign new_n22744_ = ~\b[8]  & ~new_n22743_;
  assign new_n22745_ = ~new_n21988_ & new_n22055_;
  assign new_n22746_ = ~new_n22051_ & new_n22745_;
  assign new_n22747_ = ~new_n22052_ & ~new_n22055_;
  assign new_n22748_ = ~new_n22746_ & ~new_n22747_;
  assign new_n22749_ = \quotient[8]  & ~new_n22748_;
  assign new_n22750_ = ~new_n21978_ & ~new_n22311_;
  assign new_n22751_ = ~new_n22310_ & new_n22750_;
  assign new_n22752_ = ~new_n22749_ & ~new_n22751_;
  assign new_n22753_ = ~\b[7]  & ~new_n22752_;
  assign new_n22754_ = ~new_n21997_ & new_n22050_;
  assign new_n22755_ = ~new_n22046_ & new_n22754_;
  assign new_n22756_ = ~new_n22047_ & ~new_n22050_;
  assign new_n22757_ = ~new_n22755_ & ~new_n22756_;
  assign new_n22758_ = \quotient[8]  & ~new_n22757_;
  assign new_n22759_ = ~new_n21987_ & ~new_n22311_;
  assign new_n22760_ = ~new_n22310_ & new_n22759_;
  assign new_n22761_ = ~new_n22758_ & ~new_n22760_;
  assign new_n22762_ = ~\b[6]  & ~new_n22761_;
  assign new_n22763_ = ~new_n22006_ & new_n22045_;
  assign new_n22764_ = ~new_n22041_ & new_n22763_;
  assign new_n22765_ = ~new_n22042_ & ~new_n22045_;
  assign new_n22766_ = ~new_n22764_ & ~new_n22765_;
  assign new_n22767_ = \quotient[8]  & ~new_n22766_;
  assign new_n22768_ = ~new_n21996_ & ~new_n22311_;
  assign new_n22769_ = ~new_n22310_ & new_n22768_;
  assign new_n22770_ = ~new_n22767_ & ~new_n22769_;
  assign new_n22771_ = ~\b[5]  & ~new_n22770_;
  assign new_n22772_ = ~new_n22014_ & new_n22040_;
  assign new_n22773_ = ~new_n22036_ & new_n22772_;
  assign new_n22774_ = ~new_n22037_ & ~new_n22040_;
  assign new_n22775_ = ~new_n22773_ & ~new_n22774_;
  assign new_n22776_ = \quotient[8]  & ~new_n22775_;
  assign new_n22777_ = ~new_n22005_ & ~new_n22311_;
  assign new_n22778_ = ~new_n22310_ & new_n22777_;
  assign new_n22779_ = ~new_n22776_ & ~new_n22778_;
  assign new_n22780_ = ~\b[4]  & ~new_n22779_;
  assign new_n22781_ = ~new_n22031_ & new_n22035_;
  assign new_n22782_ = ~new_n22030_ & new_n22781_;
  assign new_n22783_ = ~new_n22032_ & ~new_n22035_;
  assign new_n22784_ = ~new_n22782_ & ~new_n22783_;
  assign new_n22785_ = \quotient[8]  & ~new_n22784_;
  assign new_n22786_ = ~new_n22013_ & ~new_n22311_;
  assign new_n22787_ = ~new_n22310_ & new_n22786_;
  assign new_n22788_ = ~new_n22785_ & ~new_n22787_;
  assign new_n22789_ = ~\b[3]  & ~new_n22788_;
  assign new_n22790_ = ~new_n22027_ & new_n22029_;
  assign new_n22791_ = ~new_n22025_ & new_n22790_;
  assign new_n22792_ = ~new_n22030_ & ~new_n22791_;
  assign new_n22793_ = \quotient[8]  & new_n22792_;
  assign new_n22794_ = ~new_n22024_ & ~new_n22311_;
  assign new_n22795_ = ~new_n22310_ & new_n22794_;
  assign new_n22796_ = ~new_n22793_ & ~new_n22795_;
  assign new_n22797_ = ~\b[2]  & ~new_n22796_;
  assign new_n22798_ = \b[0]  & \quotient[8] ;
  assign new_n22799_ = \a[8]  & ~new_n22798_;
  assign new_n22800_ = new_n22029_ & \quotient[8] ;
  assign new_n22801_ = ~new_n22799_ & ~new_n22800_;
  assign new_n22802_ = \b[1]  & ~new_n22801_;
  assign new_n22803_ = ~\b[1]  & ~new_n22800_;
  assign new_n22804_ = ~new_n22799_ & new_n22803_;
  assign new_n22805_ = ~new_n22802_ & ~new_n22804_;
  assign new_n22806_ = ~\a[7]  & \b[0] ;
  assign new_n22807_ = ~new_n22805_ & ~new_n22806_;
  assign new_n22808_ = ~\b[1]  & ~new_n22801_;
  assign new_n22809_ = ~new_n22807_ & ~new_n22808_;
  assign new_n22810_ = \b[2]  & ~new_n22795_;
  assign new_n22811_ = ~new_n22793_ & new_n22810_;
  assign new_n22812_ = ~new_n22797_ & ~new_n22811_;
  assign new_n22813_ = ~new_n22809_ & new_n22812_;
  assign new_n22814_ = ~new_n22797_ & ~new_n22813_;
  assign new_n22815_ = \b[3]  & ~new_n22787_;
  assign new_n22816_ = ~new_n22785_ & new_n22815_;
  assign new_n22817_ = ~new_n22789_ & ~new_n22816_;
  assign new_n22818_ = ~new_n22814_ & new_n22817_;
  assign new_n22819_ = ~new_n22789_ & ~new_n22818_;
  assign new_n22820_ = \b[4]  & ~new_n22778_;
  assign new_n22821_ = ~new_n22776_ & new_n22820_;
  assign new_n22822_ = ~new_n22780_ & ~new_n22821_;
  assign new_n22823_ = ~new_n22819_ & new_n22822_;
  assign new_n22824_ = ~new_n22780_ & ~new_n22823_;
  assign new_n22825_ = \b[5]  & ~new_n22769_;
  assign new_n22826_ = ~new_n22767_ & new_n22825_;
  assign new_n22827_ = ~new_n22771_ & ~new_n22826_;
  assign new_n22828_ = ~new_n22824_ & new_n22827_;
  assign new_n22829_ = ~new_n22771_ & ~new_n22828_;
  assign new_n22830_ = \b[6]  & ~new_n22760_;
  assign new_n22831_ = ~new_n22758_ & new_n22830_;
  assign new_n22832_ = ~new_n22762_ & ~new_n22831_;
  assign new_n22833_ = ~new_n22829_ & new_n22832_;
  assign new_n22834_ = ~new_n22762_ & ~new_n22833_;
  assign new_n22835_ = \b[7]  & ~new_n22751_;
  assign new_n22836_ = ~new_n22749_ & new_n22835_;
  assign new_n22837_ = ~new_n22753_ & ~new_n22836_;
  assign new_n22838_ = ~new_n22834_ & new_n22837_;
  assign new_n22839_ = ~new_n22753_ & ~new_n22838_;
  assign new_n22840_ = \b[8]  & ~new_n22742_;
  assign new_n22841_ = ~new_n22740_ & new_n22840_;
  assign new_n22842_ = ~new_n22744_ & ~new_n22841_;
  assign new_n22843_ = ~new_n22839_ & new_n22842_;
  assign new_n22844_ = ~new_n22744_ & ~new_n22843_;
  assign new_n22845_ = \b[9]  & ~new_n22733_;
  assign new_n22846_ = ~new_n22731_ & new_n22845_;
  assign new_n22847_ = ~new_n22735_ & ~new_n22846_;
  assign new_n22848_ = ~new_n22844_ & new_n22847_;
  assign new_n22849_ = ~new_n22735_ & ~new_n22848_;
  assign new_n22850_ = \b[10]  & ~new_n22724_;
  assign new_n22851_ = ~new_n22722_ & new_n22850_;
  assign new_n22852_ = ~new_n22726_ & ~new_n22851_;
  assign new_n22853_ = ~new_n22849_ & new_n22852_;
  assign new_n22854_ = ~new_n22726_ & ~new_n22853_;
  assign new_n22855_ = \b[11]  & ~new_n22715_;
  assign new_n22856_ = ~new_n22713_ & new_n22855_;
  assign new_n22857_ = ~new_n22717_ & ~new_n22856_;
  assign new_n22858_ = ~new_n22854_ & new_n22857_;
  assign new_n22859_ = ~new_n22717_ & ~new_n22858_;
  assign new_n22860_ = \b[12]  & ~new_n22706_;
  assign new_n22861_ = ~new_n22704_ & new_n22860_;
  assign new_n22862_ = ~new_n22708_ & ~new_n22861_;
  assign new_n22863_ = ~new_n22859_ & new_n22862_;
  assign new_n22864_ = ~new_n22708_ & ~new_n22863_;
  assign new_n22865_ = \b[13]  & ~new_n22697_;
  assign new_n22866_ = ~new_n22695_ & new_n22865_;
  assign new_n22867_ = ~new_n22699_ & ~new_n22866_;
  assign new_n22868_ = ~new_n22864_ & new_n22867_;
  assign new_n22869_ = ~new_n22699_ & ~new_n22868_;
  assign new_n22870_ = \b[14]  & ~new_n22688_;
  assign new_n22871_ = ~new_n22686_ & new_n22870_;
  assign new_n22872_ = ~new_n22690_ & ~new_n22871_;
  assign new_n22873_ = ~new_n22869_ & new_n22872_;
  assign new_n22874_ = ~new_n22690_ & ~new_n22873_;
  assign new_n22875_ = \b[15]  & ~new_n22679_;
  assign new_n22876_ = ~new_n22677_ & new_n22875_;
  assign new_n22877_ = ~new_n22681_ & ~new_n22876_;
  assign new_n22878_ = ~new_n22874_ & new_n22877_;
  assign new_n22879_ = ~new_n22681_ & ~new_n22878_;
  assign new_n22880_ = \b[16]  & ~new_n22670_;
  assign new_n22881_ = ~new_n22668_ & new_n22880_;
  assign new_n22882_ = ~new_n22672_ & ~new_n22881_;
  assign new_n22883_ = ~new_n22879_ & new_n22882_;
  assign new_n22884_ = ~new_n22672_ & ~new_n22883_;
  assign new_n22885_ = \b[17]  & ~new_n22661_;
  assign new_n22886_ = ~new_n22659_ & new_n22885_;
  assign new_n22887_ = ~new_n22663_ & ~new_n22886_;
  assign new_n22888_ = ~new_n22884_ & new_n22887_;
  assign new_n22889_ = ~new_n22663_ & ~new_n22888_;
  assign new_n22890_ = \b[18]  & ~new_n22652_;
  assign new_n22891_ = ~new_n22650_ & new_n22890_;
  assign new_n22892_ = ~new_n22654_ & ~new_n22891_;
  assign new_n22893_ = ~new_n22889_ & new_n22892_;
  assign new_n22894_ = ~new_n22654_ & ~new_n22893_;
  assign new_n22895_ = \b[19]  & ~new_n22643_;
  assign new_n22896_ = ~new_n22641_ & new_n22895_;
  assign new_n22897_ = ~new_n22645_ & ~new_n22896_;
  assign new_n22898_ = ~new_n22894_ & new_n22897_;
  assign new_n22899_ = ~new_n22645_ & ~new_n22898_;
  assign new_n22900_ = \b[20]  & ~new_n22634_;
  assign new_n22901_ = ~new_n22632_ & new_n22900_;
  assign new_n22902_ = ~new_n22636_ & ~new_n22901_;
  assign new_n22903_ = ~new_n22899_ & new_n22902_;
  assign new_n22904_ = ~new_n22636_ & ~new_n22903_;
  assign new_n22905_ = \b[21]  & ~new_n22625_;
  assign new_n22906_ = ~new_n22623_ & new_n22905_;
  assign new_n22907_ = ~new_n22627_ & ~new_n22906_;
  assign new_n22908_ = ~new_n22904_ & new_n22907_;
  assign new_n22909_ = ~new_n22627_ & ~new_n22908_;
  assign new_n22910_ = \b[22]  & ~new_n22616_;
  assign new_n22911_ = ~new_n22614_ & new_n22910_;
  assign new_n22912_ = ~new_n22618_ & ~new_n22911_;
  assign new_n22913_ = ~new_n22909_ & new_n22912_;
  assign new_n22914_ = ~new_n22618_ & ~new_n22913_;
  assign new_n22915_ = \b[23]  & ~new_n22607_;
  assign new_n22916_ = ~new_n22605_ & new_n22915_;
  assign new_n22917_ = ~new_n22609_ & ~new_n22916_;
  assign new_n22918_ = ~new_n22914_ & new_n22917_;
  assign new_n22919_ = ~new_n22609_ & ~new_n22918_;
  assign new_n22920_ = \b[24]  & ~new_n22598_;
  assign new_n22921_ = ~new_n22596_ & new_n22920_;
  assign new_n22922_ = ~new_n22600_ & ~new_n22921_;
  assign new_n22923_ = ~new_n22919_ & new_n22922_;
  assign new_n22924_ = ~new_n22600_ & ~new_n22923_;
  assign new_n22925_ = \b[25]  & ~new_n22589_;
  assign new_n22926_ = ~new_n22587_ & new_n22925_;
  assign new_n22927_ = ~new_n22591_ & ~new_n22926_;
  assign new_n22928_ = ~new_n22924_ & new_n22927_;
  assign new_n22929_ = ~new_n22591_ & ~new_n22928_;
  assign new_n22930_ = \b[26]  & ~new_n22580_;
  assign new_n22931_ = ~new_n22578_ & new_n22930_;
  assign new_n22932_ = ~new_n22582_ & ~new_n22931_;
  assign new_n22933_ = ~new_n22929_ & new_n22932_;
  assign new_n22934_ = ~new_n22582_ & ~new_n22933_;
  assign new_n22935_ = \b[27]  & ~new_n22571_;
  assign new_n22936_ = ~new_n22569_ & new_n22935_;
  assign new_n22937_ = ~new_n22573_ & ~new_n22936_;
  assign new_n22938_ = ~new_n22934_ & new_n22937_;
  assign new_n22939_ = ~new_n22573_ & ~new_n22938_;
  assign new_n22940_ = \b[28]  & ~new_n22562_;
  assign new_n22941_ = ~new_n22560_ & new_n22940_;
  assign new_n22942_ = ~new_n22564_ & ~new_n22941_;
  assign new_n22943_ = ~new_n22939_ & new_n22942_;
  assign new_n22944_ = ~new_n22564_ & ~new_n22943_;
  assign new_n22945_ = \b[29]  & ~new_n22553_;
  assign new_n22946_ = ~new_n22551_ & new_n22945_;
  assign new_n22947_ = ~new_n22555_ & ~new_n22946_;
  assign new_n22948_ = ~new_n22944_ & new_n22947_;
  assign new_n22949_ = ~new_n22555_ & ~new_n22948_;
  assign new_n22950_ = \b[30]  & ~new_n22544_;
  assign new_n22951_ = ~new_n22542_ & new_n22950_;
  assign new_n22952_ = ~new_n22546_ & ~new_n22951_;
  assign new_n22953_ = ~new_n22949_ & new_n22952_;
  assign new_n22954_ = ~new_n22546_ & ~new_n22953_;
  assign new_n22955_ = \b[31]  & ~new_n22535_;
  assign new_n22956_ = ~new_n22533_ & new_n22955_;
  assign new_n22957_ = ~new_n22537_ & ~new_n22956_;
  assign new_n22958_ = ~new_n22954_ & new_n22957_;
  assign new_n22959_ = ~new_n22537_ & ~new_n22958_;
  assign new_n22960_ = \b[32]  & ~new_n22526_;
  assign new_n22961_ = ~new_n22524_ & new_n22960_;
  assign new_n22962_ = ~new_n22528_ & ~new_n22961_;
  assign new_n22963_ = ~new_n22959_ & new_n22962_;
  assign new_n22964_ = ~new_n22528_ & ~new_n22963_;
  assign new_n22965_ = \b[33]  & ~new_n22517_;
  assign new_n22966_ = ~new_n22515_ & new_n22965_;
  assign new_n22967_ = ~new_n22519_ & ~new_n22966_;
  assign new_n22968_ = ~new_n22964_ & new_n22967_;
  assign new_n22969_ = ~new_n22519_ & ~new_n22968_;
  assign new_n22970_ = \b[34]  & ~new_n22508_;
  assign new_n22971_ = ~new_n22506_ & new_n22970_;
  assign new_n22972_ = ~new_n22510_ & ~new_n22971_;
  assign new_n22973_ = ~new_n22969_ & new_n22972_;
  assign new_n22974_ = ~new_n22510_ & ~new_n22973_;
  assign new_n22975_ = \b[35]  & ~new_n22499_;
  assign new_n22976_ = ~new_n22497_ & new_n22975_;
  assign new_n22977_ = ~new_n22501_ & ~new_n22976_;
  assign new_n22978_ = ~new_n22974_ & new_n22977_;
  assign new_n22979_ = ~new_n22501_ & ~new_n22978_;
  assign new_n22980_ = \b[36]  & ~new_n22490_;
  assign new_n22981_ = ~new_n22488_ & new_n22980_;
  assign new_n22982_ = ~new_n22492_ & ~new_n22981_;
  assign new_n22983_ = ~new_n22979_ & new_n22982_;
  assign new_n22984_ = ~new_n22492_ & ~new_n22983_;
  assign new_n22985_ = \b[37]  & ~new_n22481_;
  assign new_n22986_ = ~new_n22479_ & new_n22985_;
  assign new_n22987_ = ~new_n22483_ & ~new_n22986_;
  assign new_n22988_ = ~new_n22984_ & new_n22987_;
  assign new_n22989_ = ~new_n22483_ & ~new_n22988_;
  assign new_n22990_ = \b[38]  & ~new_n22472_;
  assign new_n22991_ = ~new_n22470_ & new_n22990_;
  assign new_n22992_ = ~new_n22474_ & ~new_n22991_;
  assign new_n22993_ = ~new_n22989_ & new_n22992_;
  assign new_n22994_ = ~new_n22474_ & ~new_n22993_;
  assign new_n22995_ = \b[39]  & ~new_n22463_;
  assign new_n22996_ = ~new_n22461_ & new_n22995_;
  assign new_n22997_ = ~new_n22465_ & ~new_n22996_;
  assign new_n22998_ = ~new_n22994_ & new_n22997_;
  assign new_n22999_ = ~new_n22465_ & ~new_n22998_;
  assign new_n23000_ = \b[40]  & ~new_n22454_;
  assign new_n23001_ = ~new_n22452_ & new_n23000_;
  assign new_n23002_ = ~new_n22456_ & ~new_n23001_;
  assign new_n23003_ = ~new_n22999_ & new_n23002_;
  assign new_n23004_ = ~new_n22456_ & ~new_n23003_;
  assign new_n23005_ = \b[41]  & ~new_n22445_;
  assign new_n23006_ = ~new_n22443_ & new_n23005_;
  assign new_n23007_ = ~new_n22447_ & ~new_n23006_;
  assign new_n23008_ = ~new_n23004_ & new_n23007_;
  assign new_n23009_ = ~new_n22447_ & ~new_n23008_;
  assign new_n23010_ = \b[42]  & ~new_n22436_;
  assign new_n23011_ = ~new_n22434_ & new_n23010_;
  assign new_n23012_ = ~new_n22438_ & ~new_n23011_;
  assign new_n23013_ = ~new_n23009_ & new_n23012_;
  assign new_n23014_ = ~new_n22438_ & ~new_n23013_;
  assign new_n23015_ = \b[43]  & ~new_n22427_;
  assign new_n23016_ = ~new_n22425_ & new_n23015_;
  assign new_n23017_ = ~new_n22429_ & ~new_n23016_;
  assign new_n23018_ = ~new_n23014_ & new_n23017_;
  assign new_n23019_ = ~new_n22429_ & ~new_n23018_;
  assign new_n23020_ = \b[44]  & ~new_n22418_;
  assign new_n23021_ = ~new_n22416_ & new_n23020_;
  assign new_n23022_ = ~new_n22420_ & ~new_n23021_;
  assign new_n23023_ = ~new_n23019_ & new_n23022_;
  assign new_n23024_ = ~new_n22420_ & ~new_n23023_;
  assign new_n23025_ = \b[45]  & ~new_n22409_;
  assign new_n23026_ = ~new_n22407_ & new_n23025_;
  assign new_n23027_ = ~new_n22411_ & ~new_n23026_;
  assign new_n23028_ = ~new_n23024_ & new_n23027_;
  assign new_n23029_ = ~new_n22411_ & ~new_n23028_;
  assign new_n23030_ = \b[46]  & ~new_n22400_;
  assign new_n23031_ = ~new_n22398_ & new_n23030_;
  assign new_n23032_ = ~new_n22402_ & ~new_n23031_;
  assign new_n23033_ = ~new_n23029_ & new_n23032_;
  assign new_n23034_ = ~new_n22402_ & ~new_n23033_;
  assign new_n23035_ = \b[47]  & ~new_n22391_;
  assign new_n23036_ = ~new_n22389_ & new_n23035_;
  assign new_n23037_ = ~new_n22393_ & ~new_n23036_;
  assign new_n23038_ = ~new_n23034_ & new_n23037_;
  assign new_n23039_ = ~new_n22393_ & ~new_n23038_;
  assign new_n23040_ = \b[48]  & ~new_n22382_;
  assign new_n23041_ = ~new_n22380_ & new_n23040_;
  assign new_n23042_ = ~new_n22384_ & ~new_n23041_;
  assign new_n23043_ = ~new_n23039_ & new_n23042_;
  assign new_n23044_ = ~new_n22384_ & ~new_n23043_;
  assign new_n23045_ = \b[49]  & ~new_n22373_;
  assign new_n23046_ = ~new_n22371_ & new_n23045_;
  assign new_n23047_ = ~new_n22375_ & ~new_n23046_;
  assign new_n23048_ = ~new_n23044_ & new_n23047_;
  assign new_n23049_ = ~new_n22375_ & ~new_n23048_;
  assign new_n23050_ = \b[50]  & ~new_n22364_;
  assign new_n23051_ = ~new_n22362_ & new_n23050_;
  assign new_n23052_ = ~new_n22366_ & ~new_n23051_;
  assign new_n23053_ = ~new_n23049_ & new_n23052_;
  assign new_n23054_ = ~new_n22366_ & ~new_n23053_;
  assign new_n23055_ = \b[51]  & ~new_n22355_;
  assign new_n23056_ = ~new_n22353_ & new_n23055_;
  assign new_n23057_ = ~new_n22357_ & ~new_n23056_;
  assign new_n23058_ = ~new_n23054_ & new_n23057_;
  assign new_n23059_ = ~new_n22357_ & ~new_n23058_;
  assign new_n23060_ = \b[52]  & ~new_n22346_;
  assign new_n23061_ = ~new_n22344_ & new_n23060_;
  assign new_n23062_ = ~new_n22348_ & ~new_n23061_;
  assign new_n23063_ = ~new_n23059_ & new_n23062_;
  assign new_n23064_ = ~new_n22348_ & ~new_n23063_;
  assign new_n23065_ = \b[53]  & ~new_n22337_;
  assign new_n23066_ = ~new_n22335_ & new_n23065_;
  assign new_n23067_ = ~new_n22339_ & ~new_n23066_;
  assign new_n23068_ = ~new_n23064_ & new_n23067_;
  assign new_n23069_ = ~new_n22339_ & ~new_n23068_;
  assign new_n23070_ = \b[54]  & ~new_n22328_;
  assign new_n23071_ = ~new_n22326_ & new_n23070_;
  assign new_n23072_ = ~new_n22330_ & ~new_n23071_;
  assign new_n23073_ = ~new_n23069_ & new_n23072_;
  assign new_n23074_ = ~new_n22330_ & ~new_n23073_;
  assign new_n23075_ = \b[55]  & ~new_n22319_;
  assign new_n23076_ = ~new_n22317_ & new_n23075_;
  assign new_n23077_ = ~new_n22321_ & ~new_n23076_;
  assign new_n23078_ = ~new_n23074_ & new_n23077_;
  assign new_n23079_ = ~new_n22321_ & ~new_n23078_;
  assign new_n23080_ = ~new_n21547_ & ~new_n22307_;
  assign new_n23081_ = ~new_n22305_ & new_n23080_;
  assign new_n23082_ = ~new_n22296_ & new_n23081_;
  assign new_n23083_ = ~new_n22305_ & ~new_n22307_;
  assign new_n23084_ = ~new_n22297_ & ~new_n23083_;
  assign new_n23085_ = ~new_n23082_ & ~new_n23084_;
  assign new_n23086_ = \quotient[8]  & ~new_n23085_;
  assign new_n23087_ = ~new_n22304_ & ~new_n22311_;
  assign new_n23088_ = ~new_n22310_ & new_n23087_;
  assign new_n23089_ = ~new_n23086_ & ~new_n23088_;
  assign new_n23090_ = ~\b[56]  & ~new_n23089_;
  assign new_n23091_ = \b[56]  & ~new_n23088_;
  assign new_n23092_ = ~new_n23086_ & new_n23091_;
  assign new_n23093_ = new_n407_ & ~new_n23092_;
  assign new_n23094_ = ~new_n23090_ & new_n23093_;
  assign new_n23095_ = ~new_n23079_ & new_n23094_;
  assign new_n23096_ = new_n337_ & ~new_n23089_;
  assign \quotient[7]  = new_n23095_ | new_n23096_;
  assign new_n23098_ = ~new_n22330_ & new_n23077_;
  assign new_n23099_ = ~new_n23073_ & new_n23098_;
  assign new_n23100_ = ~new_n23074_ & ~new_n23077_;
  assign new_n23101_ = ~new_n23099_ & ~new_n23100_;
  assign new_n23102_ = \quotient[7]  & ~new_n23101_;
  assign new_n23103_ = ~new_n22320_ & ~new_n23096_;
  assign new_n23104_ = ~new_n23095_ & new_n23103_;
  assign new_n23105_ = ~new_n23102_ & ~new_n23104_;
  assign new_n23106_ = ~new_n22321_ & ~new_n23092_;
  assign new_n23107_ = ~new_n23090_ & new_n23106_;
  assign new_n23108_ = ~new_n23078_ & new_n23107_;
  assign new_n23109_ = ~new_n23090_ & ~new_n23092_;
  assign new_n23110_ = ~new_n23079_ & ~new_n23109_;
  assign new_n23111_ = ~new_n23108_ & ~new_n23110_;
  assign new_n23112_ = \quotient[7]  & ~new_n23111_;
  assign new_n23113_ = ~new_n23089_ & ~new_n23096_;
  assign new_n23114_ = ~new_n23095_ & new_n23113_;
  assign new_n23115_ = ~new_n23112_ & ~new_n23114_;
  assign new_n23116_ = ~\b[57]  & ~new_n23115_;
  assign new_n23117_ = ~\b[56]  & ~new_n23105_;
  assign new_n23118_ = ~new_n22339_ & new_n23072_;
  assign new_n23119_ = ~new_n23068_ & new_n23118_;
  assign new_n23120_ = ~new_n23069_ & ~new_n23072_;
  assign new_n23121_ = ~new_n23119_ & ~new_n23120_;
  assign new_n23122_ = \quotient[7]  & ~new_n23121_;
  assign new_n23123_ = ~new_n22329_ & ~new_n23096_;
  assign new_n23124_ = ~new_n23095_ & new_n23123_;
  assign new_n23125_ = ~new_n23122_ & ~new_n23124_;
  assign new_n23126_ = ~\b[55]  & ~new_n23125_;
  assign new_n23127_ = ~new_n22348_ & new_n23067_;
  assign new_n23128_ = ~new_n23063_ & new_n23127_;
  assign new_n23129_ = ~new_n23064_ & ~new_n23067_;
  assign new_n23130_ = ~new_n23128_ & ~new_n23129_;
  assign new_n23131_ = \quotient[7]  & ~new_n23130_;
  assign new_n23132_ = ~new_n22338_ & ~new_n23096_;
  assign new_n23133_ = ~new_n23095_ & new_n23132_;
  assign new_n23134_ = ~new_n23131_ & ~new_n23133_;
  assign new_n23135_ = ~\b[54]  & ~new_n23134_;
  assign new_n23136_ = ~new_n22357_ & new_n23062_;
  assign new_n23137_ = ~new_n23058_ & new_n23136_;
  assign new_n23138_ = ~new_n23059_ & ~new_n23062_;
  assign new_n23139_ = ~new_n23137_ & ~new_n23138_;
  assign new_n23140_ = \quotient[7]  & ~new_n23139_;
  assign new_n23141_ = ~new_n22347_ & ~new_n23096_;
  assign new_n23142_ = ~new_n23095_ & new_n23141_;
  assign new_n23143_ = ~new_n23140_ & ~new_n23142_;
  assign new_n23144_ = ~\b[53]  & ~new_n23143_;
  assign new_n23145_ = ~new_n22366_ & new_n23057_;
  assign new_n23146_ = ~new_n23053_ & new_n23145_;
  assign new_n23147_ = ~new_n23054_ & ~new_n23057_;
  assign new_n23148_ = ~new_n23146_ & ~new_n23147_;
  assign new_n23149_ = \quotient[7]  & ~new_n23148_;
  assign new_n23150_ = ~new_n22356_ & ~new_n23096_;
  assign new_n23151_ = ~new_n23095_ & new_n23150_;
  assign new_n23152_ = ~new_n23149_ & ~new_n23151_;
  assign new_n23153_ = ~\b[52]  & ~new_n23152_;
  assign new_n23154_ = ~new_n22375_ & new_n23052_;
  assign new_n23155_ = ~new_n23048_ & new_n23154_;
  assign new_n23156_ = ~new_n23049_ & ~new_n23052_;
  assign new_n23157_ = ~new_n23155_ & ~new_n23156_;
  assign new_n23158_ = \quotient[7]  & ~new_n23157_;
  assign new_n23159_ = ~new_n22365_ & ~new_n23096_;
  assign new_n23160_ = ~new_n23095_ & new_n23159_;
  assign new_n23161_ = ~new_n23158_ & ~new_n23160_;
  assign new_n23162_ = ~\b[51]  & ~new_n23161_;
  assign new_n23163_ = ~new_n22384_ & new_n23047_;
  assign new_n23164_ = ~new_n23043_ & new_n23163_;
  assign new_n23165_ = ~new_n23044_ & ~new_n23047_;
  assign new_n23166_ = ~new_n23164_ & ~new_n23165_;
  assign new_n23167_ = \quotient[7]  & ~new_n23166_;
  assign new_n23168_ = ~new_n22374_ & ~new_n23096_;
  assign new_n23169_ = ~new_n23095_ & new_n23168_;
  assign new_n23170_ = ~new_n23167_ & ~new_n23169_;
  assign new_n23171_ = ~\b[50]  & ~new_n23170_;
  assign new_n23172_ = ~new_n22393_ & new_n23042_;
  assign new_n23173_ = ~new_n23038_ & new_n23172_;
  assign new_n23174_ = ~new_n23039_ & ~new_n23042_;
  assign new_n23175_ = ~new_n23173_ & ~new_n23174_;
  assign new_n23176_ = \quotient[7]  & ~new_n23175_;
  assign new_n23177_ = ~new_n22383_ & ~new_n23096_;
  assign new_n23178_ = ~new_n23095_ & new_n23177_;
  assign new_n23179_ = ~new_n23176_ & ~new_n23178_;
  assign new_n23180_ = ~\b[49]  & ~new_n23179_;
  assign new_n23181_ = ~new_n22402_ & new_n23037_;
  assign new_n23182_ = ~new_n23033_ & new_n23181_;
  assign new_n23183_ = ~new_n23034_ & ~new_n23037_;
  assign new_n23184_ = ~new_n23182_ & ~new_n23183_;
  assign new_n23185_ = \quotient[7]  & ~new_n23184_;
  assign new_n23186_ = ~new_n22392_ & ~new_n23096_;
  assign new_n23187_ = ~new_n23095_ & new_n23186_;
  assign new_n23188_ = ~new_n23185_ & ~new_n23187_;
  assign new_n23189_ = ~\b[48]  & ~new_n23188_;
  assign new_n23190_ = ~new_n22411_ & new_n23032_;
  assign new_n23191_ = ~new_n23028_ & new_n23190_;
  assign new_n23192_ = ~new_n23029_ & ~new_n23032_;
  assign new_n23193_ = ~new_n23191_ & ~new_n23192_;
  assign new_n23194_ = \quotient[7]  & ~new_n23193_;
  assign new_n23195_ = ~new_n22401_ & ~new_n23096_;
  assign new_n23196_ = ~new_n23095_ & new_n23195_;
  assign new_n23197_ = ~new_n23194_ & ~new_n23196_;
  assign new_n23198_ = ~\b[47]  & ~new_n23197_;
  assign new_n23199_ = ~new_n22420_ & new_n23027_;
  assign new_n23200_ = ~new_n23023_ & new_n23199_;
  assign new_n23201_ = ~new_n23024_ & ~new_n23027_;
  assign new_n23202_ = ~new_n23200_ & ~new_n23201_;
  assign new_n23203_ = \quotient[7]  & ~new_n23202_;
  assign new_n23204_ = ~new_n22410_ & ~new_n23096_;
  assign new_n23205_ = ~new_n23095_ & new_n23204_;
  assign new_n23206_ = ~new_n23203_ & ~new_n23205_;
  assign new_n23207_ = ~\b[46]  & ~new_n23206_;
  assign new_n23208_ = ~new_n22429_ & new_n23022_;
  assign new_n23209_ = ~new_n23018_ & new_n23208_;
  assign new_n23210_ = ~new_n23019_ & ~new_n23022_;
  assign new_n23211_ = ~new_n23209_ & ~new_n23210_;
  assign new_n23212_ = \quotient[7]  & ~new_n23211_;
  assign new_n23213_ = ~new_n22419_ & ~new_n23096_;
  assign new_n23214_ = ~new_n23095_ & new_n23213_;
  assign new_n23215_ = ~new_n23212_ & ~new_n23214_;
  assign new_n23216_ = ~\b[45]  & ~new_n23215_;
  assign new_n23217_ = ~new_n22438_ & new_n23017_;
  assign new_n23218_ = ~new_n23013_ & new_n23217_;
  assign new_n23219_ = ~new_n23014_ & ~new_n23017_;
  assign new_n23220_ = ~new_n23218_ & ~new_n23219_;
  assign new_n23221_ = \quotient[7]  & ~new_n23220_;
  assign new_n23222_ = ~new_n22428_ & ~new_n23096_;
  assign new_n23223_ = ~new_n23095_ & new_n23222_;
  assign new_n23224_ = ~new_n23221_ & ~new_n23223_;
  assign new_n23225_ = ~\b[44]  & ~new_n23224_;
  assign new_n23226_ = ~new_n22447_ & new_n23012_;
  assign new_n23227_ = ~new_n23008_ & new_n23226_;
  assign new_n23228_ = ~new_n23009_ & ~new_n23012_;
  assign new_n23229_ = ~new_n23227_ & ~new_n23228_;
  assign new_n23230_ = \quotient[7]  & ~new_n23229_;
  assign new_n23231_ = ~new_n22437_ & ~new_n23096_;
  assign new_n23232_ = ~new_n23095_ & new_n23231_;
  assign new_n23233_ = ~new_n23230_ & ~new_n23232_;
  assign new_n23234_ = ~\b[43]  & ~new_n23233_;
  assign new_n23235_ = ~new_n22456_ & new_n23007_;
  assign new_n23236_ = ~new_n23003_ & new_n23235_;
  assign new_n23237_ = ~new_n23004_ & ~new_n23007_;
  assign new_n23238_ = ~new_n23236_ & ~new_n23237_;
  assign new_n23239_ = \quotient[7]  & ~new_n23238_;
  assign new_n23240_ = ~new_n22446_ & ~new_n23096_;
  assign new_n23241_ = ~new_n23095_ & new_n23240_;
  assign new_n23242_ = ~new_n23239_ & ~new_n23241_;
  assign new_n23243_ = ~\b[42]  & ~new_n23242_;
  assign new_n23244_ = ~new_n22465_ & new_n23002_;
  assign new_n23245_ = ~new_n22998_ & new_n23244_;
  assign new_n23246_ = ~new_n22999_ & ~new_n23002_;
  assign new_n23247_ = ~new_n23245_ & ~new_n23246_;
  assign new_n23248_ = \quotient[7]  & ~new_n23247_;
  assign new_n23249_ = ~new_n22455_ & ~new_n23096_;
  assign new_n23250_ = ~new_n23095_ & new_n23249_;
  assign new_n23251_ = ~new_n23248_ & ~new_n23250_;
  assign new_n23252_ = ~\b[41]  & ~new_n23251_;
  assign new_n23253_ = ~new_n22474_ & new_n22997_;
  assign new_n23254_ = ~new_n22993_ & new_n23253_;
  assign new_n23255_ = ~new_n22994_ & ~new_n22997_;
  assign new_n23256_ = ~new_n23254_ & ~new_n23255_;
  assign new_n23257_ = \quotient[7]  & ~new_n23256_;
  assign new_n23258_ = ~new_n22464_ & ~new_n23096_;
  assign new_n23259_ = ~new_n23095_ & new_n23258_;
  assign new_n23260_ = ~new_n23257_ & ~new_n23259_;
  assign new_n23261_ = ~\b[40]  & ~new_n23260_;
  assign new_n23262_ = ~new_n22483_ & new_n22992_;
  assign new_n23263_ = ~new_n22988_ & new_n23262_;
  assign new_n23264_ = ~new_n22989_ & ~new_n22992_;
  assign new_n23265_ = ~new_n23263_ & ~new_n23264_;
  assign new_n23266_ = \quotient[7]  & ~new_n23265_;
  assign new_n23267_ = ~new_n22473_ & ~new_n23096_;
  assign new_n23268_ = ~new_n23095_ & new_n23267_;
  assign new_n23269_ = ~new_n23266_ & ~new_n23268_;
  assign new_n23270_ = ~\b[39]  & ~new_n23269_;
  assign new_n23271_ = ~new_n22492_ & new_n22987_;
  assign new_n23272_ = ~new_n22983_ & new_n23271_;
  assign new_n23273_ = ~new_n22984_ & ~new_n22987_;
  assign new_n23274_ = ~new_n23272_ & ~new_n23273_;
  assign new_n23275_ = \quotient[7]  & ~new_n23274_;
  assign new_n23276_ = ~new_n22482_ & ~new_n23096_;
  assign new_n23277_ = ~new_n23095_ & new_n23276_;
  assign new_n23278_ = ~new_n23275_ & ~new_n23277_;
  assign new_n23279_ = ~\b[38]  & ~new_n23278_;
  assign new_n23280_ = ~new_n22501_ & new_n22982_;
  assign new_n23281_ = ~new_n22978_ & new_n23280_;
  assign new_n23282_ = ~new_n22979_ & ~new_n22982_;
  assign new_n23283_ = ~new_n23281_ & ~new_n23282_;
  assign new_n23284_ = \quotient[7]  & ~new_n23283_;
  assign new_n23285_ = ~new_n22491_ & ~new_n23096_;
  assign new_n23286_ = ~new_n23095_ & new_n23285_;
  assign new_n23287_ = ~new_n23284_ & ~new_n23286_;
  assign new_n23288_ = ~\b[37]  & ~new_n23287_;
  assign new_n23289_ = ~new_n22510_ & new_n22977_;
  assign new_n23290_ = ~new_n22973_ & new_n23289_;
  assign new_n23291_ = ~new_n22974_ & ~new_n22977_;
  assign new_n23292_ = ~new_n23290_ & ~new_n23291_;
  assign new_n23293_ = \quotient[7]  & ~new_n23292_;
  assign new_n23294_ = ~new_n22500_ & ~new_n23096_;
  assign new_n23295_ = ~new_n23095_ & new_n23294_;
  assign new_n23296_ = ~new_n23293_ & ~new_n23295_;
  assign new_n23297_ = ~\b[36]  & ~new_n23296_;
  assign new_n23298_ = ~new_n22519_ & new_n22972_;
  assign new_n23299_ = ~new_n22968_ & new_n23298_;
  assign new_n23300_ = ~new_n22969_ & ~new_n22972_;
  assign new_n23301_ = ~new_n23299_ & ~new_n23300_;
  assign new_n23302_ = \quotient[7]  & ~new_n23301_;
  assign new_n23303_ = ~new_n22509_ & ~new_n23096_;
  assign new_n23304_ = ~new_n23095_ & new_n23303_;
  assign new_n23305_ = ~new_n23302_ & ~new_n23304_;
  assign new_n23306_ = ~\b[35]  & ~new_n23305_;
  assign new_n23307_ = ~new_n22528_ & new_n22967_;
  assign new_n23308_ = ~new_n22963_ & new_n23307_;
  assign new_n23309_ = ~new_n22964_ & ~new_n22967_;
  assign new_n23310_ = ~new_n23308_ & ~new_n23309_;
  assign new_n23311_ = \quotient[7]  & ~new_n23310_;
  assign new_n23312_ = ~new_n22518_ & ~new_n23096_;
  assign new_n23313_ = ~new_n23095_ & new_n23312_;
  assign new_n23314_ = ~new_n23311_ & ~new_n23313_;
  assign new_n23315_ = ~\b[34]  & ~new_n23314_;
  assign new_n23316_ = ~new_n22537_ & new_n22962_;
  assign new_n23317_ = ~new_n22958_ & new_n23316_;
  assign new_n23318_ = ~new_n22959_ & ~new_n22962_;
  assign new_n23319_ = ~new_n23317_ & ~new_n23318_;
  assign new_n23320_ = \quotient[7]  & ~new_n23319_;
  assign new_n23321_ = ~new_n22527_ & ~new_n23096_;
  assign new_n23322_ = ~new_n23095_ & new_n23321_;
  assign new_n23323_ = ~new_n23320_ & ~new_n23322_;
  assign new_n23324_ = ~\b[33]  & ~new_n23323_;
  assign new_n23325_ = ~new_n22546_ & new_n22957_;
  assign new_n23326_ = ~new_n22953_ & new_n23325_;
  assign new_n23327_ = ~new_n22954_ & ~new_n22957_;
  assign new_n23328_ = ~new_n23326_ & ~new_n23327_;
  assign new_n23329_ = \quotient[7]  & ~new_n23328_;
  assign new_n23330_ = ~new_n22536_ & ~new_n23096_;
  assign new_n23331_ = ~new_n23095_ & new_n23330_;
  assign new_n23332_ = ~new_n23329_ & ~new_n23331_;
  assign new_n23333_ = ~\b[32]  & ~new_n23332_;
  assign new_n23334_ = ~new_n22555_ & new_n22952_;
  assign new_n23335_ = ~new_n22948_ & new_n23334_;
  assign new_n23336_ = ~new_n22949_ & ~new_n22952_;
  assign new_n23337_ = ~new_n23335_ & ~new_n23336_;
  assign new_n23338_ = \quotient[7]  & ~new_n23337_;
  assign new_n23339_ = ~new_n22545_ & ~new_n23096_;
  assign new_n23340_ = ~new_n23095_ & new_n23339_;
  assign new_n23341_ = ~new_n23338_ & ~new_n23340_;
  assign new_n23342_ = ~\b[31]  & ~new_n23341_;
  assign new_n23343_ = ~new_n22564_ & new_n22947_;
  assign new_n23344_ = ~new_n22943_ & new_n23343_;
  assign new_n23345_ = ~new_n22944_ & ~new_n22947_;
  assign new_n23346_ = ~new_n23344_ & ~new_n23345_;
  assign new_n23347_ = \quotient[7]  & ~new_n23346_;
  assign new_n23348_ = ~new_n22554_ & ~new_n23096_;
  assign new_n23349_ = ~new_n23095_ & new_n23348_;
  assign new_n23350_ = ~new_n23347_ & ~new_n23349_;
  assign new_n23351_ = ~\b[30]  & ~new_n23350_;
  assign new_n23352_ = ~new_n22573_ & new_n22942_;
  assign new_n23353_ = ~new_n22938_ & new_n23352_;
  assign new_n23354_ = ~new_n22939_ & ~new_n22942_;
  assign new_n23355_ = ~new_n23353_ & ~new_n23354_;
  assign new_n23356_ = \quotient[7]  & ~new_n23355_;
  assign new_n23357_ = ~new_n22563_ & ~new_n23096_;
  assign new_n23358_ = ~new_n23095_ & new_n23357_;
  assign new_n23359_ = ~new_n23356_ & ~new_n23358_;
  assign new_n23360_ = ~\b[29]  & ~new_n23359_;
  assign new_n23361_ = ~new_n22582_ & new_n22937_;
  assign new_n23362_ = ~new_n22933_ & new_n23361_;
  assign new_n23363_ = ~new_n22934_ & ~new_n22937_;
  assign new_n23364_ = ~new_n23362_ & ~new_n23363_;
  assign new_n23365_ = \quotient[7]  & ~new_n23364_;
  assign new_n23366_ = ~new_n22572_ & ~new_n23096_;
  assign new_n23367_ = ~new_n23095_ & new_n23366_;
  assign new_n23368_ = ~new_n23365_ & ~new_n23367_;
  assign new_n23369_ = ~\b[28]  & ~new_n23368_;
  assign new_n23370_ = ~new_n22591_ & new_n22932_;
  assign new_n23371_ = ~new_n22928_ & new_n23370_;
  assign new_n23372_ = ~new_n22929_ & ~new_n22932_;
  assign new_n23373_ = ~new_n23371_ & ~new_n23372_;
  assign new_n23374_ = \quotient[7]  & ~new_n23373_;
  assign new_n23375_ = ~new_n22581_ & ~new_n23096_;
  assign new_n23376_ = ~new_n23095_ & new_n23375_;
  assign new_n23377_ = ~new_n23374_ & ~new_n23376_;
  assign new_n23378_ = ~\b[27]  & ~new_n23377_;
  assign new_n23379_ = ~new_n22600_ & new_n22927_;
  assign new_n23380_ = ~new_n22923_ & new_n23379_;
  assign new_n23381_ = ~new_n22924_ & ~new_n22927_;
  assign new_n23382_ = ~new_n23380_ & ~new_n23381_;
  assign new_n23383_ = \quotient[7]  & ~new_n23382_;
  assign new_n23384_ = ~new_n22590_ & ~new_n23096_;
  assign new_n23385_ = ~new_n23095_ & new_n23384_;
  assign new_n23386_ = ~new_n23383_ & ~new_n23385_;
  assign new_n23387_ = ~\b[26]  & ~new_n23386_;
  assign new_n23388_ = ~new_n22609_ & new_n22922_;
  assign new_n23389_ = ~new_n22918_ & new_n23388_;
  assign new_n23390_ = ~new_n22919_ & ~new_n22922_;
  assign new_n23391_ = ~new_n23389_ & ~new_n23390_;
  assign new_n23392_ = \quotient[7]  & ~new_n23391_;
  assign new_n23393_ = ~new_n22599_ & ~new_n23096_;
  assign new_n23394_ = ~new_n23095_ & new_n23393_;
  assign new_n23395_ = ~new_n23392_ & ~new_n23394_;
  assign new_n23396_ = ~\b[25]  & ~new_n23395_;
  assign new_n23397_ = ~new_n22618_ & new_n22917_;
  assign new_n23398_ = ~new_n22913_ & new_n23397_;
  assign new_n23399_ = ~new_n22914_ & ~new_n22917_;
  assign new_n23400_ = ~new_n23398_ & ~new_n23399_;
  assign new_n23401_ = \quotient[7]  & ~new_n23400_;
  assign new_n23402_ = ~new_n22608_ & ~new_n23096_;
  assign new_n23403_ = ~new_n23095_ & new_n23402_;
  assign new_n23404_ = ~new_n23401_ & ~new_n23403_;
  assign new_n23405_ = ~\b[24]  & ~new_n23404_;
  assign new_n23406_ = ~new_n22627_ & new_n22912_;
  assign new_n23407_ = ~new_n22908_ & new_n23406_;
  assign new_n23408_ = ~new_n22909_ & ~new_n22912_;
  assign new_n23409_ = ~new_n23407_ & ~new_n23408_;
  assign new_n23410_ = \quotient[7]  & ~new_n23409_;
  assign new_n23411_ = ~new_n22617_ & ~new_n23096_;
  assign new_n23412_ = ~new_n23095_ & new_n23411_;
  assign new_n23413_ = ~new_n23410_ & ~new_n23412_;
  assign new_n23414_ = ~\b[23]  & ~new_n23413_;
  assign new_n23415_ = ~new_n22636_ & new_n22907_;
  assign new_n23416_ = ~new_n22903_ & new_n23415_;
  assign new_n23417_ = ~new_n22904_ & ~new_n22907_;
  assign new_n23418_ = ~new_n23416_ & ~new_n23417_;
  assign new_n23419_ = \quotient[7]  & ~new_n23418_;
  assign new_n23420_ = ~new_n22626_ & ~new_n23096_;
  assign new_n23421_ = ~new_n23095_ & new_n23420_;
  assign new_n23422_ = ~new_n23419_ & ~new_n23421_;
  assign new_n23423_ = ~\b[22]  & ~new_n23422_;
  assign new_n23424_ = ~new_n22645_ & new_n22902_;
  assign new_n23425_ = ~new_n22898_ & new_n23424_;
  assign new_n23426_ = ~new_n22899_ & ~new_n22902_;
  assign new_n23427_ = ~new_n23425_ & ~new_n23426_;
  assign new_n23428_ = \quotient[7]  & ~new_n23427_;
  assign new_n23429_ = ~new_n22635_ & ~new_n23096_;
  assign new_n23430_ = ~new_n23095_ & new_n23429_;
  assign new_n23431_ = ~new_n23428_ & ~new_n23430_;
  assign new_n23432_ = ~\b[21]  & ~new_n23431_;
  assign new_n23433_ = ~new_n22654_ & new_n22897_;
  assign new_n23434_ = ~new_n22893_ & new_n23433_;
  assign new_n23435_ = ~new_n22894_ & ~new_n22897_;
  assign new_n23436_ = ~new_n23434_ & ~new_n23435_;
  assign new_n23437_ = \quotient[7]  & ~new_n23436_;
  assign new_n23438_ = ~new_n22644_ & ~new_n23096_;
  assign new_n23439_ = ~new_n23095_ & new_n23438_;
  assign new_n23440_ = ~new_n23437_ & ~new_n23439_;
  assign new_n23441_ = ~\b[20]  & ~new_n23440_;
  assign new_n23442_ = ~new_n22663_ & new_n22892_;
  assign new_n23443_ = ~new_n22888_ & new_n23442_;
  assign new_n23444_ = ~new_n22889_ & ~new_n22892_;
  assign new_n23445_ = ~new_n23443_ & ~new_n23444_;
  assign new_n23446_ = \quotient[7]  & ~new_n23445_;
  assign new_n23447_ = ~new_n22653_ & ~new_n23096_;
  assign new_n23448_ = ~new_n23095_ & new_n23447_;
  assign new_n23449_ = ~new_n23446_ & ~new_n23448_;
  assign new_n23450_ = ~\b[19]  & ~new_n23449_;
  assign new_n23451_ = ~new_n22672_ & new_n22887_;
  assign new_n23452_ = ~new_n22883_ & new_n23451_;
  assign new_n23453_ = ~new_n22884_ & ~new_n22887_;
  assign new_n23454_ = ~new_n23452_ & ~new_n23453_;
  assign new_n23455_ = \quotient[7]  & ~new_n23454_;
  assign new_n23456_ = ~new_n22662_ & ~new_n23096_;
  assign new_n23457_ = ~new_n23095_ & new_n23456_;
  assign new_n23458_ = ~new_n23455_ & ~new_n23457_;
  assign new_n23459_ = ~\b[18]  & ~new_n23458_;
  assign new_n23460_ = ~new_n22681_ & new_n22882_;
  assign new_n23461_ = ~new_n22878_ & new_n23460_;
  assign new_n23462_ = ~new_n22879_ & ~new_n22882_;
  assign new_n23463_ = ~new_n23461_ & ~new_n23462_;
  assign new_n23464_ = \quotient[7]  & ~new_n23463_;
  assign new_n23465_ = ~new_n22671_ & ~new_n23096_;
  assign new_n23466_ = ~new_n23095_ & new_n23465_;
  assign new_n23467_ = ~new_n23464_ & ~new_n23466_;
  assign new_n23468_ = ~\b[17]  & ~new_n23467_;
  assign new_n23469_ = ~new_n22690_ & new_n22877_;
  assign new_n23470_ = ~new_n22873_ & new_n23469_;
  assign new_n23471_ = ~new_n22874_ & ~new_n22877_;
  assign new_n23472_ = ~new_n23470_ & ~new_n23471_;
  assign new_n23473_ = \quotient[7]  & ~new_n23472_;
  assign new_n23474_ = ~new_n22680_ & ~new_n23096_;
  assign new_n23475_ = ~new_n23095_ & new_n23474_;
  assign new_n23476_ = ~new_n23473_ & ~new_n23475_;
  assign new_n23477_ = ~\b[16]  & ~new_n23476_;
  assign new_n23478_ = ~new_n22699_ & new_n22872_;
  assign new_n23479_ = ~new_n22868_ & new_n23478_;
  assign new_n23480_ = ~new_n22869_ & ~new_n22872_;
  assign new_n23481_ = ~new_n23479_ & ~new_n23480_;
  assign new_n23482_ = \quotient[7]  & ~new_n23481_;
  assign new_n23483_ = ~new_n22689_ & ~new_n23096_;
  assign new_n23484_ = ~new_n23095_ & new_n23483_;
  assign new_n23485_ = ~new_n23482_ & ~new_n23484_;
  assign new_n23486_ = ~\b[15]  & ~new_n23485_;
  assign new_n23487_ = ~new_n22708_ & new_n22867_;
  assign new_n23488_ = ~new_n22863_ & new_n23487_;
  assign new_n23489_ = ~new_n22864_ & ~new_n22867_;
  assign new_n23490_ = ~new_n23488_ & ~new_n23489_;
  assign new_n23491_ = \quotient[7]  & ~new_n23490_;
  assign new_n23492_ = ~new_n22698_ & ~new_n23096_;
  assign new_n23493_ = ~new_n23095_ & new_n23492_;
  assign new_n23494_ = ~new_n23491_ & ~new_n23493_;
  assign new_n23495_ = ~\b[14]  & ~new_n23494_;
  assign new_n23496_ = ~new_n22717_ & new_n22862_;
  assign new_n23497_ = ~new_n22858_ & new_n23496_;
  assign new_n23498_ = ~new_n22859_ & ~new_n22862_;
  assign new_n23499_ = ~new_n23497_ & ~new_n23498_;
  assign new_n23500_ = \quotient[7]  & ~new_n23499_;
  assign new_n23501_ = ~new_n22707_ & ~new_n23096_;
  assign new_n23502_ = ~new_n23095_ & new_n23501_;
  assign new_n23503_ = ~new_n23500_ & ~new_n23502_;
  assign new_n23504_ = ~\b[13]  & ~new_n23503_;
  assign new_n23505_ = ~new_n22726_ & new_n22857_;
  assign new_n23506_ = ~new_n22853_ & new_n23505_;
  assign new_n23507_ = ~new_n22854_ & ~new_n22857_;
  assign new_n23508_ = ~new_n23506_ & ~new_n23507_;
  assign new_n23509_ = \quotient[7]  & ~new_n23508_;
  assign new_n23510_ = ~new_n22716_ & ~new_n23096_;
  assign new_n23511_ = ~new_n23095_ & new_n23510_;
  assign new_n23512_ = ~new_n23509_ & ~new_n23511_;
  assign new_n23513_ = ~\b[12]  & ~new_n23512_;
  assign new_n23514_ = ~new_n22735_ & new_n22852_;
  assign new_n23515_ = ~new_n22848_ & new_n23514_;
  assign new_n23516_ = ~new_n22849_ & ~new_n22852_;
  assign new_n23517_ = ~new_n23515_ & ~new_n23516_;
  assign new_n23518_ = \quotient[7]  & ~new_n23517_;
  assign new_n23519_ = ~new_n22725_ & ~new_n23096_;
  assign new_n23520_ = ~new_n23095_ & new_n23519_;
  assign new_n23521_ = ~new_n23518_ & ~new_n23520_;
  assign new_n23522_ = ~\b[11]  & ~new_n23521_;
  assign new_n23523_ = ~new_n22744_ & new_n22847_;
  assign new_n23524_ = ~new_n22843_ & new_n23523_;
  assign new_n23525_ = ~new_n22844_ & ~new_n22847_;
  assign new_n23526_ = ~new_n23524_ & ~new_n23525_;
  assign new_n23527_ = \quotient[7]  & ~new_n23526_;
  assign new_n23528_ = ~new_n22734_ & ~new_n23096_;
  assign new_n23529_ = ~new_n23095_ & new_n23528_;
  assign new_n23530_ = ~new_n23527_ & ~new_n23529_;
  assign new_n23531_ = ~\b[10]  & ~new_n23530_;
  assign new_n23532_ = ~new_n22753_ & new_n22842_;
  assign new_n23533_ = ~new_n22838_ & new_n23532_;
  assign new_n23534_ = ~new_n22839_ & ~new_n22842_;
  assign new_n23535_ = ~new_n23533_ & ~new_n23534_;
  assign new_n23536_ = \quotient[7]  & ~new_n23535_;
  assign new_n23537_ = ~new_n22743_ & ~new_n23096_;
  assign new_n23538_ = ~new_n23095_ & new_n23537_;
  assign new_n23539_ = ~new_n23536_ & ~new_n23538_;
  assign new_n23540_ = ~\b[9]  & ~new_n23539_;
  assign new_n23541_ = ~new_n22762_ & new_n22837_;
  assign new_n23542_ = ~new_n22833_ & new_n23541_;
  assign new_n23543_ = ~new_n22834_ & ~new_n22837_;
  assign new_n23544_ = ~new_n23542_ & ~new_n23543_;
  assign new_n23545_ = \quotient[7]  & ~new_n23544_;
  assign new_n23546_ = ~new_n22752_ & ~new_n23096_;
  assign new_n23547_ = ~new_n23095_ & new_n23546_;
  assign new_n23548_ = ~new_n23545_ & ~new_n23547_;
  assign new_n23549_ = ~\b[8]  & ~new_n23548_;
  assign new_n23550_ = ~new_n22771_ & new_n22832_;
  assign new_n23551_ = ~new_n22828_ & new_n23550_;
  assign new_n23552_ = ~new_n22829_ & ~new_n22832_;
  assign new_n23553_ = ~new_n23551_ & ~new_n23552_;
  assign new_n23554_ = \quotient[7]  & ~new_n23553_;
  assign new_n23555_ = ~new_n22761_ & ~new_n23096_;
  assign new_n23556_ = ~new_n23095_ & new_n23555_;
  assign new_n23557_ = ~new_n23554_ & ~new_n23556_;
  assign new_n23558_ = ~\b[7]  & ~new_n23557_;
  assign new_n23559_ = ~new_n22780_ & new_n22827_;
  assign new_n23560_ = ~new_n22823_ & new_n23559_;
  assign new_n23561_ = ~new_n22824_ & ~new_n22827_;
  assign new_n23562_ = ~new_n23560_ & ~new_n23561_;
  assign new_n23563_ = \quotient[7]  & ~new_n23562_;
  assign new_n23564_ = ~new_n22770_ & ~new_n23096_;
  assign new_n23565_ = ~new_n23095_ & new_n23564_;
  assign new_n23566_ = ~new_n23563_ & ~new_n23565_;
  assign new_n23567_ = ~\b[6]  & ~new_n23566_;
  assign new_n23568_ = ~new_n22789_ & new_n22822_;
  assign new_n23569_ = ~new_n22818_ & new_n23568_;
  assign new_n23570_ = ~new_n22819_ & ~new_n22822_;
  assign new_n23571_ = ~new_n23569_ & ~new_n23570_;
  assign new_n23572_ = \quotient[7]  & ~new_n23571_;
  assign new_n23573_ = ~new_n22779_ & ~new_n23096_;
  assign new_n23574_ = ~new_n23095_ & new_n23573_;
  assign new_n23575_ = ~new_n23572_ & ~new_n23574_;
  assign new_n23576_ = ~\b[5]  & ~new_n23575_;
  assign new_n23577_ = ~new_n22797_ & new_n22817_;
  assign new_n23578_ = ~new_n22813_ & new_n23577_;
  assign new_n23579_ = ~new_n22814_ & ~new_n22817_;
  assign new_n23580_ = ~new_n23578_ & ~new_n23579_;
  assign new_n23581_ = \quotient[7]  & ~new_n23580_;
  assign new_n23582_ = ~new_n22788_ & ~new_n23096_;
  assign new_n23583_ = ~new_n23095_ & new_n23582_;
  assign new_n23584_ = ~new_n23581_ & ~new_n23583_;
  assign new_n23585_ = ~\b[4]  & ~new_n23584_;
  assign new_n23586_ = ~new_n22808_ & new_n22812_;
  assign new_n23587_ = ~new_n22807_ & new_n23586_;
  assign new_n23588_ = ~new_n22809_ & ~new_n22812_;
  assign new_n23589_ = ~new_n23587_ & ~new_n23588_;
  assign new_n23590_ = \quotient[7]  & ~new_n23589_;
  assign new_n23591_ = ~new_n22796_ & ~new_n23096_;
  assign new_n23592_ = ~new_n23095_ & new_n23591_;
  assign new_n23593_ = ~new_n23590_ & ~new_n23592_;
  assign new_n23594_ = ~\b[3]  & ~new_n23593_;
  assign new_n23595_ = ~new_n22804_ & new_n22806_;
  assign new_n23596_ = ~new_n22802_ & new_n23595_;
  assign new_n23597_ = ~new_n22807_ & ~new_n23596_;
  assign new_n23598_ = \quotient[7]  & new_n23597_;
  assign new_n23599_ = ~new_n22801_ & ~new_n23096_;
  assign new_n23600_ = ~new_n23095_ & new_n23599_;
  assign new_n23601_ = ~new_n23598_ & ~new_n23600_;
  assign new_n23602_ = ~\b[2]  & ~new_n23601_;
  assign new_n23603_ = \b[0]  & \quotient[7] ;
  assign new_n23604_ = \a[7]  & ~new_n23603_;
  assign new_n23605_ = new_n22806_ & \quotient[7] ;
  assign new_n23606_ = ~new_n23604_ & ~new_n23605_;
  assign new_n23607_ = \b[1]  & ~new_n23606_;
  assign new_n23608_ = ~\b[1]  & ~new_n23605_;
  assign new_n23609_ = ~new_n23604_ & new_n23608_;
  assign new_n23610_ = ~new_n23607_ & ~new_n23609_;
  assign new_n23611_ = ~\a[6]  & \b[0] ;
  assign new_n23612_ = ~new_n23610_ & ~new_n23611_;
  assign new_n23613_ = ~\b[1]  & ~new_n23606_;
  assign new_n23614_ = ~new_n23612_ & ~new_n23613_;
  assign new_n23615_ = \b[2]  & ~new_n23600_;
  assign new_n23616_ = ~new_n23598_ & new_n23615_;
  assign new_n23617_ = ~new_n23602_ & ~new_n23616_;
  assign new_n23618_ = ~new_n23614_ & new_n23617_;
  assign new_n23619_ = ~new_n23602_ & ~new_n23618_;
  assign new_n23620_ = \b[3]  & ~new_n23592_;
  assign new_n23621_ = ~new_n23590_ & new_n23620_;
  assign new_n23622_ = ~new_n23594_ & ~new_n23621_;
  assign new_n23623_ = ~new_n23619_ & new_n23622_;
  assign new_n23624_ = ~new_n23594_ & ~new_n23623_;
  assign new_n23625_ = \b[4]  & ~new_n23583_;
  assign new_n23626_ = ~new_n23581_ & new_n23625_;
  assign new_n23627_ = ~new_n23585_ & ~new_n23626_;
  assign new_n23628_ = ~new_n23624_ & new_n23627_;
  assign new_n23629_ = ~new_n23585_ & ~new_n23628_;
  assign new_n23630_ = \b[5]  & ~new_n23574_;
  assign new_n23631_ = ~new_n23572_ & new_n23630_;
  assign new_n23632_ = ~new_n23576_ & ~new_n23631_;
  assign new_n23633_ = ~new_n23629_ & new_n23632_;
  assign new_n23634_ = ~new_n23576_ & ~new_n23633_;
  assign new_n23635_ = \b[6]  & ~new_n23565_;
  assign new_n23636_ = ~new_n23563_ & new_n23635_;
  assign new_n23637_ = ~new_n23567_ & ~new_n23636_;
  assign new_n23638_ = ~new_n23634_ & new_n23637_;
  assign new_n23639_ = ~new_n23567_ & ~new_n23638_;
  assign new_n23640_ = \b[7]  & ~new_n23556_;
  assign new_n23641_ = ~new_n23554_ & new_n23640_;
  assign new_n23642_ = ~new_n23558_ & ~new_n23641_;
  assign new_n23643_ = ~new_n23639_ & new_n23642_;
  assign new_n23644_ = ~new_n23558_ & ~new_n23643_;
  assign new_n23645_ = \b[8]  & ~new_n23547_;
  assign new_n23646_ = ~new_n23545_ & new_n23645_;
  assign new_n23647_ = ~new_n23549_ & ~new_n23646_;
  assign new_n23648_ = ~new_n23644_ & new_n23647_;
  assign new_n23649_ = ~new_n23549_ & ~new_n23648_;
  assign new_n23650_ = \b[9]  & ~new_n23538_;
  assign new_n23651_ = ~new_n23536_ & new_n23650_;
  assign new_n23652_ = ~new_n23540_ & ~new_n23651_;
  assign new_n23653_ = ~new_n23649_ & new_n23652_;
  assign new_n23654_ = ~new_n23540_ & ~new_n23653_;
  assign new_n23655_ = \b[10]  & ~new_n23529_;
  assign new_n23656_ = ~new_n23527_ & new_n23655_;
  assign new_n23657_ = ~new_n23531_ & ~new_n23656_;
  assign new_n23658_ = ~new_n23654_ & new_n23657_;
  assign new_n23659_ = ~new_n23531_ & ~new_n23658_;
  assign new_n23660_ = \b[11]  & ~new_n23520_;
  assign new_n23661_ = ~new_n23518_ & new_n23660_;
  assign new_n23662_ = ~new_n23522_ & ~new_n23661_;
  assign new_n23663_ = ~new_n23659_ & new_n23662_;
  assign new_n23664_ = ~new_n23522_ & ~new_n23663_;
  assign new_n23665_ = \b[12]  & ~new_n23511_;
  assign new_n23666_ = ~new_n23509_ & new_n23665_;
  assign new_n23667_ = ~new_n23513_ & ~new_n23666_;
  assign new_n23668_ = ~new_n23664_ & new_n23667_;
  assign new_n23669_ = ~new_n23513_ & ~new_n23668_;
  assign new_n23670_ = \b[13]  & ~new_n23502_;
  assign new_n23671_ = ~new_n23500_ & new_n23670_;
  assign new_n23672_ = ~new_n23504_ & ~new_n23671_;
  assign new_n23673_ = ~new_n23669_ & new_n23672_;
  assign new_n23674_ = ~new_n23504_ & ~new_n23673_;
  assign new_n23675_ = \b[14]  & ~new_n23493_;
  assign new_n23676_ = ~new_n23491_ & new_n23675_;
  assign new_n23677_ = ~new_n23495_ & ~new_n23676_;
  assign new_n23678_ = ~new_n23674_ & new_n23677_;
  assign new_n23679_ = ~new_n23495_ & ~new_n23678_;
  assign new_n23680_ = \b[15]  & ~new_n23484_;
  assign new_n23681_ = ~new_n23482_ & new_n23680_;
  assign new_n23682_ = ~new_n23486_ & ~new_n23681_;
  assign new_n23683_ = ~new_n23679_ & new_n23682_;
  assign new_n23684_ = ~new_n23486_ & ~new_n23683_;
  assign new_n23685_ = \b[16]  & ~new_n23475_;
  assign new_n23686_ = ~new_n23473_ & new_n23685_;
  assign new_n23687_ = ~new_n23477_ & ~new_n23686_;
  assign new_n23688_ = ~new_n23684_ & new_n23687_;
  assign new_n23689_ = ~new_n23477_ & ~new_n23688_;
  assign new_n23690_ = \b[17]  & ~new_n23466_;
  assign new_n23691_ = ~new_n23464_ & new_n23690_;
  assign new_n23692_ = ~new_n23468_ & ~new_n23691_;
  assign new_n23693_ = ~new_n23689_ & new_n23692_;
  assign new_n23694_ = ~new_n23468_ & ~new_n23693_;
  assign new_n23695_ = \b[18]  & ~new_n23457_;
  assign new_n23696_ = ~new_n23455_ & new_n23695_;
  assign new_n23697_ = ~new_n23459_ & ~new_n23696_;
  assign new_n23698_ = ~new_n23694_ & new_n23697_;
  assign new_n23699_ = ~new_n23459_ & ~new_n23698_;
  assign new_n23700_ = \b[19]  & ~new_n23448_;
  assign new_n23701_ = ~new_n23446_ & new_n23700_;
  assign new_n23702_ = ~new_n23450_ & ~new_n23701_;
  assign new_n23703_ = ~new_n23699_ & new_n23702_;
  assign new_n23704_ = ~new_n23450_ & ~new_n23703_;
  assign new_n23705_ = \b[20]  & ~new_n23439_;
  assign new_n23706_ = ~new_n23437_ & new_n23705_;
  assign new_n23707_ = ~new_n23441_ & ~new_n23706_;
  assign new_n23708_ = ~new_n23704_ & new_n23707_;
  assign new_n23709_ = ~new_n23441_ & ~new_n23708_;
  assign new_n23710_ = \b[21]  & ~new_n23430_;
  assign new_n23711_ = ~new_n23428_ & new_n23710_;
  assign new_n23712_ = ~new_n23432_ & ~new_n23711_;
  assign new_n23713_ = ~new_n23709_ & new_n23712_;
  assign new_n23714_ = ~new_n23432_ & ~new_n23713_;
  assign new_n23715_ = \b[22]  & ~new_n23421_;
  assign new_n23716_ = ~new_n23419_ & new_n23715_;
  assign new_n23717_ = ~new_n23423_ & ~new_n23716_;
  assign new_n23718_ = ~new_n23714_ & new_n23717_;
  assign new_n23719_ = ~new_n23423_ & ~new_n23718_;
  assign new_n23720_ = \b[23]  & ~new_n23412_;
  assign new_n23721_ = ~new_n23410_ & new_n23720_;
  assign new_n23722_ = ~new_n23414_ & ~new_n23721_;
  assign new_n23723_ = ~new_n23719_ & new_n23722_;
  assign new_n23724_ = ~new_n23414_ & ~new_n23723_;
  assign new_n23725_ = \b[24]  & ~new_n23403_;
  assign new_n23726_ = ~new_n23401_ & new_n23725_;
  assign new_n23727_ = ~new_n23405_ & ~new_n23726_;
  assign new_n23728_ = ~new_n23724_ & new_n23727_;
  assign new_n23729_ = ~new_n23405_ & ~new_n23728_;
  assign new_n23730_ = \b[25]  & ~new_n23394_;
  assign new_n23731_ = ~new_n23392_ & new_n23730_;
  assign new_n23732_ = ~new_n23396_ & ~new_n23731_;
  assign new_n23733_ = ~new_n23729_ & new_n23732_;
  assign new_n23734_ = ~new_n23396_ & ~new_n23733_;
  assign new_n23735_ = \b[26]  & ~new_n23385_;
  assign new_n23736_ = ~new_n23383_ & new_n23735_;
  assign new_n23737_ = ~new_n23387_ & ~new_n23736_;
  assign new_n23738_ = ~new_n23734_ & new_n23737_;
  assign new_n23739_ = ~new_n23387_ & ~new_n23738_;
  assign new_n23740_ = \b[27]  & ~new_n23376_;
  assign new_n23741_ = ~new_n23374_ & new_n23740_;
  assign new_n23742_ = ~new_n23378_ & ~new_n23741_;
  assign new_n23743_ = ~new_n23739_ & new_n23742_;
  assign new_n23744_ = ~new_n23378_ & ~new_n23743_;
  assign new_n23745_ = \b[28]  & ~new_n23367_;
  assign new_n23746_ = ~new_n23365_ & new_n23745_;
  assign new_n23747_ = ~new_n23369_ & ~new_n23746_;
  assign new_n23748_ = ~new_n23744_ & new_n23747_;
  assign new_n23749_ = ~new_n23369_ & ~new_n23748_;
  assign new_n23750_ = \b[29]  & ~new_n23358_;
  assign new_n23751_ = ~new_n23356_ & new_n23750_;
  assign new_n23752_ = ~new_n23360_ & ~new_n23751_;
  assign new_n23753_ = ~new_n23749_ & new_n23752_;
  assign new_n23754_ = ~new_n23360_ & ~new_n23753_;
  assign new_n23755_ = \b[30]  & ~new_n23349_;
  assign new_n23756_ = ~new_n23347_ & new_n23755_;
  assign new_n23757_ = ~new_n23351_ & ~new_n23756_;
  assign new_n23758_ = ~new_n23754_ & new_n23757_;
  assign new_n23759_ = ~new_n23351_ & ~new_n23758_;
  assign new_n23760_ = \b[31]  & ~new_n23340_;
  assign new_n23761_ = ~new_n23338_ & new_n23760_;
  assign new_n23762_ = ~new_n23342_ & ~new_n23761_;
  assign new_n23763_ = ~new_n23759_ & new_n23762_;
  assign new_n23764_ = ~new_n23342_ & ~new_n23763_;
  assign new_n23765_ = \b[32]  & ~new_n23331_;
  assign new_n23766_ = ~new_n23329_ & new_n23765_;
  assign new_n23767_ = ~new_n23333_ & ~new_n23766_;
  assign new_n23768_ = ~new_n23764_ & new_n23767_;
  assign new_n23769_ = ~new_n23333_ & ~new_n23768_;
  assign new_n23770_ = \b[33]  & ~new_n23322_;
  assign new_n23771_ = ~new_n23320_ & new_n23770_;
  assign new_n23772_ = ~new_n23324_ & ~new_n23771_;
  assign new_n23773_ = ~new_n23769_ & new_n23772_;
  assign new_n23774_ = ~new_n23324_ & ~new_n23773_;
  assign new_n23775_ = \b[34]  & ~new_n23313_;
  assign new_n23776_ = ~new_n23311_ & new_n23775_;
  assign new_n23777_ = ~new_n23315_ & ~new_n23776_;
  assign new_n23778_ = ~new_n23774_ & new_n23777_;
  assign new_n23779_ = ~new_n23315_ & ~new_n23778_;
  assign new_n23780_ = \b[35]  & ~new_n23304_;
  assign new_n23781_ = ~new_n23302_ & new_n23780_;
  assign new_n23782_ = ~new_n23306_ & ~new_n23781_;
  assign new_n23783_ = ~new_n23779_ & new_n23782_;
  assign new_n23784_ = ~new_n23306_ & ~new_n23783_;
  assign new_n23785_ = \b[36]  & ~new_n23295_;
  assign new_n23786_ = ~new_n23293_ & new_n23785_;
  assign new_n23787_ = ~new_n23297_ & ~new_n23786_;
  assign new_n23788_ = ~new_n23784_ & new_n23787_;
  assign new_n23789_ = ~new_n23297_ & ~new_n23788_;
  assign new_n23790_ = \b[37]  & ~new_n23286_;
  assign new_n23791_ = ~new_n23284_ & new_n23790_;
  assign new_n23792_ = ~new_n23288_ & ~new_n23791_;
  assign new_n23793_ = ~new_n23789_ & new_n23792_;
  assign new_n23794_ = ~new_n23288_ & ~new_n23793_;
  assign new_n23795_ = \b[38]  & ~new_n23277_;
  assign new_n23796_ = ~new_n23275_ & new_n23795_;
  assign new_n23797_ = ~new_n23279_ & ~new_n23796_;
  assign new_n23798_ = ~new_n23794_ & new_n23797_;
  assign new_n23799_ = ~new_n23279_ & ~new_n23798_;
  assign new_n23800_ = \b[39]  & ~new_n23268_;
  assign new_n23801_ = ~new_n23266_ & new_n23800_;
  assign new_n23802_ = ~new_n23270_ & ~new_n23801_;
  assign new_n23803_ = ~new_n23799_ & new_n23802_;
  assign new_n23804_ = ~new_n23270_ & ~new_n23803_;
  assign new_n23805_ = \b[40]  & ~new_n23259_;
  assign new_n23806_ = ~new_n23257_ & new_n23805_;
  assign new_n23807_ = ~new_n23261_ & ~new_n23806_;
  assign new_n23808_ = ~new_n23804_ & new_n23807_;
  assign new_n23809_ = ~new_n23261_ & ~new_n23808_;
  assign new_n23810_ = \b[41]  & ~new_n23250_;
  assign new_n23811_ = ~new_n23248_ & new_n23810_;
  assign new_n23812_ = ~new_n23252_ & ~new_n23811_;
  assign new_n23813_ = ~new_n23809_ & new_n23812_;
  assign new_n23814_ = ~new_n23252_ & ~new_n23813_;
  assign new_n23815_ = \b[42]  & ~new_n23241_;
  assign new_n23816_ = ~new_n23239_ & new_n23815_;
  assign new_n23817_ = ~new_n23243_ & ~new_n23816_;
  assign new_n23818_ = ~new_n23814_ & new_n23817_;
  assign new_n23819_ = ~new_n23243_ & ~new_n23818_;
  assign new_n23820_ = \b[43]  & ~new_n23232_;
  assign new_n23821_ = ~new_n23230_ & new_n23820_;
  assign new_n23822_ = ~new_n23234_ & ~new_n23821_;
  assign new_n23823_ = ~new_n23819_ & new_n23822_;
  assign new_n23824_ = ~new_n23234_ & ~new_n23823_;
  assign new_n23825_ = \b[44]  & ~new_n23223_;
  assign new_n23826_ = ~new_n23221_ & new_n23825_;
  assign new_n23827_ = ~new_n23225_ & ~new_n23826_;
  assign new_n23828_ = ~new_n23824_ & new_n23827_;
  assign new_n23829_ = ~new_n23225_ & ~new_n23828_;
  assign new_n23830_ = \b[45]  & ~new_n23214_;
  assign new_n23831_ = ~new_n23212_ & new_n23830_;
  assign new_n23832_ = ~new_n23216_ & ~new_n23831_;
  assign new_n23833_ = ~new_n23829_ & new_n23832_;
  assign new_n23834_ = ~new_n23216_ & ~new_n23833_;
  assign new_n23835_ = \b[46]  & ~new_n23205_;
  assign new_n23836_ = ~new_n23203_ & new_n23835_;
  assign new_n23837_ = ~new_n23207_ & ~new_n23836_;
  assign new_n23838_ = ~new_n23834_ & new_n23837_;
  assign new_n23839_ = ~new_n23207_ & ~new_n23838_;
  assign new_n23840_ = \b[47]  & ~new_n23196_;
  assign new_n23841_ = ~new_n23194_ & new_n23840_;
  assign new_n23842_ = ~new_n23198_ & ~new_n23841_;
  assign new_n23843_ = ~new_n23839_ & new_n23842_;
  assign new_n23844_ = ~new_n23198_ & ~new_n23843_;
  assign new_n23845_ = \b[48]  & ~new_n23187_;
  assign new_n23846_ = ~new_n23185_ & new_n23845_;
  assign new_n23847_ = ~new_n23189_ & ~new_n23846_;
  assign new_n23848_ = ~new_n23844_ & new_n23847_;
  assign new_n23849_ = ~new_n23189_ & ~new_n23848_;
  assign new_n23850_ = \b[49]  & ~new_n23178_;
  assign new_n23851_ = ~new_n23176_ & new_n23850_;
  assign new_n23852_ = ~new_n23180_ & ~new_n23851_;
  assign new_n23853_ = ~new_n23849_ & new_n23852_;
  assign new_n23854_ = ~new_n23180_ & ~new_n23853_;
  assign new_n23855_ = \b[50]  & ~new_n23169_;
  assign new_n23856_ = ~new_n23167_ & new_n23855_;
  assign new_n23857_ = ~new_n23171_ & ~new_n23856_;
  assign new_n23858_ = ~new_n23854_ & new_n23857_;
  assign new_n23859_ = ~new_n23171_ & ~new_n23858_;
  assign new_n23860_ = \b[51]  & ~new_n23160_;
  assign new_n23861_ = ~new_n23158_ & new_n23860_;
  assign new_n23862_ = ~new_n23162_ & ~new_n23861_;
  assign new_n23863_ = ~new_n23859_ & new_n23862_;
  assign new_n23864_ = ~new_n23162_ & ~new_n23863_;
  assign new_n23865_ = \b[52]  & ~new_n23151_;
  assign new_n23866_ = ~new_n23149_ & new_n23865_;
  assign new_n23867_ = ~new_n23153_ & ~new_n23866_;
  assign new_n23868_ = ~new_n23864_ & new_n23867_;
  assign new_n23869_ = ~new_n23153_ & ~new_n23868_;
  assign new_n23870_ = \b[53]  & ~new_n23142_;
  assign new_n23871_ = ~new_n23140_ & new_n23870_;
  assign new_n23872_ = ~new_n23144_ & ~new_n23871_;
  assign new_n23873_ = ~new_n23869_ & new_n23872_;
  assign new_n23874_ = ~new_n23144_ & ~new_n23873_;
  assign new_n23875_ = \b[54]  & ~new_n23133_;
  assign new_n23876_ = ~new_n23131_ & new_n23875_;
  assign new_n23877_ = ~new_n23135_ & ~new_n23876_;
  assign new_n23878_ = ~new_n23874_ & new_n23877_;
  assign new_n23879_ = ~new_n23135_ & ~new_n23878_;
  assign new_n23880_ = \b[55]  & ~new_n23124_;
  assign new_n23881_ = ~new_n23122_ & new_n23880_;
  assign new_n23882_ = ~new_n23126_ & ~new_n23881_;
  assign new_n23883_ = ~new_n23879_ & new_n23882_;
  assign new_n23884_ = ~new_n23126_ & ~new_n23883_;
  assign new_n23885_ = \b[56]  & ~new_n23104_;
  assign new_n23886_ = ~new_n23102_ & new_n23885_;
  assign new_n23887_ = ~new_n23117_ & ~new_n23886_;
  assign new_n23888_ = ~new_n23884_ & new_n23887_;
  assign new_n23889_ = ~new_n23117_ & ~new_n23888_;
  assign new_n23890_ = \b[57]  & ~new_n23114_;
  assign new_n23891_ = ~new_n23112_ & new_n23890_;
  assign new_n23892_ = ~new_n23116_ & ~new_n23891_;
  assign new_n23893_ = ~new_n23889_ & new_n23892_;
  assign new_n23894_ = ~new_n23116_ & ~new_n23893_;
  assign new_n23895_ = new_n280_ & new_n282_;
  assign \quotient[6]  = ~new_n23894_ & new_n23895_;
  assign new_n23897_ = ~new_n23105_ & ~\quotient[6] ;
  assign new_n23898_ = ~new_n23126_ & new_n23887_;
  assign new_n23899_ = ~new_n23883_ & new_n23898_;
  assign new_n23900_ = ~new_n23884_ & ~new_n23887_;
  assign new_n23901_ = ~new_n23899_ & ~new_n23900_;
  assign new_n23902_ = new_n23895_ & ~new_n23901_;
  assign new_n23903_ = ~new_n23894_ & new_n23902_;
  assign new_n23904_ = ~new_n23897_ & ~new_n23903_;
  assign new_n23905_ = ~\b[57]  & ~new_n23904_;
  assign new_n23906_ = ~new_n23125_ & ~\quotient[6] ;
  assign new_n23907_ = ~new_n23135_ & new_n23882_;
  assign new_n23908_ = ~new_n23878_ & new_n23907_;
  assign new_n23909_ = ~new_n23879_ & ~new_n23882_;
  assign new_n23910_ = ~new_n23908_ & ~new_n23909_;
  assign new_n23911_ = new_n23895_ & ~new_n23910_;
  assign new_n23912_ = ~new_n23894_ & new_n23911_;
  assign new_n23913_ = ~new_n23906_ & ~new_n23912_;
  assign new_n23914_ = ~\b[56]  & ~new_n23913_;
  assign new_n23915_ = ~new_n23134_ & ~\quotient[6] ;
  assign new_n23916_ = ~new_n23144_ & new_n23877_;
  assign new_n23917_ = ~new_n23873_ & new_n23916_;
  assign new_n23918_ = ~new_n23874_ & ~new_n23877_;
  assign new_n23919_ = ~new_n23917_ & ~new_n23918_;
  assign new_n23920_ = new_n23895_ & ~new_n23919_;
  assign new_n23921_ = ~new_n23894_ & new_n23920_;
  assign new_n23922_ = ~new_n23915_ & ~new_n23921_;
  assign new_n23923_ = ~\b[55]  & ~new_n23922_;
  assign new_n23924_ = ~new_n23143_ & ~\quotient[6] ;
  assign new_n23925_ = ~new_n23153_ & new_n23872_;
  assign new_n23926_ = ~new_n23868_ & new_n23925_;
  assign new_n23927_ = ~new_n23869_ & ~new_n23872_;
  assign new_n23928_ = ~new_n23926_ & ~new_n23927_;
  assign new_n23929_ = new_n23895_ & ~new_n23928_;
  assign new_n23930_ = ~new_n23894_ & new_n23929_;
  assign new_n23931_ = ~new_n23924_ & ~new_n23930_;
  assign new_n23932_ = ~\b[54]  & ~new_n23931_;
  assign new_n23933_ = ~new_n23152_ & ~\quotient[6] ;
  assign new_n23934_ = ~new_n23162_ & new_n23867_;
  assign new_n23935_ = ~new_n23863_ & new_n23934_;
  assign new_n23936_ = ~new_n23864_ & ~new_n23867_;
  assign new_n23937_ = ~new_n23935_ & ~new_n23936_;
  assign new_n23938_ = new_n23895_ & ~new_n23937_;
  assign new_n23939_ = ~new_n23894_ & new_n23938_;
  assign new_n23940_ = ~new_n23933_ & ~new_n23939_;
  assign new_n23941_ = ~\b[53]  & ~new_n23940_;
  assign new_n23942_ = ~new_n23161_ & ~\quotient[6] ;
  assign new_n23943_ = ~new_n23171_ & new_n23862_;
  assign new_n23944_ = ~new_n23858_ & new_n23943_;
  assign new_n23945_ = ~new_n23859_ & ~new_n23862_;
  assign new_n23946_ = ~new_n23944_ & ~new_n23945_;
  assign new_n23947_ = new_n23895_ & ~new_n23946_;
  assign new_n23948_ = ~new_n23894_ & new_n23947_;
  assign new_n23949_ = ~new_n23942_ & ~new_n23948_;
  assign new_n23950_ = ~\b[52]  & ~new_n23949_;
  assign new_n23951_ = ~new_n23170_ & ~\quotient[6] ;
  assign new_n23952_ = ~new_n23180_ & new_n23857_;
  assign new_n23953_ = ~new_n23853_ & new_n23952_;
  assign new_n23954_ = ~new_n23854_ & ~new_n23857_;
  assign new_n23955_ = ~new_n23953_ & ~new_n23954_;
  assign new_n23956_ = new_n23895_ & ~new_n23955_;
  assign new_n23957_ = ~new_n23894_ & new_n23956_;
  assign new_n23958_ = ~new_n23951_ & ~new_n23957_;
  assign new_n23959_ = ~\b[51]  & ~new_n23958_;
  assign new_n23960_ = ~new_n23179_ & ~\quotient[6] ;
  assign new_n23961_ = ~new_n23189_ & new_n23852_;
  assign new_n23962_ = ~new_n23848_ & new_n23961_;
  assign new_n23963_ = ~new_n23849_ & ~new_n23852_;
  assign new_n23964_ = ~new_n23962_ & ~new_n23963_;
  assign new_n23965_ = new_n23895_ & ~new_n23964_;
  assign new_n23966_ = ~new_n23894_ & new_n23965_;
  assign new_n23967_ = ~new_n23960_ & ~new_n23966_;
  assign new_n23968_ = ~\b[50]  & ~new_n23967_;
  assign new_n23969_ = ~new_n23188_ & ~\quotient[6] ;
  assign new_n23970_ = ~new_n23198_ & new_n23847_;
  assign new_n23971_ = ~new_n23843_ & new_n23970_;
  assign new_n23972_ = ~new_n23844_ & ~new_n23847_;
  assign new_n23973_ = ~new_n23971_ & ~new_n23972_;
  assign new_n23974_ = new_n23895_ & ~new_n23973_;
  assign new_n23975_ = ~new_n23894_ & new_n23974_;
  assign new_n23976_ = ~new_n23969_ & ~new_n23975_;
  assign new_n23977_ = ~\b[49]  & ~new_n23976_;
  assign new_n23978_ = ~new_n23197_ & ~\quotient[6] ;
  assign new_n23979_ = ~new_n23207_ & new_n23842_;
  assign new_n23980_ = ~new_n23838_ & new_n23979_;
  assign new_n23981_ = ~new_n23839_ & ~new_n23842_;
  assign new_n23982_ = ~new_n23980_ & ~new_n23981_;
  assign new_n23983_ = new_n23895_ & ~new_n23982_;
  assign new_n23984_ = ~new_n23894_ & new_n23983_;
  assign new_n23985_ = ~new_n23978_ & ~new_n23984_;
  assign new_n23986_ = ~\b[48]  & ~new_n23985_;
  assign new_n23987_ = ~new_n23206_ & ~\quotient[6] ;
  assign new_n23988_ = ~new_n23216_ & new_n23837_;
  assign new_n23989_ = ~new_n23833_ & new_n23988_;
  assign new_n23990_ = ~new_n23834_ & ~new_n23837_;
  assign new_n23991_ = ~new_n23989_ & ~new_n23990_;
  assign new_n23992_ = new_n23895_ & ~new_n23991_;
  assign new_n23993_ = ~new_n23894_ & new_n23992_;
  assign new_n23994_ = ~new_n23987_ & ~new_n23993_;
  assign new_n23995_ = ~\b[47]  & ~new_n23994_;
  assign new_n23996_ = ~new_n23215_ & ~\quotient[6] ;
  assign new_n23997_ = ~new_n23225_ & new_n23832_;
  assign new_n23998_ = ~new_n23828_ & new_n23997_;
  assign new_n23999_ = ~new_n23829_ & ~new_n23832_;
  assign new_n24000_ = ~new_n23998_ & ~new_n23999_;
  assign new_n24001_ = new_n23895_ & ~new_n24000_;
  assign new_n24002_ = ~new_n23894_ & new_n24001_;
  assign new_n24003_ = ~new_n23996_ & ~new_n24002_;
  assign new_n24004_ = ~\b[46]  & ~new_n24003_;
  assign new_n24005_ = ~new_n23224_ & ~\quotient[6] ;
  assign new_n24006_ = ~new_n23234_ & new_n23827_;
  assign new_n24007_ = ~new_n23823_ & new_n24006_;
  assign new_n24008_ = ~new_n23824_ & ~new_n23827_;
  assign new_n24009_ = ~new_n24007_ & ~new_n24008_;
  assign new_n24010_ = new_n23895_ & ~new_n24009_;
  assign new_n24011_ = ~new_n23894_ & new_n24010_;
  assign new_n24012_ = ~new_n24005_ & ~new_n24011_;
  assign new_n24013_ = ~\b[45]  & ~new_n24012_;
  assign new_n24014_ = ~new_n23233_ & ~\quotient[6] ;
  assign new_n24015_ = ~new_n23243_ & new_n23822_;
  assign new_n24016_ = ~new_n23818_ & new_n24015_;
  assign new_n24017_ = ~new_n23819_ & ~new_n23822_;
  assign new_n24018_ = ~new_n24016_ & ~new_n24017_;
  assign new_n24019_ = new_n23895_ & ~new_n24018_;
  assign new_n24020_ = ~new_n23894_ & new_n24019_;
  assign new_n24021_ = ~new_n24014_ & ~new_n24020_;
  assign new_n24022_ = ~\b[44]  & ~new_n24021_;
  assign new_n24023_ = ~new_n23242_ & ~\quotient[6] ;
  assign new_n24024_ = ~new_n23252_ & new_n23817_;
  assign new_n24025_ = ~new_n23813_ & new_n24024_;
  assign new_n24026_ = ~new_n23814_ & ~new_n23817_;
  assign new_n24027_ = ~new_n24025_ & ~new_n24026_;
  assign new_n24028_ = new_n23895_ & ~new_n24027_;
  assign new_n24029_ = ~new_n23894_ & new_n24028_;
  assign new_n24030_ = ~new_n24023_ & ~new_n24029_;
  assign new_n24031_ = ~\b[43]  & ~new_n24030_;
  assign new_n24032_ = ~new_n23251_ & ~\quotient[6] ;
  assign new_n24033_ = ~new_n23261_ & new_n23812_;
  assign new_n24034_ = ~new_n23808_ & new_n24033_;
  assign new_n24035_ = ~new_n23809_ & ~new_n23812_;
  assign new_n24036_ = ~new_n24034_ & ~new_n24035_;
  assign new_n24037_ = new_n23895_ & ~new_n24036_;
  assign new_n24038_ = ~new_n23894_ & new_n24037_;
  assign new_n24039_ = ~new_n24032_ & ~new_n24038_;
  assign new_n24040_ = ~\b[42]  & ~new_n24039_;
  assign new_n24041_ = ~new_n23260_ & ~\quotient[6] ;
  assign new_n24042_ = ~new_n23270_ & new_n23807_;
  assign new_n24043_ = ~new_n23803_ & new_n24042_;
  assign new_n24044_ = ~new_n23804_ & ~new_n23807_;
  assign new_n24045_ = ~new_n24043_ & ~new_n24044_;
  assign new_n24046_ = new_n23895_ & ~new_n24045_;
  assign new_n24047_ = ~new_n23894_ & new_n24046_;
  assign new_n24048_ = ~new_n24041_ & ~new_n24047_;
  assign new_n24049_ = ~\b[41]  & ~new_n24048_;
  assign new_n24050_ = ~new_n23269_ & ~\quotient[6] ;
  assign new_n24051_ = ~new_n23279_ & new_n23802_;
  assign new_n24052_ = ~new_n23798_ & new_n24051_;
  assign new_n24053_ = ~new_n23799_ & ~new_n23802_;
  assign new_n24054_ = ~new_n24052_ & ~new_n24053_;
  assign new_n24055_ = new_n23895_ & ~new_n24054_;
  assign new_n24056_ = ~new_n23894_ & new_n24055_;
  assign new_n24057_ = ~new_n24050_ & ~new_n24056_;
  assign new_n24058_ = ~\b[40]  & ~new_n24057_;
  assign new_n24059_ = ~new_n23278_ & ~\quotient[6] ;
  assign new_n24060_ = ~new_n23288_ & new_n23797_;
  assign new_n24061_ = ~new_n23793_ & new_n24060_;
  assign new_n24062_ = ~new_n23794_ & ~new_n23797_;
  assign new_n24063_ = ~new_n24061_ & ~new_n24062_;
  assign new_n24064_ = new_n23895_ & ~new_n24063_;
  assign new_n24065_ = ~new_n23894_ & new_n24064_;
  assign new_n24066_ = ~new_n24059_ & ~new_n24065_;
  assign new_n24067_ = ~\b[39]  & ~new_n24066_;
  assign new_n24068_ = ~new_n23287_ & ~\quotient[6] ;
  assign new_n24069_ = ~new_n23297_ & new_n23792_;
  assign new_n24070_ = ~new_n23788_ & new_n24069_;
  assign new_n24071_ = ~new_n23789_ & ~new_n23792_;
  assign new_n24072_ = ~new_n24070_ & ~new_n24071_;
  assign new_n24073_ = new_n23895_ & ~new_n24072_;
  assign new_n24074_ = ~new_n23894_ & new_n24073_;
  assign new_n24075_ = ~new_n24068_ & ~new_n24074_;
  assign new_n24076_ = ~\b[38]  & ~new_n24075_;
  assign new_n24077_ = ~new_n23296_ & ~\quotient[6] ;
  assign new_n24078_ = ~new_n23306_ & new_n23787_;
  assign new_n24079_ = ~new_n23783_ & new_n24078_;
  assign new_n24080_ = ~new_n23784_ & ~new_n23787_;
  assign new_n24081_ = ~new_n24079_ & ~new_n24080_;
  assign new_n24082_ = new_n23895_ & ~new_n24081_;
  assign new_n24083_ = ~new_n23894_ & new_n24082_;
  assign new_n24084_ = ~new_n24077_ & ~new_n24083_;
  assign new_n24085_ = ~\b[37]  & ~new_n24084_;
  assign new_n24086_ = ~new_n23305_ & ~\quotient[6] ;
  assign new_n24087_ = ~new_n23315_ & new_n23782_;
  assign new_n24088_ = ~new_n23778_ & new_n24087_;
  assign new_n24089_ = ~new_n23779_ & ~new_n23782_;
  assign new_n24090_ = ~new_n24088_ & ~new_n24089_;
  assign new_n24091_ = new_n23895_ & ~new_n24090_;
  assign new_n24092_ = ~new_n23894_ & new_n24091_;
  assign new_n24093_ = ~new_n24086_ & ~new_n24092_;
  assign new_n24094_ = ~\b[36]  & ~new_n24093_;
  assign new_n24095_ = ~new_n23314_ & ~\quotient[6] ;
  assign new_n24096_ = ~new_n23324_ & new_n23777_;
  assign new_n24097_ = ~new_n23773_ & new_n24096_;
  assign new_n24098_ = ~new_n23774_ & ~new_n23777_;
  assign new_n24099_ = ~new_n24097_ & ~new_n24098_;
  assign new_n24100_ = new_n23895_ & ~new_n24099_;
  assign new_n24101_ = ~new_n23894_ & new_n24100_;
  assign new_n24102_ = ~new_n24095_ & ~new_n24101_;
  assign new_n24103_ = ~\b[35]  & ~new_n24102_;
  assign new_n24104_ = ~new_n23323_ & ~\quotient[6] ;
  assign new_n24105_ = ~new_n23333_ & new_n23772_;
  assign new_n24106_ = ~new_n23768_ & new_n24105_;
  assign new_n24107_ = ~new_n23769_ & ~new_n23772_;
  assign new_n24108_ = ~new_n24106_ & ~new_n24107_;
  assign new_n24109_ = new_n23895_ & ~new_n24108_;
  assign new_n24110_ = ~new_n23894_ & new_n24109_;
  assign new_n24111_ = ~new_n24104_ & ~new_n24110_;
  assign new_n24112_ = ~\b[34]  & ~new_n24111_;
  assign new_n24113_ = ~new_n23332_ & ~\quotient[6] ;
  assign new_n24114_ = ~new_n23342_ & new_n23767_;
  assign new_n24115_ = ~new_n23763_ & new_n24114_;
  assign new_n24116_ = ~new_n23764_ & ~new_n23767_;
  assign new_n24117_ = ~new_n24115_ & ~new_n24116_;
  assign new_n24118_ = new_n23895_ & ~new_n24117_;
  assign new_n24119_ = ~new_n23894_ & new_n24118_;
  assign new_n24120_ = ~new_n24113_ & ~new_n24119_;
  assign new_n24121_ = ~\b[33]  & ~new_n24120_;
  assign new_n24122_ = ~new_n23341_ & ~\quotient[6] ;
  assign new_n24123_ = ~new_n23351_ & new_n23762_;
  assign new_n24124_ = ~new_n23758_ & new_n24123_;
  assign new_n24125_ = ~new_n23759_ & ~new_n23762_;
  assign new_n24126_ = ~new_n24124_ & ~new_n24125_;
  assign new_n24127_ = new_n23895_ & ~new_n24126_;
  assign new_n24128_ = ~new_n23894_ & new_n24127_;
  assign new_n24129_ = ~new_n24122_ & ~new_n24128_;
  assign new_n24130_ = ~\b[32]  & ~new_n24129_;
  assign new_n24131_ = ~new_n23350_ & ~\quotient[6] ;
  assign new_n24132_ = ~new_n23360_ & new_n23757_;
  assign new_n24133_ = ~new_n23753_ & new_n24132_;
  assign new_n24134_ = ~new_n23754_ & ~new_n23757_;
  assign new_n24135_ = ~new_n24133_ & ~new_n24134_;
  assign new_n24136_ = new_n23895_ & ~new_n24135_;
  assign new_n24137_ = ~new_n23894_ & new_n24136_;
  assign new_n24138_ = ~new_n24131_ & ~new_n24137_;
  assign new_n24139_ = ~\b[31]  & ~new_n24138_;
  assign new_n24140_ = ~new_n23359_ & ~\quotient[6] ;
  assign new_n24141_ = ~new_n23369_ & new_n23752_;
  assign new_n24142_ = ~new_n23748_ & new_n24141_;
  assign new_n24143_ = ~new_n23749_ & ~new_n23752_;
  assign new_n24144_ = ~new_n24142_ & ~new_n24143_;
  assign new_n24145_ = new_n23895_ & ~new_n24144_;
  assign new_n24146_ = ~new_n23894_ & new_n24145_;
  assign new_n24147_ = ~new_n24140_ & ~new_n24146_;
  assign new_n24148_ = ~\b[30]  & ~new_n24147_;
  assign new_n24149_ = ~new_n23368_ & ~\quotient[6] ;
  assign new_n24150_ = ~new_n23378_ & new_n23747_;
  assign new_n24151_ = ~new_n23743_ & new_n24150_;
  assign new_n24152_ = ~new_n23744_ & ~new_n23747_;
  assign new_n24153_ = ~new_n24151_ & ~new_n24152_;
  assign new_n24154_ = new_n23895_ & ~new_n24153_;
  assign new_n24155_ = ~new_n23894_ & new_n24154_;
  assign new_n24156_ = ~new_n24149_ & ~new_n24155_;
  assign new_n24157_ = ~\b[29]  & ~new_n24156_;
  assign new_n24158_ = ~new_n23377_ & ~\quotient[6] ;
  assign new_n24159_ = ~new_n23387_ & new_n23742_;
  assign new_n24160_ = ~new_n23738_ & new_n24159_;
  assign new_n24161_ = ~new_n23739_ & ~new_n23742_;
  assign new_n24162_ = ~new_n24160_ & ~new_n24161_;
  assign new_n24163_ = new_n23895_ & ~new_n24162_;
  assign new_n24164_ = ~new_n23894_ & new_n24163_;
  assign new_n24165_ = ~new_n24158_ & ~new_n24164_;
  assign new_n24166_ = ~\b[28]  & ~new_n24165_;
  assign new_n24167_ = ~new_n23386_ & ~\quotient[6] ;
  assign new_n24168_ = ~new_n23396_ & new_n23737_;
  assign new_n24169_ = ~new_n23733_ & new_n24168_;
  assign new_n24170_ = ~new_n23734_ & ~new_n23737_;
  assign new_n24171_ = ~new_n24169_ & ~new_n24170_;
  assign new_n24172_ = new_n23895_ & ~new_n24171_;
  assign new_n24173_ = ~new_n23894_ & new_n24172_;
  assign new_n24174_ = ~new_n24167_ & ~new_n24173_;
  assign new_n24175_ = ~\b[27]  & ~new_n24174_;
  assign new_n24176_ = ~new_n23395_ & ~\quotient[6] ;
  assign new_n24177_ = ~new_n23405_ & new_n23732_;
  assign new_n24178_ = ~new_n23728_ & new_n24177_;
  assign new_n24179_ = ~new_n23729_ & ~new_n23732_;
  assign new_n24180_ = ~new_n24178_ & ~new_n24179_;
  assign new_n24181_ = new_n23895_ & ~new_n24180_;
  assign new_n24182_ = ~new_n23894_ & new_n24181_;
  assign new_n24183_ = ~new_n24176_ & ~new_n24182_;
  assign new_n24184_ = ~\b[26]  & ~new_n24183_;
  assign new_n24185_ = ~new_n23404_ & ~\quotient[6] ;
  assign new_n24186_ = ~new_n23414_ & new_n23727_;
  assign new_n24187_ = ~new_n23723_ & new_n24186_;
  assign new_n24188_ = ~new_n23724_ & ~new_n23727_;
  assign new_n24189_ = ~new_n24187_ & ~new_n24188_;
  assign new_n24190_ = new_n23895_ & ~new_n24189_;
  assign new_n24191_ = ~new_n23894_ & new_n24190_;
  assign new_n24192_ = ~new_n24185_ & ~new_n24191_;
  assign new_n24193_ = ~\b[25]  & ~new_n24192_;
  assign new_n24194_ = ~new_n23413_ & ~\quotient[6] ;
  assign new_n24195_ = ~new_n23423_ & new_n23722_;
  assign new_n24196_ = ~new_n23718_ & new_n24195_;
  assign new_n24197_ = ~new_n23719_ & ~new_n23722_;
  assign new_n24198_ = ~new_n24196_ & ~new_n24197_;
  assign new_n24199_ = new_n23895_ & ~new_n24198_;
  assign new_n24200_ = ~new_n23894_ & new_n24199_;
  assign new_n24201_ = ~new_n24194_ & ~new_n24200_;
  assign new_n24202_ = ~\b[24]  & ~new_n24201_;
  assign new_n24203_ = ~new_n23422_ & ~\quotient[6] ;
  assign new_n24204_ = ~new_n23432_ & new_n23717_;
  assign new_n24205_ = ~new_n23713_ & new_n24204_;
  assign new_n24206_ = ~new_n23714_ & ~new_n23717_;
  assign new_n24207_ = ~new_n24205_ & ~new_n24206_;
  assign new_n24208_ = new_n23895_ & ~new_n24207_;
  assign new_n24209_ = ~new_n23894_ & new_n24208_;
  assign new_n24210_ = ~new_n24203_ & ~new_n24209_;
  assign new_n24211_ = ~\b[23]  & ~new_n24210_;
  assign new_n24212_ = ~new_n23431_ & ~\quotient[6] ;
  assign new_n24213_ = ~new_n23441_ & new_n23712_;
  assign new_n24214_ = ~new_n23708_ & new_n24213_;
  assign new_n24215_ = ~new_n23709_ & ~new_n23712_;
  assign new_n24216_ = ~new_n24214_ & ~new_n24215_;
  assign new_n24217_ = new_n23895_ & ~new_n24216_;
  assign new_n24218_ = ~new_n23894_ & new_n24217_;
  assign new_n24219_ = ~new_n24212_ & ~new_n24218_;
  assign new_n24220_ = ~\b[22]  & ~new_n24219_;
  assign new_n24221_ = ~new_n23440_ & ~\quotient[6] ;
  assign new_n24222_ = ~new_n23450_ & new_n23707_;
  assign new_n24223_ = ~new_n23703_ & new_n24222_;
  assign new_n24224_ = ~new_n23704_ & ~new_n23707_;
  assign new_n24225_ = ~new_n24223_ & ~new_n24224_;
  assign new_n24226_ = new_n23895_ & ~new_n24225_;
  assign new_n24227_ = ~new_n23894_ & new_n24226_;
  assign new_n24228_ = ~new_n24221_ & ~new_n24227_;
  assign new_n24229_ = ~\b[21]  & ~new_n24228_;
  assign new_n24230_ = ~new_n23449_ & ~\quotient[6] ;
  assign new_n24231_ = ~new_n23459_ & new_n23702_;
  assign new_n24232_ = ~new_n23698_ & new_n24231_;
  assign new_n24233_ = ~new_n23699_ & ~new_n23702_;
  assign new_n24234_ = ~new_n24232_ & ~new_n24233_;
  assign new_n24235_ = new_n23895_ & ~new_n24234_;
  assign new_n24236_ = ~new_n23894_ & new_n24235_;
  assign new_n24237_ = ~new_n24230_ & ~new_n24236_;
  assign new_n24238_ = ~\b[20]  & ~new_n24237_;
  assign new_n24239_ = ~new_n23458_ & ~\quotient[6] ;
  assign new_n24240_ = ~new_n23468_ & new_n23697_;
  assign new_n24241_ = ~new_n23693_ & new_n24240_;
  assign new_n24242_ = ~new_n23694_ & ~new_n23697_;
  assign new_n24243_ = ~new_n24241_ & ~new_n24242_;
  assign new_n24244_ = new_n23895_ & ~new_n24243_;
  assign new_n24245_ = ~new_n23894_ & new_n24244_;
  assign new_n24246_ = ~new_n24239_ & ~new_n24245_;
  assign new_n24247_ = ~\b[19]  & ~new_n24246_;
  assign new_n24248_ = ~new_n23467_ & ~\quotient[6] ;
  assign new_n24249_ = ~new_n23477_ & new_n23692_;
  assign new_n24250_ = ~new_n23688_ & new_n24249_;
  assign new_n24251_ = ~new_n23689_ & ~new_n23692_;
  assign new_n24252_ = ~new_n24250_ & ~new_n24251_;
  assign new_n24253_ = new_n23895_ & ~new_n24252_;
  assign new_n24254_ = ~new_n23894_ & new_n24253_;
  assign new_n24255_ = ~new_n24248_ & ~new_n24254_;
  assign new_n24256_ = ~\b[18]  & ~new_n24255_;
  assign new_n24257_ = ~new_n23476_ & ~\quotient[6] ;
  assign new_n24258_ = ~new_n23486_ & new_n23687_;
  assign new_n24259_ = ~new_n23683_ & new_n24258_;
  assign new_n24260_ = ~new_n23684_ & ~new_n23687_;
  assign new_n24261_ = ~new_n24259_ & ~new_n24260_;
  assign new_n24262_ = new_n23895_ & ~new_n24261_;
  assign new_n24263_ = ~new_n23894_ & new_n24262_;
  assign new_n24264_ = ~new_n24257_ & ~new_n24263_;
  assign new_n24265_ = ~\b[17]  & ~new_n24264_;
  assign new_n24266_ = ~new_n23485_ & ~\quotient[6] ;
  assign new_n24267_ = ~new_n23495_ & new_n23682_;
  assign new_n24268_ = ~new_n23678_ & new_n24267_;
  assign new_n24269_ = ~new_n23679_ & ~new_n23682_;
  assign new_n24270_ = ~new_n24268_ & ~new_n24269_;
  assign new_n24271_ = new_n23895_ & ~new_n24270_;
  assign new_n24272_ = ~new_n23894_ & new_n24271_;
  assign new_n24273_ = ~new_n24266_ & ~new_n24272_;
  assign new_n24274_ = ~\b[16]  & ~new_n24273_;
  assign new_n24275_ = ~new_n23494_ & ~\quotient[6] ;
  assign new_n24276_ = ~new_n23504_ & new_n23677_;
  assign new_n24277_ = ~new_n23673_ & new_n24276_;
  assign new_n24278_ = ~new_n23674_ & ~new_n23677_;
  assign new_n24279_ = ~new_n24277_ & ~new_n24278_;
  assign new_n24280_ = new_n23895_ & ~new_n24279_;
  assign new_n24281_ = ~new_n23894_ & new_n24280_;
  assign new_n24282_ = ~new_n24275_ & ~new_n24281_;
  assign new_n24283_ = ~\b[15]  & ~new_n24282_;
  assign new_n24284_ = ~new_n23503_ & ~\quotient[6] ;
  assign new_n24285_ = ~new_n23513_ & new_n23672_;
  assign new_n24286_ = ~new_n23668_ & new_n24285_;
  assign new_n24287_ = ~new_n23669_ & ~new_n23672_;
  assign new_n24288_ = ~new_n24286_ & ~new_n24287_;
  assign new_n24289_ = new_n23895_ & ~new_n24288_;
  assign new_n24290_ = ~new_n23894_ & new_n24289_;
  assign new_n24291_ = ~new_n24284_ & ~new_n24290_;
  assign new_n24292_ = ~\b[14]  & ~new_n24291_;
  assign new_n24293_ = ~new_n23512_ & ~\quotient[6] ;
  assign new_n24294_ = ~new_n23522_ & new_n23667_;
  assign new_n24295_ = ~new_n23663_ & new_n24294_;
  assign new_n24296_ = ~new_n23664_ & ~new_n23667_;
  assign new_n24297_ = ~new_n24295_ & ~new_n24296_;
  assign new_n24298_ = new_n23895_ & ~new_n24297_;
  assign new_n24299_ = ~new_n23894_ & new_n24298_;
  assign new_n24300_ = ~new_n24293_ & ~new_n24299_;
  assign new_n24301_ = ~\b[13]  & ~new_n24300_;
  assign new_n24302_ = ~new_n23521_ & ~\quotient[6] ;
  assign new_n24303_ = ~new_n23531_ & new_n23662_;
  assign new_n24304_ = ~new_n23658_ & new_n24303_;
  assign new_n24305_ = ~new_n23659_ & ~new_n23662_;
  assign new_n24306_ = ~new_n24304_ & ~new_n24305_;
  assign new_n24307_ = new_n23895_ & ~new_n24306_;
  assign new_n24308_ = ~new_n23894_ & new_n24307_;
  assign new_n24309_ = ~new_n24302_ & ~new_n24308_;
  assign new_n24310_ = ~\b[12]  & ~new_n24309_;
  assign new_n24311_ = ~new_n23530_ & ~\quotient[6] ;
  assign new_n24312_ = ~new_n23540_ & new_n23657_;
  assign new_n24313_ = ~new_n23653_ & new_n24312_;
  assign new_n24314_ = ~new_n23654_ & ~new_n23657_;
  assign new_n24315_ = ~new_n24313_ & ~new_n24314_;
  assign new_n24316_ = new_n23895_ & ~new_n24315_;
  assign new_n24317_ = ~new_n23894_ & new_n24316_;
  assign new_n24318_ = ~new_n24311_ & ~new_n24317_;
  assign new_n24319_ = ~\b[11]  & ~new_n24318_;
  assign new_n24320_ = ~new_n23539_ & ~\quotient[6] ;
  assign new_n24321_ = ~new_n23549_ & new_n23652_;
  assign new_n24322_ = ~new_n23648_ & new_n24321_;
  assign new_n24323_ = ~new_n23649_ & ~new_n23652_;
  assign new_n24324_ = ~new_n24322_ & ~new_n24323_;
  assign new_n24325_ = new_n23895_ & ~new_n24324_;
  assign new_n24326_ = ~new_n23894_ & new_n24325_;
  assign new_n24327_ = ~new_n24320_ & ~new_n24326_;
  assign new_n24328_ = ~\b[10]  & ~new_n24327_;
  assign new_n24329_ = ~new_n23548_ & ~\quotient[6] ;
  assign new_n24330_ = ~new_n23558_ & new_n23647_;
  assign new_n24331_ = ~new_n23643_ & new_n24330_;
  assign new_n24332_ = ~new_n23644_ & ~new_n23647_;
  assign new_n24333_ = ~new_n24331_ & ~new_n24332_;
  assign new_n24334_ = new_n23895_ & ~new_n24333_;
  assign new_n24335_ = ~new_n23894_ & new_n24334_;
  assign new_n24336_ = ~new_n24329_ & ~new_n24335_;
  assign new_n24337_ = ~\b[9]  & ~new_n24336_;
  assign new_n24338_ = ~new_n23557_ & ~\quotient[6] ;
  assign new_n24339_ = ~new_n23567_ & new_n23642_;
  assign new_n24340_ = ~new_n23638_ & new_n24339_;
  assign new_n24341_ = ~new_n23639_ & ~new_n23642_;
  assign new_n24342_ = ~new_n24340_ & ~new_n24341_;
  assign new_n24343_ = new_n23895_ & ~new_n24342_;
  assign new_n24344_ = ~new_n23894_ & new_n24343_;
  assign new_n24345_ = ~new_n24338_ & ~new_n24344_;
  assign new_n24346_ = ~\b[8]  & ~new_n24345_;
  assign new_n24347_ = ~new_n23566_ & ~\quotient[6] ;
  assign new_n24348_ = ~new_n23576_ & new_n23637_;
  assign new_n24349_ = ~new_n23633_ & new_n24348_;
  assign new_n24350_ = ~new_n23634_ & ~new_n23637_;
  assign new_n24351_ = ~new_n24349_ & ~new_n24350_;
  assign new_n24352_ = new_n23895_ & ~new_n24351_;
  assign new_n24353_ = ~new_n23894_ & new_n24352_;
  assign new_n24354_ = ~new_n24347_ & ~new_n24353_;
  assign new_n24355_ = ~\b[7]  & ~new_n24354_;
  assign new_n24356_ = ~new_n23575_ & ~\quotient[6] ;
  assign new_n24357_ = ~new_n23585_ & new_n23632_;
  assign new_n24358_ = ~new_n23628_ & new_n24357_;
  assign new_n24359_ = ~new_n23629_ & ~new_n23632_;
  assign new_n24360_ = ~new_n24358_ & ~new_n24359_;
  assign new_n24361_ = new_n23895_ & ~new_n24360_;
  assign new_n24362_ = ~new_n23894_ & new_n24361_;
  assign new_n24363_ = ~new_n24356_ & ~new_n24362_;
  assign new_n24364_ = ~\b[6]  & ~new_n24363_;
  assign new_n24365_ = ~new_n23584_ & ~\quotient[6] ;
  assign new_n24366_ = ~new_n23594_ & new_n23627_;
  assign new_n24367_ = ~new_n23623_ & new_n24366_;
  assign new_n24368_ = ~new_n23624_ & ~new_n23627_;
  assign new_n24369_ = ~new_n24367_ & ~new_n24368_;
  assign new_n24370_ = new_n23895_ & ~new_n24369_;
  assign new_n24371_ = ~new_n23894_ & new_n24370_;
  assign new_n24372_ = ~new_n24365_ & ~new_n24371_;
  assign new_n24373_ = ~\b[5]  & ~new_n24372_;
  assign new_n24374_ = ~new_n23593_ & ~\quotient[6] ;
  assign new_n24375_ = ~new_n23602_ & new_n23622_;
  assign new_n24376_ = ~new_n23618_ & new_n24375_;
  assign new_n24377_ = ~new_n23619_ & ~new_n23622_;
  assign new_n24378_ = ~new_n24376_ & ~new_n24377_;
  assign new_n24379_ = new_n23895_ & ~new_n24378_;
  assign new_n24380_ = ~new_n23894_ & new_n24379_;
  assign new_n24381_ = ~new_n24374_ & ~new_n24380_;
  assign new_n24382_ = ~\b[4]  & ~new_n24381_;
  assign new_n24383_ = ~new_n23601_ & ~\quotient[6] ;
  assign new_n24384_ = ~new_n23613_ & new_n23617_;
  assign new_n24385_ = ~new_n23612_ & new_n24384_;
  assign new_n24386_ = ~new_n23614_ & ~new_n23617_;
  assign new_n24387_ = ~new_n24385_ & ~new_n24386_;
  assign new_n24388_ = new_n23895_ & ~new_n24387_;
  assign new_n24389_ = ~new_n23894_ & new_n24388_;
  assign new_n24390_ = ~new_n24383_ & ~new_n24389_;
  assign new_n24391_ = ~\b[3]  & ~new_n24390_;
  assign new_n24392_ = ~new_n23606_ & ~\quotient[6] ;
  assign new_n24393_ = ~new_n23609_ & new_n23611_;
  assign new_n24394_ = ~new_n23607_ & new_n24393_;
  assign new_n24395_ = new_n23895_ & ~new_n24394_;
  assign new_n24396_ = ~new_n23612_ & new_n24395_;
  assign new_n24397_ = ~new_n23894_ & new_n24396_;
  assign new_n24398_ = ~new_n24392_ & ~new_n24397_;
  assign new_n24399_ = ~\b[2]  & ~new_n24398_;
  assign new_n24400_ = \b[0]  & ~\b[58] ;
  assign new_n24401_ = new_n405_ & new_n24400_;
  assign new_n24402_ = new_n403_ & new_n24401_;
  assign new_n24403_ = ~new_n23894_ & new_n24402_;
  assign new_n24404_ = \a[6]  & ~new_n24403_;
  assign new_n24405_ = new_n282_ & new_n23611_;
  assign new_n24406_ = new_n280_ & new_n24405_;
  assign new_n24407_ = ~new_n23894_ & new_n24406_;
  assign new_n24408_ = ~new_n24404_ & ~new_n24407_;
  assign new_n24409_ = \b[1]  & ~new_n24408_;
  assign new_n24410_ = ~\b[1]  & ~new_n24407_;
  assign new_n24411_ = ~new_n24404_ & new_n24410_;
  assign new_n24412_ = ~new_n24409_ & ~new_n24411_;
  assign new_n24413_ = ~\a[5]  & \b[0] ;
  assign new_n24414_ = ~new_n24412_ & ~new_n24413_;
  assign new_n24415_ = ~\b[1]  & ~new_n24408_;
  assign new_n24416_ = ~new_n24414_ & ~new_n24415_;
  assign new_n24417_ = \b[2]  & ~new_n24397_;
  assign new_n24418_ = ~new_n24392_ & new_n24417_;
  assign new_n24419_ = ~new_n24399_ & ~new_n24418_;
  assign new_n24420_ = ~new_n24416_ & new_n24419_;
  assign new_n24421_ = ~new_n24399_ & ~new_n24420_;
  assign new_n24422_ = \b[3]  & ~new_n24389_;
  assign new_n24423_ = ~new_n24383_ & new_n24422_;
  assign new_n24424_ = ~new_n24391_ & ~new_n24423_;
  assign new_n24425_ = ~new_n24421_ & new_n24424_;
  assign new_n24426_ = ~new_n24391_ & ~new_n24425_;
  assign new_n24427_ = \b[4]  & ~new_n24380_;
  assign new_n24428_ = ~new_n24374_ & new_n24427_;
  assign new_n24429_ = ~new_n24382_ & ~new_n24428_;
  assign new_n24430_ = ~new_n24426_ & new_n24429_;
  assign new_n24431_ = ~new_n24382_ & ~new_n24430_;
  assign new_n24432_ = \b[5]  & ~new_n24371_;
  assign new_n24433_ = ~new_n24365_ & new_n24432_;
  assign new_n24434_ = ~new_n24373_ & ~new_n24433_;
  assign new_n24435_ = ~new_n24431_ & new_n24434_;
  assign new_n24436_ = ~new_n24373_ & ~new_n24435_;
  assign new_n24437_ = \b[6]  & ~new_n24362_;
  assign new_n24438_ = ~new_n24356_ & new_n24437_;
  assign new_n24439_ = ~new_n24364_ & ~new_n24438_;
  assign new_n24440_ = ~new_n24436_ & new_n24439_;
  assign new_n24441_ = ~new_n24364_ & ~new_n24440_;
  assign new_n24442_ = \b[7]  & ~new_n24353_;
  assign new_n24443_ = ~new_n24347_ & new_n24442_;
  assign new_n24444_ = ~new_n24355_ & ~new_n24443_;
  assign new_n24445_ = ~new_n24441_ & new_n24444_;
  assign new_n24446_ = ~new_n24355_ & ~new_n24445_;
  assign new_n24447_ = \b[8]  & ~new_n24344_;
  assign new_n24448_ = ~new_n24338_ & new_n24447_;
  assign new_n24449_ = ~new_n24346_ & ~new_n24448_;
  assign new_n24450_ = ~new_n24446_ & new_n24449_;
  assign new_n24451_ = ~new_n24346_ & ~new_n24450_;
  assign new_n24452_ = \b[9]  & ~new_n24335_;
  assign new_n24453_ = ~new_n24329_ & new_n24452_;
  assign new_n24454_ = ~new_n24337_ & ~new_n24453_;
  assign new_n24455_ = ~new_n24451_ & new_n24454_;
  assign new_n24456_ = ~new_n24337_ & ~new_n24455_;
  assign new_n24457_ = \b[10]  & ~new_n24326_;
  assign new_n24458_ = ~new_n24320_ & new_n24457_;
  assign new_n24459_ = ~new_n24328_ & ~new_n24458_;
  assign new_n24460_ = ~new_n24456_ & new_n24459_;
  assign new_n24461_ = ~new_n24328_ & ~new_n24460_;
  assign new_n24462_ = \b[11]  & ~new_n24317_;
  assign new_n24463_ = ~new_n24311_ & new_n24462_;
  assign new_n24464_ = ~new_n24319_ & ~new_n24463_;
  assign new_n24465_ = ~new_n24461_ & new_n24464_;
  assign new_n24466_ = ~new_n24319_ & ~new_n24465_;
  assign new_n24467_ = \b[12]  & ~new_n24308_;
  assign new_n24468_ = ~new_n24302_ & new_n24467_;
  assign new_n24469_ = ~new_n24310_ & ~new_n24468_;
  assign new_n24470_ = ~new_n24466_ & new_n24469_;
  assign new_n24471_ = ~new_n24310_ & ~new_n24470_;
  assign new_n24472_ = \b[13]  & ~new_n24299_;
  assign new_n24473_ = ~new_n24293_ & new_n24472_;
  assign new_n24474_ = ~new_n24301_ & ~new_n24473_;
  assign new_n24475_ = ~new_n24471_ & new_n24474_;
  assign new_n24476_ = ~new_n24301_ & ~new_n24475_;
  assign new_n24477_ = \b[14]  & ~new_n24290_;
  assign new_n24478_ = ~new_n24284_ & new_n24477_;
  assign new_n24479_ = ~new_n24292_ & ~new_n24478_;
  assign new_n24480_ = ~new_n24476_ & new_n24479_;
  assign new_n24481_ = ~new_n24292_ & ~new_n24480_;
  assign new_n24482_ = \b[15]  & ~new_n24281_;
  assign new_n24483_ = ~new_n24275_ & new_n24482_;
  assign new_n24484_ = ~new_n24283_ & ~new_n24483_;
  assign new_n24485_ = ~new_n24481_ & new_n24484_;
  assign new_n24486_ = ~new_n24283_ & ~new_n24485_;
  assign new_n24487_ = \b[16]  & ~new_n24272_;
  assign new_n24488_ = ~new_n24266_ & new_n24487_;
  assign new_n24489_ = ~new_n24274_ & ~new_n24488_;
  assign new_n24490_ = ~new_n24486_ & new_n24489_;
  assign new_n24491_ = ~new_n24274_ & ~new_n24490_;
  assign new_n24492_ = \b[17]  & ~new_n24263_;
  assign new_n24493_ = ~new_n24257_ & new_n24492_;
  assign new_n24494_ = ~new_n24265_ & ~new_n24493_;
  assign new_n24495_ = ~new_n24491_ & new_n24494_;
  assign new_n24496_ = ~new_n24265_ & ~new_n24495_;
  assign new_n24497_ = \b[18]  & ~new_n24254_;
  assign new_n24498_ = ~new_n24248_ & new_n24497_;
  assign new_n24499_ = ~new_n24256_ & ~new_n24498_;
  assign new_n24500_ = ~new_n24496_ & new_n24499_;
  assign new_n24501_ = ~new_n24256_ & ~new_n24500_;
  assign new_n24502_ = \b[19]  & ~new_n24245_;
  assign new_n24503_ = ~new_n24239_ & new_n24502_;
  assign new_n24504_ = ~new_n24247_ & ~new_n24503_;
  assign new_n24505_ = ~new_n24501_ & new_n24504_;
  assign new_n24506_ = ~new_n24247_ & ~new_n24505_;
  assign new_n24507_ = \b[20]  & ~new_n24236_;
  assign new_n24508_ = ~new_n24230_ & new_n24507_;
  assign new_n24509_ = ~new_n24238_ & ~new_n24508_;
  assign new_n24510_ = ~new_n24506_ & new_n24509_;
  assign new_n24511_ = ~new_n24238_ & ~new_n24510_;
  assign new_n24512_ = \b[21]  & ~new_n24227_;
  assign new_n24513_ = ~new_n24221_ & new_n24512_;
  assign new_n24514_ = ~new_n24229_ & ~new_n24513_;
  assign new_n24515_ = ~new_n24511_ & new_n24514_;
  assign new_n24516_ = ~new_n24229_ & ~new_n24515_;
  assign new_n24517_ = \b[22]  & ~new_n24218_;
  assign new_n24518_ = ~new_n24212_ & new_n24517_;
  assign new_n24519_ = ~new_n24220_ & ~new_n24518_;
  assign new_n24520_ = ~new_n24516_ & new_n24519_;
  assign new_n24521_ = ~new_n24220_ & ~new_n24520_;
  assign new_n24522_ = \b[23]  & ~new_n24209_;
  assign new_n24523_ = ~new_n24203_ & new_n24522_;
  assign new_n24524_ = ~new_n24211_ & ~new_n24523_;
  assign new_n24525_ = ~new_n24521_ & new_n24524_;
  assign new_n24526_ = ~new_n24211_ & ~new_n24525_;
  assign new_n24527_ = \b[24]  & ~new_n24200_;
  assign new_n24528_ = ~new_n24194_ & new_n24527_;
  assign new_n24529_ = ~new_n24202_ & ~new_n24528_;
  assign new_n24530_ = ~new_n24526_ & new_n24529_;
  assign new_n24531_ = ~new_n24202_ & ~new_n24530_;
  assign new_n24532_ = \b[25]  & ~new_n24191_;
  assign new_n24533_ = ~new_n24185_ & new_n24532_;
  assign new_n24534_ = ~new_n24193_ & ~new_n24533_;
  assign new_n24535_ = ~new_n24531_ & new_n24534_;
  assign new_n24536_ = ~new_n24193_ & ~new_n24535_;
  assign new_n24537_ = \b[26]  & ~new_n24182_;
  assign new_n24538_ = ~new_n24176_ & new_n24537_;
  assign new_n24539_ = ~new_n24184_ & ~new_n24538_;
  assign new_n24540_ = ~new_n24536_ & new_n24539_;
  assign new_n24541_ = ~new_n24184_ & ~new_n24540_;
  assign new_n24542_ = \b[27]  & ~new_n24173_;
  assign new_n24543_ = ~new_n24167_ & new_n24542_;
  assign new_n24544_ = ~new_n24175_ & ~new_n24543_;
  assign new_n24545_ = ~new_n24541_ & new_n24544_;
  assign new_n24546_ = ~new_n24175_ & ~new_n24545_;
  assign new_n24547_ = \b[28]  & ~new_n24164_;
  assign new_n24548_ = ~new_n24158_ & new_n24547_;
  assign new_n24549_ = ~new_n24166_ & ~new_n24548_;
  assign new_n24550_ = ~new_n24546_ & new_n24549_;
  assign new_n24551_ = ~new_n24166_ & ~new_n24550_;
  assign new_n24552_ = \b[29]  & ~new_n24155_;
  assign new_n24553_ = ~new_n24149_ & new_n24552_;
  assign new_n24554_ = ~new_n24157_ & ~new_n24553_;
  assign new_n24555_ = ~new_n24551_ & new_n24554_;
  assign new_n24556_ = ~new_n24157_ & ~new_n24555_;
  assign new_n24557_ = \b[30]  & ~new_n24146_;
  assign new_n24558_ = ~new_n24140_ & new_n24557_;
  assign new_n24559_ = ~new_n24148_ & ~new_n24558_;
  assign new_n24560_ = ~new_n24556_ & new_n24559_;
  assign new_n24561_ = ~new_n24148_ & ~new_n24560_;
  assign new_n24562_ = \b[31]  & ~new_n24137_;
  assign new_n24563_ = ~new_n24131_ & new_n24562_;
  assign new_n24564_ = ~new_n24139_ & ~new_n24563_;
  assign new_n24565_ = ~new_n24561_ & new_n24564_;
  assign new_n24566_ = ~new_n24139_ & ~new_n24565_;
  assign new_n24567_ = \b[32]  & ~new_n24128_;
  assign new_n24568_ = ~new_n24122_ & new_n24567_;
  assign new_n24569_ = ~new_n24130_ & ~new_n24568_;
  assign new_n24570_ = ~new_n24566_ & new_n24569_;
  assign new_n24571_ = ~new_n24130_ & ~new_n24570_;
  assign new_n24572_ = \b[33]  & ~new_n24119_;
  assign new_n24573_ = ~new_n24113_ & new_n24572_;
  assign new_n24574_ = ~new_n24121_ & ~new_n24573_;
  assign new_n24575_ = ~new_n24571_ & new_n24574_;
  assign new_n24576_ = ~new_n24121_ & ~new_n24575_;
  assign new_n24577_ = \b[34]  & ~new_n24110_;
  assign new_n24578_ = ~new_n24104_ & new_n24577_;
  assign new_n24579_ = ~new_n24112_ & ~new_n24578_;
  assign new_n24580_ = ~new_n24576_ & new_n24579_;
  assign new_n24581_ = ~new_n24112_ & ~new_n24580_;
  assign new_n24582_ = \b[35]  & ~new_n24101_;
  assign new_n24583_ = ~new_n24095_ & new_n24582_;
  assign new_n24584_ = ~new_n24103_ & ~new_n24583_;
  assign new_n24585_ = ~new_n24581_ & new_n24584_;
  assign new_n24586_ = ~new_n24103_ & ~new_n24585_;
  assign new_n24587_ = \b[36]  & ~new_n24092_;
  assign new_n24588_ = ~new_n24086_ & new_n24587_;
  assign new_n24589_ = ~new_n24094_ & ~new_n24588_;
  assign new_n24590_ = ~new_n24586_ & new_n24589_;
  assign new_n24591_ = ~new_n24094_ & ~new_n24590_;
  assign new_n24592_ = \b[37]  & ~new_n24083_;
  assign new_n24593_ = ~new_n24077_ & new_n24592_;
  assign new_n24594_ = ~new_n24085_ & ~new_n24593_;
  assign new_n24595_ = ~new_n24591_ & new_n24594_;
  assign new_n24596_ = ~new_n24085_ & ~new_n24595_;
  assign new_n24597_ = \b[38]  & ~new_n24074_;
  assign new_n24598_ = ~new_n24068_ & new_n24597_;
  assign new_n24599_ = ~new_n24076_ & ~new_n24598_;
  assign new_n24600_ = ~new_n24596_ & new_n24599_;
  assign new_n24601_ = ~new_n24076_ & ~new_n24600_;
  assign new_n24602_ = \b[39]  & ~new_n24065_;
  assign new_n24603_ = ~new_n24059_ & new_n24602_;
  assign new_n24604_ = ~new_n24067_ & ~new_n24603_;
  assign new_n24605_ = ~new_n24601_ & new_n24604_;
  assign new_n24606_ = ~new_n24067_ & ~new_n24605_;
  assign new_n24607_ = \b[40]  & ~new_n24056_;
  assign new_n24608_ = ~new_n24050_ & new_n24607_;
  assign new_n24609_ = ~new_n24058_ & ~new_n24608_;
  assign new_n24610_ = ~new_n24606_ & new_n24609_;
  assign new_n24611_ = ~new_n24058_ & ~new_n24610_;
  assign new_n24612_ = \b[41]  & ~new_n24047_;
  assign new_n24613_ = ~new_n24041_ & new_n24612_;
  assign new_n24614_ = ~new_n24049_ & ~new_n24613_;
  assign new_n24615_ = ~new_n24611_ & new_n24614_;
  assign new_n24616_ = ~new_n24049_ & ~new_n24615_;
  assign new_n24617_ = \b[42]  & ~new_n24038_;
  assign new_n24618_ = ~new_n24032_ & new_n24617_;
  assign new_n24619_ = ~new_n24040_ & ~new_n24618_;
  assign new_n24620_ = ~new_n24616_ & new_n24619_;
  assign new_n24621_ = ~new_n24040_ & ~new_n24620_;
  assign new_n24622_ = \b[43]  & ~new_n24029_;
  assign new_n24623_ = ~new_n24023_ & new_n24622_;
  assign new_n24624_ = ~new_n24031_ & ~new_n24623_;
  assign new_n24625_ = ~new_n24621_ & new_n24624_;
  assign new_n24626_ = ~new_n24031_ & ~new_n24625_;
  assign new_n24627_ = \b[44]  & ~new_n24020_;
  assign new_n24628_ = ~new_n24014_ & new_n24627_;
  assign new_n24629_ = ~new_n24022_ & ~new_n24628_;
  assign new_n24630_ = ~new_n24626_ & new_n24629_;
  assign new_n24631_ = ~new_n24022_ & ~new_n24630_;
  assign new_n24632_ = \b[45]  & ~new_n24011_;
  assign new_n24633_ = ~new_n24005_ & new_n24632_;
  assign new_n24634_ = ~new_n24013_ & ~new_n24633_;
  assign new_n24635_ = ~new_n24631_ & new_n24634_;
  assign new_n24636_ = ~new_n24013_ & ~new_n24635_;
  assign new_n24637_ = \b[46]  & ~new_n24002_;
  assign new_n24638_ = ~new_n23996_ & new_n24637_;
  assign new_n24639_ = ~new_n24004_ & ~new_n24638_;
  assign new_n24640_ = ~new_n24636_ & new_n24639_;
  assign new_n24641_ = ~new_n24004_ & ~new_n24640_;
  assign new_n24642_ = \b[47]  & ~new_n23993_;
  assign new_n24643_ = ~new_n23987_ & new_n24642_;
  assign new_n24644_ = ~new_n23995_ & ~new_n24643_;
  assign new_n24645_ = ~new_n24641_ & new_n24644_;
  assign new_n24646_ = ~new_n23995_ & ~new_n24645_;
  assign new_n24647_ = \b[48]  & ~new_n23984_;
  assign new_n24648_ = ~new_n23978_ & new_n24647_;
  assign new_n24649_ = ~new_n23986_ & ~new_n24648_;
  assign new_n24650_ = ~new_n24646_ & new_n24649_;
  assign new_n24651_ = ~new_n23986_ & ~new_n24650_;
  assign new_n24652_ = \b[49]  & ~new_n23975_;
  assign new_n24653_ = ~new_n23969_ & new_n24652_;
  assign new_n24654_ = ~new_n23977_ & ~new_n24653_;
  assign new_n24655_ = ~new_n24651_ & new_n24654_;
  assign new_n24656_ = ~new_n23977_ & ~new_n24655_;
  assign new_n24657_ = \b[50]  & ~new_n23966_;
  assign new_n24658_ = ~new_n23960_ & new_n24657_;
  assign new_n24659_ = ~new_n23968_ & ~new_n24658_;
  assign new_n24660_ = ~new_n24656_ & new_n24659_;
  assign new_n24661_ = ~new_n23968_ & ~new_n24660_;
  assign new_n24662_ = \b[51]  & ~new_n23957_;
  assign new_n24663_ = ~new_n23951_ & new_n24662_;
  assign new_n24664_ = ~new_n23959_ & ~new_n24663_;
  assign new_n24665_ = ~new_n24661_ & new_n24664_;
  assign new_n24666_ = ~new_n23959_ & ~new_n24665_;
  assign new_n24667_ = \b[52]  & ~new_n23948_;
  assign new_n24668_ = ~new_n23942_ & new_n24667_;
  assign new_n24669_ = ~new_n23950_ & ~new_n24668_;
  assign new_n24670_ = ~new_n24666_ & new_n24669_;
  assign new_n24671_ = ~new_n23950_ & ~new_n24670_;
  assign new_n24672_ = \b[53]  & ~new_n23939_;
  assign new_n24673_ = ~new_n23933_ & new_n24672_;
  assign new_n24674_ = ~new_n23941_ & ~new_n24673_;
  assign new_n24675_ = ~new_n24671_ & new_n24674_;
  assign new_n24676_ = ~new_n23941_ & ~new_n24675_;
  assign new_n24677_ = \b[54]  & ~new_n23930_;
  assign new_n24678_ = ~new_n23924_ & new_n24677_;
  assign new_n24679_ = ~new_n23932_ & ~new_n24678_;
  assign new_n24680_ = ~new_n24676_ & new_n24679_;
  assign new_n24681_ = ~new_n23932_ & ~new_n24680_;
  assign new_n24682_ = \b[55]  & ~new_n23921_;
  assign new_n24683_ = ~new_n23915_ & new_n24682_;
  assign new_n24684_ = ~new_n23923_ & ~new_n24683_;
  assign new_n24685_ = ~new_n24681_ & new_n24684_;
  assign new_n24686_ = ~new_n23923_ & ~new_n24685_;
  assign new_n24687_ = \b[56]  & ~new_n23912_;
  assign new_n24688_ = ~new_n23906_ & new_n24687_;
  assign new_n24689_ = ~new_n23914_ & ~new_n24688_;
  assign new_n24690_ = ~new_n24686_ & new_n24689_;
  assign new_n24691_ = ~new_n23914_ & ~new_n24690_;
  assign new_n24692_ = \b[57]  & ~new_n23903_;
  assign new_n24693_ = ~new_n23897_ & new_n24692_;
  assign new_n24694_ = ~new_n23905_ & ~new_n24693_;
  assign new_n24695_ = ~new_n24691_ & new_n24694_;
  assign new_n24696_ = ~new_n23905_ & ~new_n24695_;
  assign new_n24697_ = ~new_n23115_ & ~\quotient[6] ;
  assign new_n24698_ = ~new_n23117_ & new_n23892_;
  assign new_n24699_ = ~new_n23888_ & new_n24698_;
  assign new_n24700_ = ~new_n23889_ & ~new_n23892_;
  assign new_n24701_ = ~new_n24699_ & ~new_n24700_;
  assign new_n24702_ = \quotient[6]  & ~new_n24701_;
  assign new_n24703_ = ~new_n24697_ & ~new_n24702_;
  assign new_n24704_ = ~\b[58]  & ~new_n24703_;
  assign new_n24705_ = \b[58]  & ~new_n24697_;
  assign new_n24706_ = ~new_n24702_ & new_n24705_;
  assign new_n24707_ = new_n403_ & new_n405_;
  assign new_n24708_ = ~new_n24706_ & new_n24707_;
  assign new_n24709_ = ~new_n24704_ & new_n24708_;
  assign new_n24710_ = ~new_n24696_ & new_n24709_;
  assign new_n24711_ = new_n23895_ & ~new_n24703_;
  assign \quotient[5]  = new_n24710_ | new_n24711_;
  assign new_n24713_ = ~new_n23914_ & new_n24694_;
  assign new_n24714_ = ~new_n24690_ & new_n24713_;
  assign new_n24715_ = ~new_n24691_ & ~new_n24694_;
  assign new_n24716_ = ~new_n24714_ & ~new_n24715_;
  assign new_n24717_ = \quotient[5]  & ~new_n24716_;
  assign new_n24718_ = ~new_n23904_ & ~new_n24711_;
  assign new_n24719_ = ~new_n24710_ & new_n24718_;
  assign new_n24720_ = ~new_n24717_ & ~new_n24719_;
  assign new_n24721_ = ~\b[58]  & ~new_n24720_;
  assign new_n24722_ = ~new_n23923_ & new_n24689_;
  assign new_n24723_ = ~new_n24685_ & new_n24722_;
  assign new_n24724_ = ~new_n24686_ & ~new_n24689_;
  assign new_n24725_ = ~new_n24723_ & ~new_n24724_;
  assign new_n24726_ = \quotient[5]  & ~new_n24725_;
  assign new_n24727_ = ~new_n23913_ & ~new_n24711_;
  assign new_n24728_ = ~new_n24710_ & new_n24727_;
  assign new_n24729_ = ~new_n24726_ & ~new_n24728_;
  assign new_n24730_ = ~\b[57]  & ~new_n24729_;
  assign new_n24731_ = ~new_n23932_ & new_n24684_;
  assign new_n24732_ = ~new_n24680_ & new_n24731_;
  assign new_n24733_ = ~new_n24681_ & ~new_n24684_;
  assign new_n24734_ = ~new_n24732_ & ~new_n24733_;
  assign new_n24735_ = \quotient[5]  & ~new_n24734_;
  assign new_n24736_ = ~new_n23922_ & ~new_n24711_;
  assign new_n24737_ = ~new_n24710_ & new_n24736_;
  assign new_n24738_ = ~new_n24735_ & ~new_n24737_;
  assign new_n24739_ = ~\b[56]  & ~new_n24738_;
  assign new_n24740_ = ~new_n23941_ & new_n24679_;
  assign new_n24741_ = ~new_n24675_ & new_n24740_;
  assign new_n24742_ = ~new_n24676_ & ~new_n24679_;
  assign new_n24743_ = ~new_n24741_ & ~new_n24742_;
  assign new_n24744_ = \quotient[5]  & ~new_n24743_;
  assign new_n24745_ = ~new_n23931_ & ~new_n24711_;
  assign new_n24746_ = ~new_n24710_ & new_n24745_;
  assign new_n24747_ = ~new_n24744_ & ~new_n24746_;
  assign new_n24748_ = ~\b[55]  & ~new_n24747_;
  assign new_n24749_ = ~new_n23950_ & new_n24674_;
  assign new_n24750_ = ~new_n24670_ & new_n24749_;
  assign new_n24751_ = ~new_n24671_ & ~new_n24674_;
  assign new_n24752_ = ~new_n24750_ & ~new_n24751_;
  assign new_n24753_ = \quotient[5]  & ~new_n24752_;
  assign new_n24754_ = ~new_n23940_ & ~new_n24711_;
  assign new_n24755_ = ~new_n24710_ & new_n24754_;
  assign new_n24756_ = ~new_n24753_ & ~new_n24755_;
  assign new_n24757_ = ~\b[54]  & ~new_n24756_;
  assign new_n24758_ = ~new_n23959_ & new_n24669_;
  assign new_n24759_ = ~new_n24665_ & new_n24758_;
  assign new_n24760_ = ~new_n24666_ & ~new_n24669_;
  assign new_n24761_ = ~new_n24759_ & ~new_n24760_;
  assign new_n24762_ = \quotient[5]  & ~new_n24761_;
  assign new_n24763_ = ~new_n23949_ & ~new_n24711_;
  assign new_n24764_ = ~new_n24710_ & new_n24763_;
  assign new_n24765_ = ~new_n24762_ & ~new_n24764_;
  assign new_n24766_ = ~\b[53]  & ~new_n24765_;
  assign new_n24767_ = ~new_n23968_ & new_n24664_;
  assign new_n24768_ = ~new_n24660_ & new_n24767_;
  assign new_n24769_ = ~new_n24661_ & ~new_n24664_;
  assign new_n24770_ = ~new_n24768_ & ~new_n24769_;
  assign new_n24771_ = \quotient[5]  & ~new_n24770_;
  assign new_n24772_ = ~new_n23958_ & ~new_n24711_;
  assign new_n24773_ = ~new_n24710_ & new_n24772_;
  assign new_n24774_ = ~new_n24771_ & ~new_n24773_;
  assign new_n24775_ = ~\b[52]  & ~new_n24774_;
  assign new_n24776_ = ~new_n23977_ & new_n24659_;
  assign new_n24777_ = ~new_n24655_ & new_n24776_;
  assign new_n24778_ = ~new_n24656_ & ~new_n24659_;
  assign new_n24779_ = ~new_n24777_ & ~new_n24778_;
  assign new_n24780_ = \quotient[5]  & ~new_n24779_;
  assign new_n24781_ = ~new_n23967_ & ~new_n24711_;
  assign new_n24782_ = ~new_n24710_ & new_n24781_;
  assign new_n24783_ = ~new_n24780_ & ~new_n24782_;
  assign new_n24784_ = ~\b[51]  & ~new_n24783_;
  assign new_n24785_ = ~new_n23986_ & new_n24654_;
  assign new_n24786_ = ~new_n24650_ & new_n24785_;
  assign new_n24787_ = ~new_n24651_ & ~new_n24654_;
  assign new_n24788_ = ~new_n24786_ & ~new_n24787_;
  assign new_n24789_ = \quotient[5]  & ~new_n24788_;
  assign new_n24790_ = ~new_n23976_ & ~new_n24711_;
  assign new_n24791_ = ~new_n24710_ & new_n24790_;
  assign new_n24792_ = ~new_n24789_ & ~new_n24791_;
  assign new_n24793_ = ~\b[50]  & ~new_n24792_;
  assign new_n24794_ = ~new_n23995_ & new_n24649_;
  assign new_n24795_ = ~new_n24645_ & new_n24794_;
  assign new_n24796_ = ~new_n24646_ & ~new_n24649_;
  assign new_n24797_ = ~new_n24795_ & ~new_n24796_;
  assign new_n24798_ = \quotient[5]  & ~new_n24797_;
  assign new_n24799_ = ~new_n23985_ & ~new_n24711_;
  assign new_n24800_ = ~new_n24710_ & new_n24799_;
  assign new_n24801_ = ~new_n24798_ & ~new_n24800_;
  assign new_n24802_ = ~\b[49]  & ~new_n24801_;
  assign new_n24803_ = ~new_n24004_ & new_n24644_;
  assign new_n24804_ = ~new_n24640_ & new_n24803_;
  assign new_n24805_ = ~new_n24641_ & ~new_n24644_;
  assign new_n24806_ = ~new_n24804_ & ~new_n24805_;
  assign new_n24807_ = \quotient[5]  & ~new_n24806_;
  assign new_n24808_ = ~new_n23994_ & ~new_n24711_;
  assign new_n24809_ = ~new_n24710_ & new_n24808_;
  assign new_n24810_ = ~new_n24807_ & ~new_n24809_;
  assign new_n24811_ = ~\b[48]  & ~new_n24810_;
  assign new_n24812_ = ~new_n24013_ & new_n24639_;
  assign new_n24813_ = ~new_n24635_ & new_n24812_;
  assign new_n24814_ = ~new_n24636_ & ~new_n24639_;
  assign new_n24815_ = ~new_n24813_ & ~new_n24814_;
  assign new_n24816_ = \quotient[5]  & ~new_n24815_;
  assign new_n24817_ = ~new_n24003_ & ~new_n24711_;
  assign new_n24818_ = ~new_n24710_ & new_n24817_;
  assign new_n24819_ = ~new_n24816_ & ~new_n24818_;
  assign new_n24820_ = ~\b[47]  & ~new_n24819_;
  assign new_n24821_ = ~new_n24022_ & new_n24634_;
  assign new_n24822_ = ~new_n24630_ & new_n24821_;
  assign new_n24823_ = ~new_n24631_ & ~new_n24634_;
  assign new_n24824_ = ~new_n24822_ & ~new_n24823_;
  assign new_n24825_ = \quotient[5]  & ~new_n24824_;
  assign new_n24826_ = ~new_n24012_ & ~new_n24711_;
  assign new_n24827_ = ~new_n24710_ & new_n24826_;
  assign new_n24828_ = ~new_n24825_ & ~new_n24827_;
  assign new_n24829_ = ~\b[46]  & ~new_n24828_;
  assign new_n24830_ = ~new_n24031_ & new_n24629_;
  assign new_n24831_ = ~new_n24625_ & new_n24830_;
  assign new_n24832_ = ~new_n24626_ & ~new_n24629_;
  assign new_n24833_ = ~new_n24831_ & ~new_n24832_;
  assign new_n24834_ = \quotient[5]  & ~new_n24833_;
  assign new_n24835_ = ~new_n24021_ & ~new_n24711_;
  assign new_n24836_ = ~new_n24710_ & new_n24835_;
  assign new_n24837_ = ~new_n24834_ & ~new_n24836_;
  assign new_n24838_ = ~\b[45]  & ~new_n24837_;
  assign new_n24839_ = ~new_n24040_ & new_n24624_;
  assign new_n24840_ = ~new_n24620_ & new_n24839_;
  assign new_n24841_ = ~new_n24621_ & ~new_n24624_;
  assign new_n24842_ = ~new_n24840_ & ~new_n24841_;
  assign new_n24843_ = \quotient[5]  & ~new_n24842_;
  assign new_n24844_ = ~new_n24030_ & ~new_n24711_;
  assign new_n24845_ = ~new_n24710_ & new_n24844_;
  assign new_n24846_ = ~new_n24843_ & ~new_n24845_;
  assign new_n24847_ = ~\b[44]  & ~new_n24846_;
  assign new_n24848_ = ~new_n24049_ & new_n24619_;
  assign new_n24849_ = ~new_n24615_ & new_n24848_;
  assign new_n24850_ = ~new_n24616_ & ~new_n24619_;
  assign new_n24851_ = ~new_n24849_ & ~new_n24850_;
  assign new_n24852_ = \quotient[5]  & ~new_n24851_;
  assign new_n24853_ = ~new_n24039_ & ~new_n24711_;
  assign new_n24854_ = ~new_n24710_ & new_n24853_;
  assign new_n24855_ = ~new_n24852_ & ~new_n24854_;
  assign new_n24856_ = ~\b[43]  & ~new_n24855_;
  assign new_n24857_ = ~new_n24058_ & new_n24614_;
  assign new_n24858_ = ~new_n24610_ & new_n24857_;
  assign new_n24859_ = ~new_n24611_ & ~new_n24614_;
  assign new_n24860_ = ~new_n24858_ & ~new_n24859_;
  assign new_n24861_ = \quotient[5]  & ~new_n24860_;
  assign new_n24862_ = ~new_n24048_ & ~new_n24711_;
  assign new_n24863_ = ~new_n24710_ & new_n24862_;
  assign new_n24864_ = ~new_n24861_ & ~new_n24863_;
  assign new_n24865_ = ~\b[42]  & ~new_n24864_;
  assign new_n24866_ = ~new_n24067_ & new_n24609_;
  assign new_n24867_ = ~new_n24605_ & new_n24866_;
  assign new_n24868_ = ~new_n24606_ & ~new_n24609_;
  assign new_n24869_ = ~new_n24867_ & ~new_n24868_;
  assign new_n24870_ = \quotient[5]  & ~new_n24869_;
  assign new_n24871_ = ~new_n24057_ & ~new_n24711_;
  assign new_n24872_ = ~new_n24710_ & new_n24871_;
  assign new_n24873_ = ~new_n24870_ & ~new_n24872_;
  assign new_n24874_ = ~\b[41]  & ~new_n24873_;
  assign new_n24875_ = ~new_n24076_ & new_n24604_;
  assign new_n24876_ = ~new_n24600_ & new_n24875_;
  assign new_n24877_ = ~new_n24601_ & ~new_n24604_;
  assign new_n24878_ = ~new_n24876_ & ~new_n24877_;
  assign new_n24879_ = \quotient[5]  & ~new_n24878_;
  assign new_n24880_ = ~new_n24066_ & ~new_n24711_;
  assign new_n24881_ = ~new_n24710_ & new_n24880_;
  assign new_n24882_ = ~new_n24879_ & ~new_n24881_;
  assign new_n24883_ = ~\b[40]  & ~new_n24882_;
  assign new_n24884_ = ~new_n24085_ & new_n24599_;
  assign new_n24885_ = ~new_n24595_ & new_n24884_;
  assign new_n24886_ = ~new_n24596_ & ~new_n24599_;
  assign new_n24887_ = ~new_n24885_ & ~new_n24886_;
  assign new_n24888_ = \quotient[5]  & ~new_n24887_;
  assign new_n24889_ = ~new_n24075_ & ~new_n24711_;
  assign new_n24890_ = ~new_n24710_ & new_n24889_;
  assign new_n24891_ = ~new_n24888_ & ~new_n24890_;
  assign new_n24892_ = ~\b[39]  & ~new_n24891_;
  assign new_n24893_ = ~new_n24094_ & new_n24594_;
  assign new_n24894_ = ~new_n24590_ & new_n24893_;
  assign new_n24895_ = ~new_n24591_ & ~new_n24594_;
  assign new_n24896_ = ~new_n24894_ & ~new_n24895_;
  assign new_n24897_ = \quotient[5]  & ~new_n24896_;
  assign new_n24898_ = ~new_n24084_ & ~new_n24711_;
  assign new_n24899_ = ~new_n24710_ & new_n24898_;
  assign new_n24900_ = ~new_n24897_ & ~new_n24899_;
  assign new_n24901_ = ~\b[38]  & ~new_n24900_;
  assign new_n24902_ = ~new_n24103_ & new_n24589_;
  assign new_n24903_ = ~new_n24585_ & new_n24902_;
  assign new_n24904_ = ~new_n24586_ & ~new_n24589_;
  assign new_n24905_ = ~new_n24903_ & ~new_n24904_;
  assign new_n24906_ = \quotient[5]  & ~new_n24905_;
  assign new_n24907_ = ~new_n24093_ & ~new_n24711_;
  assign new_n24908_ = ~new_n24710_ & new_n24907_;
  assign new_n24909_ = ~new_n24906_ & ~new_n24908_;
  assign new_n24910_ = ~\b[37]  & ~new_n24909_;
  assign new_n24911_ = ~new_n24112_ & new_n24584_;
  assign new_n24912_ = ~new_n24580_ & new_n24911_;
  assign new_n24913_ = ~new_n24581_ & ~new_n24584_;
  assign new_n24914_ = ~new_n24912_ & ~new_n24913_;
  assign new_n24915_ = \quotient[5]  & ~new_n24914_;
  assign new_n24916_ = ~new_n24102_ & ~new_n24711_;
  assign new_n24917_ = ~new_n24710_ & new_n24916_;
  assign new_n24918_ = ~new_n24915_ & ~new_n24917_;
  assign new_n24919_ = ~\b[36]  & ~new_n24918_;
  assign new_n24920_ = ~new_n24121_ & new_n24579_;
  assign new_n24921_ = ~new_n24575_ & new_n24920_;
  assign new_n24922_ = ~new_n24576_ & ~new_n24579_;
  assign new_n24923_ = ~new_n24921_ & ~new_n24922_;
  assign new_n24924_ = \quotient[5]  & ~new_n24923_;
  assign new_n24925_ = ~new_n24111_ & ~new_n24711_;
  assign new_n24926_ = ~new_n24710_ & new_n24925_;
  assign new_n24927_ = ~new_n24924_ & ~new_n24926_;
  assign new_n24928_ = ~\b[35]  & ~new_n24927_;
  assign new_n24929_ = ~new_n24130_ & new_n24574_;
  assign new_n24930_ = ~new_n24570_ & new_n24929_;
  assign new_n24931_ = ~new_n24571_ & ~new_n24574_;
  assign new_n24932_ = ~new_n24930_ & ~new_n24931_;
  assign new_n24933_ = \quotient[5]  & ~new_n24932_;
  assign new_n24934_ = ~new_n24120_ & ~new_n24711_;
  assign new_n24935_ = ~new_n24710_ & new_n24934_;
  assign new_n24936_ = ~new_n24933_ & ~new_n24935_;
  assign new_n24937_ = ~\b[34]  & ~new_n24936_;
  assign new_n24938_ = ~new_n24139_ & new_n24569_;
  assign new_n24939_ = ~new_n24565_ & new_n24938_;
  assign new_n24940_ = ~new_n24566_ & ~new_n24569_;
  assign new_n24941_ = ~new_n24939_ & ~new_n24940_;
  assign new_n24942_ = \quotient[5]  & ~new_n24941_;
  assign new_n24943_ = ~new_n24129_ & ~new_n24711_;
  assign new_n24944_ = ~new_n24710_ & new_n24943_;
  assign new_n24945_ = ~new_n24942_ & ~new_n24944_;
  assign new_n24946_ = ~\b[33]  & ~new_n24945_;
  assign new_n24947_ = ~new_n24148_ & new_n24564_;
  assign new_n24948_ = ~new_n24560_ & new_n24947_;
  assign new_n24949_ = ~new_n24561_ & ~new_n24564_;
  assign new_n24950_ = ~new_n24948_ & ~new_n24949_;
  assign new_n24951_ = \quotient[5]  & ~new_n24950_;
  assign new_n24952_ = ~new_n24138_ & ~new_n24711_;
  assign new_n24953_ = ~new_n24710_ & new_n24952_;
  assign new_n24954_ = ~new_n24951_ & ~new_n24953_;
  assign new_n24955_ = ~\b[32]  & ~new_n24954_;
  assign new_n24956_ = ~new_n24157_ & new_n24559_;
  assign new_n24957_ = ~new_n24555_ & new_n24956_;
  assign new_n24958_ = ~new_n24556_ & ~new_n24559_;
  assign new_n24959_ = ~new_n24957_ & ~new_n24958_;
  assign new_n24960_ = \quotient[5]  & ~new_n24959_;
  assign new_n24961_ = ~new_n24147_ & ~new_n24711_;
  assign new_n24962_ = ~new_n24710_ & new_n24961_;
  assign new_n24963_ = ~new_n24960_ & ~new_n24962_;
  assign new_n24964_ = ~\b[31]  & ~new_n24963_;
  assign new_n24965_ = ~new_n24166_ & new_n24554_;
  assign new_n24966_ = ~new_n24550_ & new_n24965_;
  assign new_n24967_ = ~new_n24551_ & ~new_n24554_;
  assign new_n24968_ = ~new_n24966_ & ~new_n24967_;
  assign new_n24969_ = \quotient[5]  & ~new_n24968_;
  assign new_n24970_ = ~new_n24156_ & ~new_n24711_;
  assign new_n24971_ = ~new_n24710_ & new_n24970_;
  assign new_n24972_ = ~new_n24969_ & ~new_n24971_;
  assign new_n24973_ = ~\b[30]  & ~new_n24972_;
  assign new_n24974_ = ~new_n24175_ & new_n24549_;
  assign new_n24975_ = ~new_n24545_ & new_n24974_;
  assign new_n24976_ = ~new_n24546_ & ~new_n24549_;
  assign new_n24977_ = ~new_n24975_ & ~new_n24976_;
  assign new_n24978_ = \quotient[5]  & ~new_n24977_;
  assign new_n24979_ = ~new_n24165_ & ~new_n24711_;
  assign new_n24980_ = ~new_n24710_ & new_n24979_;
  assign new_n24981_ = ~new_n24978_ & ~new_n24980_;
  assign new_n24982_ = ~\b[29]  & ~new_n24981_;
  assign new_n24983_ = ~new_n24184_ & new_n24544_;
  assign new_n24984_ = ~new_n24540_ & new_n24983_;
  assign new_n24985_ = ~new_n24541_ & ~new_n24544_;
  assign new_n24986_ = ~new_n24984_ & ~new_n24985_;
  assign new_n24987_ = \quotient[5]  & ~new_n24986_;
  assign new_n24988_ = ~new_n24174_ & ~new_n24711_;
  assign new_n24989_ = ~new_n24710_ & new_n24988_;
  assign new_n24990_ = ~new_n24987_ & ~new_n24989_;
  assign new_n24991_ = ~\b[28]  & ~new_n24990_;
  assign new_n24992_ = ~new_n24193_ & new_n24539_;
  assign new_n24993_ = ~new_n24535_ & new_n24992_;
  assign new_n24994_ = ~new_n24536_ & ~new_n24539_;
  assign new_n24995_ = ~new_n24993_ & ~new_n24994_;
  assign new_n24996_ = \quotient[5]  & ~new_n24995_;
  assign new_n24997_ = ~new_n24183_ & ~new_n24711_;
  assign new_n24998_ = ~new_n24710_ & new_n24997_;
  assign new_n24999_ = ~new_n24996_ & ~new_n24998_;
  assign new_n25000_ = ~\b[27]  & ~new_n24999_;
  assign new_n25001_ = ~new_n24202_ & new_n24534_;
  assign new_n25002_ = ~new_n24530_ & new_n25001_;
  assign new_n25003_ = ~new_n24531_ & ~new_n24534_;
  assign new_n25004_ = ~new_n25002_ & ~new_n25003_;
  assign new_n25005_ = \quotient[5]  & ~new_n25004_;
  assign new_n25006_ = ~new_n24192_ & ~new_n24711_;
  assign new_n25007_ = ~new_n24710_ & new_n25006_;
  assign new_n25008_ = ~new_n25005_ & ~new_n25007_;
  assign new_n25009_ = ~\b[26]  & ~new_n25008_;
  assign new_n25010_ = ~new_n24211_ & new_n24529_;
  assign new_n25011_ = ~new_n24525_ & new_n25010_;
  assign new_n25012_ = ~new_n24526_ & ~new_n24529_;
  assign new_n25013_ = ~new_n25011_ & ~new_n25012_;
  assign new_n25014_ = \quotient[5]  & ~new_n25013_;
  assign new_n25015_ = ~new_n24201_ & ~new_n24711_;
  assign new_n25016_ = ~new_n24710_ & new_n25015_;
  assign new_n25017_ = ~new_n25014_ & ~new_n25016_;
  assign new_n25018_ = ~\b[25]  & ~new_n25017_;
  assign new_n25019_ = ~new_n24220_ & new_n24524_;
  assign new_n25020_ = ~new_n24520_ & new_n25019_;
  assign new_n25021_ = ~new_n24521_ & ~new_n24524_;
  assign new_n25022_ = ~new_n25020_ & ~new_n25021_;
  assign new_n25023_ = \quotient[5]  & ~new_n25022_;
  assign new_n25024_ = ~new_n24210_ & ~new_n24711_;
  assign new_n25025_ = ~new_n24710_ & new_n25024_;
  assign new_n25026_ = ~new_n25023_ & ~new_n25025_;
  assign new_n25027_ = ~\b[24]  & ~new_n25026_;
  assign new_n25028_ = ~new_n24229_ & new_n24519_;
  assign new_n25029_ = ~new_n24515_ & new_n25028_;
  assign new_n25030_ = ~new_n24516_ & ~new_n24519_;
  assign new_n25031_ = ~new_n25029_ & ~new_n25030_;
  assign new_n25032_ = \quotient[5]  & ~new_n25031_;
  assign new_n25033_ = ~new_n24219_ & ~new_n24711_;
  assign new_n25034_ = ~new_n24710_ & new_n25033_;
  assign new_n25035_ = ~new_n25032_ & ~new_n25034_;
  assign new_n25036_ = ~\b[23]  & ~new_n25035_;
  assign new_n25037_ = ~new_n24238_ & new_n24514_;
  assign new_n25038_ = ~new_n24510_ & new_n25037_;
  assign new_n25039_ = ~new_n24511_ & ~new_n24514_;
  assign new_n25040_ = ~new_n25038_ & ~new_n25039_;
  assign new_n25041_ = \quotient[5]  & ~new_n25040_;
  assign new_n25042_ = ~new_n24228_ & ~new_n24711_;
  assign new_n25043_ = ~new_n24710_ & new_n25042_;
  assign new_n25044_ = ~new_n25041_ & ~new_n25043_;
  assign new_n25045_ = ~\b[22]  & ~new_n25044_;
  assign new_n25046_ = ~new_n24247_ & new_n24509_;
  assign new_n25047_ = ~new_n24505_ & new_n25046_;
  assign new_n25048_ = ~new_n24506_ & ~new_n24509_;
  assign new_n25049_ = ~new_n25047_ & ~new_n25048_;
  assign new_n25050_ = \quotient[5]  & ~new_n25049_;
  assign new_n25051_ = ~new_n24237_ & ~new_n24711_;
  assign new_n25052_ = ~new_n24710_ & new_n25051_;
  assign new_n25053_ = ~new_n25050_ & ~new_n25052_;
  assign new_n25054_ = ~\b[21]  & ~new_n25053_;
  assign new_n25055_ = ~new_n24256_ & new_n24504_;
  assign new_n25056_ = ~new_n24500_ & new_n25055_;
  assign new_n25057_ = ~new_n24501_ & ~new_n24504_;
  assign new_n25058_ = ~new_n25056_ & ~new_n25057_;
  assign new_n25059_ = \quotient[5]  & ~new_n25058_;
  assign new_n25060_ = ~new_n24246_ & ~new_n24711_;
  assign new_n25061_ = ~new_n24710_ & new_n25060_;
  assign new_n25062_ = ~new_n25059_ & ~new_n25061_;
  assign new_n25063_ = ~\b[20]  & ~new_n25062_;
  assign new_n25064_ = ~new_n24265_ & new_n24499_;
  assign new_n25065_ = ~new_n24495_ & new_n25064_;
  assign new_n25066_ = ~new_n24496_ & ~new_n24499_;
  assign new_n25067_ = ~new_n25065_ & ~new_n25066_;
  assign new_n25068_ = \quotient[5]  & ~new_n25067_;
  assign new_n25069_ = ~new_n24255_ & ~new_n24711_;
  assign new_n25070_ = ~new_n24710_ & new_n25069_;
  assign new_n25071_ = ~new_n25068_ & ~new_n25070_;
  assign new_n25072_ = ~\b[19]  & ~new_n25071_;
  assign new_n25073_ = ~new_n24274_ & new_n24494_;
  assign new_n25074_ = ~new_n24490_ & new_n25073_;
  assign new_n25075_ = ~new_n24491_ & ~new_n24494_;
  assign new_n25076_ = ~new_n25074_ & ~new_n25075_;
  assign new_n25077_ = \quotient[5]  & ~new_n25076_;
  assign new_n25078_ = ~new_n24264_ & ~new_n24711_;
  assign new_n25079_ = ~new_n24710_ & new_n25078_;
  assign new_n25080_ = ~new_n25077_ & ~new_n25079_;
  assign new_n25081_ = ~\b[18]  & ~new_n25080_;
  assign new_n25082_ = ~new_n24283_ & new_n24489_;
  assign new_n25083_ = ~new_n24485_ & new_n25082_;
  assign new_n25084_ = ~new_n24486_ & ~new_n24489_;
  assign new_n25085_ = ~new_n25083_ & ~new_n25084_;
  assign new_n25086_ = \quotient[5]  & ~new_n25085_;
  assign new_n25087_ = ~new_n24273_ & ~new_n24711_;
  assign new_n25088_ = ~new_n24710_ & new_n25087_;
  assign new_n25089_ = ~new_n25086_ & ~new_n25088_;
  assign new_n25090_ = ~\b[17]  & ~new_n25089_;
  assign new_n25091_ = ~new_n24292_ & new_n24484_;
  assign new_n25092_ = ~new_n24480_ & new_n25091_;
  assign new_n25093_ = ~new_n24481_ & ~new_n24484_;
  assign new_n25094_ = ~new_n25092_ & ~new_n25093_;
  assign new_n25095_ = \quotient[5]  & ~new_n25094_;
  assign new_n25096_ = ~new_n24282_ & ~new_n24711_;
  assign new_n25097_ = ~new_n24710_ & new_n25096_;
  assign new_n25098_ = ~new_n25095_ & ~new_n25097_;
  assign new_n25099_ = ~\b[16]  & ~new_n25098_;
  assign new_n25100_ = ~new_n24301_ & new_n24479_;
  assign new_n25101_ = ~new_n24475_ & new_n25100_;
  assign new_n25102_ = ~new_n24476_ & ~new_n24479_;
  assign new_n25103_ = ~new_n25101_ & ~new_n25102_;
  assign new_n25104_ = \quotient[5]  & ~new_n25103_;
  assign new_n25105_ = ~new_n24291_ & ~new_n24711_;
  assign new_n25106_ = ~new_n24710_ & new_n25105_;
  assign new_n25107_ = ~new_n25104_ & ~new_n25106_;
  assign new_n25108_ = ~\b[15]  & ~new_n25107_;
  assign new_n25109_ = ~new_n24310_ & new_n24474_;
  assign new_n25110_ = ~new_n24470_ & new_n25109_;
  assign new_n25111_ = ~new_n24471_ & ~new_n24474_;
  assign new_n25112_ = ~new_n25110_ & ~new_n25111_;
  assign new_n25113_ = \quotient[5]  & ~new_n25112_;
  assign new_n25114_ = ~new_n24300_ & ~new_n24711_;
  assign new_n25115_ = ~new_n24710_ & new_n25114_;
  assign new_n25116_ = ~new_n25113_ & ~new_n25115_;
  assign new_n25117_ = ~\b[14]  & ~new_n25116_;
  assign new_n25118_ = ~new_n24319_ & new_n24469_;
  assign new_n25119_ = ~new_n24465_ & new_n25118_;
  assign new_n25120_ = ~new_n24466_ & ~new_n24469_;
  assign new_n25121_ = ~new_n25119_ & ~new_n25120_;
  assign new_n25122_ = \quotient[5]  & ~new_n25121_;
  assign new_n25123_ = ~new_n24309_ & ~new_n24711_;
  assign new_n25124_ = ~new_n24710_ & new_n25123_;
  assign new_n25125_ = ~new_n25122_ & ~new_n25124_;
  assign new_n25126_ = ~\b[13]  & ~new_n25125_;
  assign new_n25127_ = ~new_n24328_ & new_n24464_;
  assign new_n25128_ = ~new_n24460_ & new_n25127_;
  assign new_n25129_ = ~new_n24461_ & ~new_n24464_;
  assign new_n25130_ = ~new_n25128_ & ~new_n25129_;
  assign new_n25131_ = \quotient[5]  & ~new_n25130_;
  assign new_n25132_ = ~new_n24318_ & ~new_n24711_;
  assign new_n25133_ = ~new_n24710_ & new_n25132_;
  assign new_n25134_ = ~new_n25131_ & ~new_n25133_;
  assign new_n25135_ = ~\b[12]  & ~new_n25134_;
  assign new_n25136_ = ~new_n24337_ & new_n24459_;
  assign new_n25137_ = ~new_n24455_ & new_n25136_;
  assign new_n25138_ = ~new_n24456_ & ~new_n24459_;
  assign new_n25139_ = ~new_n25137_ & ~new_n25138_;
  assign new_n25140_ = \quotient[5]  & ~new_n25139_;
  assign new_n25141_ = ~new_n24327_ & ~new_n24711_;
  assign new_n25142_ = ~new_n24710_ & new_n25141_;
  assign new_n25143_ = ~new_n25140_ & ~new_n25142_;
  assign new_n25144_ = ~\b[11]  & ~new_n25143_;
  assign new_n25145_ = ~new_n24346_ & new_n24454_;
  assign new_n25146_ = ~new_n24450_ & new_n25145_;
  assign new_n25147_ = ~new_n24451_ & ~new_n24454_;
  assign new_n25148_ = ~new_n25146_ & ~new_n25147_;
  assign new_n25149_ = \quotient[5]  & ~new_n25148_;
  assign new_n25150_ = ~new_n24336_ & ~new_n24711_;
  assign new_n25151_ = ~new_n24710_ & new_n25150_;
  assign new_n25152_ = ~new_n25149_ & ~new_n25151_;
  assign new_n25153_ = ~\b[10]  & ~new_n25152_;
  assign new_n25154_ = ~new_n24355_ & new_n24449_;
  assign new_n25155_ = ~new_n24445_ & new_n25154_;
  assign new_n25156_ = ~new_n24446_ & ~new_n24449_;
  assign new_n25157_ = ~new_n25155_ & ~new_n25156_;
  assign new_n25158_ = \quotient[5]  & ~new_n25157_;
  assign new_n25159_ = ~new_n24345_ & ~new_n24711_;
  assign new_n25160_ = ~new_n24710_ & new_n25159_;
  assign new_n25161_ = ~new_n25158_ & ~new_n25160_;
  assign new_n25162_ = ~\b[9]  & ~new_n25161_;
  assign new_n25163_ = ~new_n24364_ & new_n24444_;
  assign new_n25164_ = ~new_n24440_ & new_n25163_;
  assign new_n25165_ = ~new_n24441_ & ~new_n24444_;
  assign new_n25166_ = ~new_n25164_ & ~new_n25165_;
  assign new_n25167_ = \quotient[5]  & ~new_n25166_;
  assign new_n25168_ = ~new_n24354_ & ~new_n24711_;
  assign new_n25169_ = ~new_n24710_ & new_n25168_;
  assign new_n25170_ = ~new_n25167_ & ~new_n25169_;
  assign new_n25171_ = ~\b[8]  & ~new_n25170_;
  assign new_n25172_ = ~new_n24373_ & new_n24439_;
  assign new_n25173_ = ~new_n24435_ & new_n25172_;
  assign new_n25174_ = ~new_n24436_ & ~new_n24439_;
  assign new_n25175_ = ~new_n25173_ & ~new_n25174_;
  assign new_n25176_ = \quotient[5]  & ~new_n25175_;
  assign new_n25177_ = ~new_n24363_ & ~new_n24711_;
  assign new_n25178_ = ~new_n24710_ & new_n25177_;
  assign new_n25179_ = ~new_n25176_ & ~new_n25178_;
  assign new_n25180_ = ~\b[7]  & ~new_n25179_;
  assign new_n25181_ = ~new_n24382_ & new_n24434_;
  assign new_n25182_ = ~new_n24430_ & new_n25181_;
  assign new_n25183_ = ~new_n24431_ & ~new_n24434_;
  assign new_n25184_ = ~new_n25182_ & ~new_n25183_;
  assign new_n25185_ = \quotient[5]  & ~new_n25184_;
  assign new_n25186_ = ~new_n24372_ & ~new_n24711_;
  assign new_n25187_ = ~new_n24710_ & new_n25186_;
  assign new_n25188_ = ~new_n25185_ & ~new_n25187_;
  assign new_n25189_ = ~\b[6]  & ~new_n25188_;
  assign new_n25190_ = ~new_n24391_ & new_n24429_;
  assign new_n25191_ = ~new_n24425_ & new_n25190_;
  assign new_n25192_ = ~new_n24426_ & ~new_n24429_;
  assign new_n25193_ = ~new_n25191_ & ~new_n25192_;
  assign new_n25194_ = \quotient[5]  & ~new_n25193_;
  assign new_n25195_ = ~new_n24381_ & ~new_n24711_;
  assign new_n25196_ = ~new_n24710_ & new_n25195_;
  assign new_n25197_ = ~new_n25194_ & ~new_n25196_;
  assign new_n25198_ = ~\b[5]  & ~new_n25197_;
  assign new_n25199_ = ~new_n24399_ & new_n24424_;
  assign new_n25200_ = ~new_n24420_ & new_n25199_;
  assign new_n25201_ = ~new_n24421_ & ~new_n24424_;
  assign new_n25202_ = ~new_n25200_ & ~new_n25201_;
  assign new_n25203_ = \quotient[5]  & ~new_n25202_;
  assign new_n25204_ = ~new_n24390_ & ~new_n24711_;
  assign new_n25205_ = ~new_n24710_ & new_n25204_;
  assign new_n25206_ = ~new_n25203_ & ~new_n25205_;
  assign new_n25207_ = ~\b[4]  & ~new_n25206_;
  assign new_n25208_ = ~new_n24415_ & new_n24419_;
  assign new_n25209_ = ~new_n24414_ & new_n25208_;
  assign new_n25210_ = ~new_n24416_ & ~new_n24419_;
  assign new_n25211_ = ~new_n25209_ & ~new_n25210_;
  assign new_n25212_ = \quotient[5]  & ~new_n25211_;
  assign new_n25213_ = ~new_n24398_ & ~new_n24711_;
  assign new_n25214_ = ~new_n24710_ & new_n25213_;
  assign new_n25215_ = ~new_n25212_ & ~new_n25214_;
  assign new_n25216_ = ~\b[3]  & ~new_n25215_;
  assign new_n25217_ = ~new_n24411_ & new_n24413_;
  assign new_n25218_ = ~new_n24409_ & new_n25217_;
  assign new_n25219_ = ~new_n24414_ & ~new_n25218_;
  assign new_n25220_ = \quotient[5]  & new_n25219_;
  assign new_n25221_ = ~new_n24408_ & ~new_n24711_;
  assign new_n25222_ = ~new_n24710_ & new_n25221_;
  assign new_n25223_ = ~new_n25220_ & ~new_n25222_;
  assign new_n25224_ = ~\b[2]  & ~new_n25223_;
  assign new_n25225_ = \b[0]  & \quotient[5] ;
  assign new_n25226_ = \a[5]  & ~new_n25225_;
  assign new_n25227_ = new_n24413_ & \quotient[5] ;
  assign new_n25228_ = ~new_n25226_ & ~new_n25227_;
  assign new_n25229_ = \b[1]  & ~new_n25228_;
  assign new_n25230_ = ~\b[1]  & ~new_n25227_;
  assign new_n25231_ = ~new_n25226_ & new_n25230_;
  assign new_n25232_ = ~new_n25229_ & ~new_n25231_;
  assign new_n25233_ = ~\a[4]  & \b[0] ;
  assign new_n25234_ = ~new_n25232_ & ~new_n25233_;
  assign new_n25235_ = ~\b[1]  & ~new_n25228_;
  assign new_n25236_ = ~new_n25234_ & ~new_n25235_;
  assign new_n25237_ = \b[2]  & ~new_n25222_;
  assign new_n25238_ = ~new_n25220_ & new_n25237_;
  assign new_n25239_ = ~new_n25224_ & ~new_n25238_;
  assign new_n25240_ = ~new_n25236_ & new_n25239_;
  assign new_n25241_ = ~new_n25224_ & ~new_n25240_;
  assign new_n25242_ = \b[3]  & ~new_n25214_;
  assign new_n25243_ = ~new_n25212_ & new_n25242_;
  assign new_n25244_ = ~new_n25216_ & ~new_n25243_;
  assign new_n25245_ = ~new_n25241_ & new_n25244_;
  assign new_n25246_ = ~new_n25216_ & ~new_n25245_;
  assign new_n25247_ = \b[4]  & ~new_n25205_;
  assign new_n25248_ = ~new_n25203_ & new_n25247_;
  assign new_n25249_ = ~new_n25207_ & ~new_n25248_;
  assign new_n25250_ = ~new_n25246_ & new_n25249_;
  assign new_n25251_ = ~new_n25207_ & ~new_n25250_;
  assign new_n25252_ = \b[5]  & ~new_n25196_;
  assign new_n25253_ = ~new_n25194_ & new_n25252_;
  assign new_n25254_ = ~new_n25198_ & ~new_n25253_;
  assign new_n25255_ = ~new_n25251_ & new_n25254_;
  assign new_n25256_ = ~new_n25198_ & ~new_n25255_;
  assign new_n25257_ = \b[6]  & ~new_n25187_;
  assign new_n25258_ = ~new_n25185_ & new_n25257_;
  assign new_n25259_ = ~new_n25189_ & ~new_n25258_;
  assign new_n25260_ = ~new_n25256_ & new_n25259_;
  assign new_n25261_ = ~new_n25189_ & ~new_n25260_;
  assign new_n25262_ = \b[7]  & ~new_n25178_;
  assign new_n25263_ = ~new_n25176_ & new_n25262_;
  assign new_n25264_ = ~new_n25180_ & ~new_n25263_;
  assign new_n25265_ = ~new_n25261_ & new_n25264_;
  assign new_n25266_ = ~new_n25180_ & ~new_n25265_;
  assign new_n25267_ = \b[8]  & ~new_n25169_;
  assign new_n25268_ = ~new_n25167_ & new_n25267_;
  assign new_n25269_ = ~new_n25171_ & ~new_n25268_;
  assign new_n25270_ = ~new_n25266_ & new_n25269_;
  assign new_n25271_ = ~new_n25171_ & ~new_n25270_;
  assign new_n25272_ = \b[9]  & ~new_n25160_;
  assign new_n25273_ = ~new_n25158_ & new_n25272_;
  assign new_n25274_ = ~new_n25162_ & ~new_n25273_;
  assign new_n25275_ = ~new_n25271_ & new_n25274_;
  assign new_n25276_ = ~new_n25162_ & ~new_n25275_;
  assign new_n25277_ = \b[10]  & ~new_n25151_;
  assign new_n25278_ = ~new_n25149_ & new_n25277_;
  assign new_n25279_ = ~new_n25153_ & ~new_n25278_;
  assign new_n25280_ = ~new_n25276_ & new_n25279_;
  assign new_n25281_ = ~new_n25153_ & ~new_n25280_;
  assign new_n25282_ = \b[11]  & ~new_n25142_;
  assign new_n25283_ = ~new_n25140_ & new_n25282_;
  assign new_n25284_ = ~new_n25144_ & ~new_n25283_;
  assign new_n25285_ = ~new_n25281_ & new_n25284_;
  assign new_n25286_ = ~new_n25144_ & ~new_n25285_;
  assign new_n25287_ = \b[12]  & ~new_n25133_;
  assign new_n25288_ = ~new_n25131_ & new_n25287_;
  assign new_n25289_ = ~new_n25135_ & ~new_n25288_;
  assign new_n25290_ = ~new_n25286_ & new_n25289_;
  assign new_n25291_ = ~new_n25135_ & ~new_n25290_;
  assign new_n25292_ = \b[13]  & ~new_n25124_;
  assign new_n25293_ = ~new_n25122_ & new_n25292_;
  assign new_n25294_ = ~new_n25126_ & ~new_n25293_;
  assign new_n25295_ = ~new_n25291_ & new_n25294_;
  assign new_n25296_ = ~new_n25126_ & ~new_n25295_;
  assign new_n25297_ = \b[14]  & ~new_n25115_;
  assign new_n25298_ = ~new_n25113_ & new_n25297_;
  assign new_n25299_ = ~new_n25117_ & ~new_n25298_;
  assign new_n25300_ = ~new_n25296_ & new_n25299_;
  assign new_n25301_ = ~new_n25117_ & ~new_n25300_;
  assign new_n25302_ = \b[15]  & ~new_n25106_;
  assign new_n25303_ = ~new_n25104_ & new_n25302_;
  assign new_n25304_ = ~new_n25108_ & ~new_n25303_;
  assign new_n25305_ = ~new_n25301_ & new_n25304_;
  assign new_n25306_ = ~new_n25108_ & ~new_n25305_;
  assign new_n25307_ = \b[16]  & ~new_n25097_;
  assign new_n25308_ = ~new_n25095_ & new_n25307_;
  assign new_n25309_ = ~new_n25099_ & ~new_n25308_;
  assign new_n25310_ = ~new_n25306_ & new_n25309_;
  assign new_n25311_ = ~new_n25099_ & ~new_n25310_;
  assign new_n25312_ = \b[17]  & ~new_n25088_;
  assign new_n25313_ = ~new_n25086_ & new_n25312_;
  assign new_n25314_ = ~new_n25090_ & ~new_n25313_;
  assign new_n25315_ = ~new_n25311_ & new_n25314_;
  assign new_n25316_ = ~new_n25090_ & ~new_n25315_;
  assign new_n25317_ = \b[18]  & ~new_n25079_;
  assign new_n25318_ = ~new_n25077_ & new_n25317_;
  assign new_n25319_ = ~new_n25081_ & ~new_n25318_;
  assign new_n25320_ = ~new_n25316_ & new_n25319_;
  assign new_n25321_ = ~new_n25081_ & ~new_n25320_;
  assign new_n25322_ = \b[19]  & ~new_n25070_;
  assign new_n25323_ = ~new_n25068_ & new_n25322_;
  assign new_n25324_ = ~new_n25072_ & ~new_n25323_;
  assign new_n25325_ = ~new_n25321_ & new_n25324_;
  assign new_n25326_ = ~new_n25072_ & ~new_n25325_;
  assign new_n25327_ = \b[20]  & ~new_n25061_;
  assign new_n25328_ = ~new_n25059_ & new_n25327_;
  assign new_n25329_ = ~new_n25063_ & ~new_n25328_;
  assign new_n25330_ = ~new_n25326_ & new_n25329_;
  assign new_n25331_ = ~new_n25063_ & ~new_n25330_;
  assign new_n25332_ = \b[21]  & ~new_n25052_;
  assign new_n25333_ = ~new_n25050_ & new_n25332_;
  assign new_n25334_ = ~new_n25054_ & ~new_n25333_;
  assign new_n25335_ = ~new_n25331_ & new_n25334_;
  assign new_n25336_ = ~new_n25054_ & ~new_n25335_;
  assign new_n25337_ = \b[22]  & ~new_n25043_;
  assign new_n25338_ = ~new_n25041_ & new_n25337_;
  assign new_n25339_ = ~new_n25045_ & ~new_n25338_;
  assign new_n25340_ = ~new_n25336_ & new_n25339_;
  assign new_n25341_ = ~new_n25045_ & ~new_n25340_;
  assign new_n25342_ = \b[23]  & ~new_n25034_;
  assign new_n25343_ = ~new_n25032_ & new_n25342_;
  assign new_n25344_ = ~new_n25036_ & ~new_n25343_;
  assign new_n25345_ = ~new_n25341_ & new_n25344_;
  assign new_n25346_ = ~new_n25036_ & ~new_n25345_;
  assign new_n25347_ = \b[24]  & ~new_n25025_;
  assign new_n25348_ = ~new_n25023_ & new_n25347_;
  assign new_n25349_ = ~new_n25027_ & ~new_n25348_;
  assign new_n25350_ = ~new_n25346_ & new_n25349_;
  assign new_n25351_ = ~new_n25027_ & ~new_n25350_;
  assign new_n25352_ = \b[25]  & ~new_n25016_;
  assign new_n25353_ = ~new_n25014_ & new_n25352_;
  assign new_n25354_ = ~new_n25018_ & ~new_n25353_;
  assign new_n25355_ = ~new_n25351_ & new_n25354_;
  assign new_n25356_ = ~new_n25018_ & ~new_n25355_;
  assign new_n25357_ = \b[26]  & ~new_n25007_;
  assign new_n25358_ = ~new_n25005_ & new_n25357_;
  assign new_n25359_ = ~new_n25009_ & ~new_n25358_;
  assign new_n25360_ = ~new_n25356_ & new_n25359_;
  assign new_n25361_ = ~new_n25009_ & ~new_n25360_;
  assign new_n25362_ = \b[27]  & ~new_n24998_;
  assign new_n25363_ = ~new_n24996_ & new_n25362_;
  assign new_n25364_ = ~new_n25000_ & ~new_n25363_;
  assign new_n25365_ = ~new_n25361_ & new_n25364_;
  assign new_n25366_ = ~new_n25000_ & ~new_n25365_;
  assign new_n25367_ = \b[28]  & ~new_n24989_;
  assign new_n25368_ = ~new_n24987_ & new_n25367_;
  assign new_n25369_ = ~new_n24991_ & ~new_n25368_;
  assign new_n25370_ = ~new_n25366_ & new_n25369_;
  assign new_n25371_ = ~new_n24991_ & ~new_n25370_;
  assign new_n25372_ = \b[29]  & ~new_n24980_;
  assign new_n25373_ = ~new_n24978_ & new_n25372_;
  assign new_n25374_ = ~new_n24982_ & ~new_n25373_;
  assign new_n25375_ = ~new_n25371_ & new_n25374_;
  assign new_n25376_ = ~new_n24982_ & ~new_n25375_;
  assign new_n25377_ = \b[30]  & ~new_n24971_;
  assign new_n25378_ = ~new_n24969_ & new_n25377_;
  assign new_n25379_ = ~new_n24973_ & ~new_n25378_;
  assign new_n25380_ = ~new_n25376_ & new_n25379_;
  assign new_n25381_ = ~new_n24973_ & ~new_n25380_;
  assign new_n25382_ = \b[31]  & ~new_n24962_;
  assign new_n25383_ = ~new_n24960_ & new_n25382_;
  assign new_n25384_ = ~new_n24964_ & ~new_n25383_;
  assign new_n25385_ = ~new_n25381_ & new_n25384_;
  assign new_n25386_ = ~new_n24964_ & ~new_n25385_;
  assign new_n25387_ = \b[32]  & ~new_n24953_;
  assign new_n25388_ = ~new_n24951_ & new_n25387_;
  assign new_n25389_ = ~new_n24955_ & ~new_n25388_;
  assign new_n25390_ = ~new_n25386_ & new_n25389_;
  assign new_n25391_ = ~new_n24955_ & ~new_n25390_;
  assign new_n25392_ = \b[33]  & ~new_n24944_;
  assign new_n25393_ = ~new_n24942_ & new_n25392_;
  assign new_n25394_ = ~new_n24946_ & ~new_n25393_;
  assign new_n25395_ = ~new_n25391_ & new_n25394_;
  assign new_n25396_ = ~new_n24946_ & ~new_n25395_;
  assign new_n25397_ = \b[34]  & ~new_n24935_;
  assign new_n25398_ = ~new_n24933_ & new_n25397_;
  assign new_n25399_ = ~new_n24937_ & ~new_n25398_;
  assign new_n25400_ = ~new_n25396_ & new_n25399_;
  assign new_n25401_ = ~new_n24937_ & ~new_n25400_;
  assign new_n25402_ = \b[35]  & ~new_n24926_;
  assign new_n25403_ = ~new_n24924_ & new_n25402_;
  assign new_n25404_ = ~new_n24928_ & ~new_n25403_;
  assign new_n25405_ = ~new_n25401_ & new_n25404_;
  assign new_n25406_ = ~new_n24928_ & ~new_n25405_;
  assign new_n25407_ = \b[36]  & ~new_n24917_;
  assign new_n25408_ = ~new_n24915_ & new_n25407_;
  assign new_n25409_ = ~new_n24919_ & ~new_n25408_;
  assign new_n25410_ = ~new_n25406_ & new_n25409_;
  assign new_n25411_ = ~new_n24919_ & ~new_n25410_;
  assign new_n25412_ = \b[37]  & ~new_n24908_;
  assign new_n25413_ = ~new_n24906_ & new_n25412_;
  assign new_n25414_ = ~new_n24910_ & ~new_n25413_;
  assign new_n25415_ = ~new_n25411_ & new_n25414_;
  assign new_n25416_ = ~new_n24910_ & ~new_n25415_;
  assign new_n25417_ = \b[38]  & ~new_n24899_;
  assign new_n25418_ = ~new_n24897_ & new_n25417_;
  assign new_n25419_ = ~new_n24901_ & ~new_n25418_;
  assign new_n25420_ = ~new_n25416_ & new_n25419_;
  assign new_n25421_ = ~new_n24901_ & ~new_n25420_;
  assign new_n25422_ = \b[39]  & ~new_n24890_;
  assign new_n25423_ = ~new_n24888_ & new_n25422_;
  assign new_n25424_ = ~new_n24892_ & ~new_n25423_;
  assign new_n25425_ = ~new_n25421_ & new_n25424_;
  assign new_n25426_ = ~new_n24892_ & ~new_n25425_;
  assign new_n25427_ = \b[40]  & ~new_n24881_;
  assign new_n25428_ = ~new_n24879_ & new_n25427_;
  assign new_n25429_ = ~new_n24883_ & ~new_n25428_;
  assign new_n25430_ = ~new_n25426_ & new_n25429_;
  assign new_n25431_ = ~new_n24883_ & ~new_n25430_;
  assign new_n25432_ = \b[41]  & ~new_n24872_;
  assign new_n25433_ = ~new_n24870_ & new_n25432_;
  assign new_n25434_ = ~new_n24874_ & ~new_n25433_;
  assign new_n25435_ = ~new_n25431_ & new_n25434_;
  assign new_n25436_ = ~new_n24874_ & ~new_n25435_;
  assign new_n25437_ = \b[42]  & ~new_n24863_;
  assign new_n25438_ = ~new_n24861_ & new_n25437_;
  assign new_n25439_ = ~new_n24865_ & ~new_n25438_;
  assign new_n25440_ = ~new_n25436_ & new_n25439_;
  assign new_n25441_ = ~new_n24865_ & ~new_n25440_;
  assign new_n25442_ = \b[43]  & ~new_n24854_;
  assign new_n25443_ = ~new_n24852_ & new_n25442_;
  assign new_n25444_ = ~new_n24856_ & ~new_n25443_;
  assign new_n25445_ = ~new_n25441_ & new_n25444_;
  assign new_n25446_ = ~new_n24856_ & ~new_n25445_;
  assign new_n25447_ = \b[44]  & ~new_n24845_;
  assign new_n25448_ = ~new_n24843_ & new_n25447_;
  assign new_n25449_ = ~new_n24847_ & ~new_n25448_;
  assign new_n25450_ = ~new_n25446_ & new_n25449_;
  assign new_n25451_ = ~new_n24847_ & ~new_n25450_;
  assign new_n25452_ = \b[45]  & ~new_n24836_;
  assign new_n25453_ = ~new_n24834_ & new_n25452_;
  assign new_n25454_ = ~new_n24838_ & ~new_n25453_;
  assign new_n25455_ = ~new_n25451_ & new_n25454_;
  assign new_n25456_ = ~new_n24838_ & ~new_n25455_;
  assign new_n25457_ = \b[46]  & ~new_n24827_;
  assign new_n25458_ = ~new_n24825_ & new_n25457_;
  assign new_n25459_ = ~new_n24829_ & ~new_n25458_;
  assign new_n25460_ = ~new_n25456_ & new_n25459_;
  assign new_n25461_ = ~new_n24829_ & ~new_n25460_;
  assign new_n25462_ = \b[47]  & ~new_n24818_;
  assign new_n25463_ = ~new_n24816_ & new_n25462_;
  assign new_n25464_ = ~new_n24820_ & ~new_n25463_;
  assign new_n25465_ = ~new_n25461_ & new_n25464_;
  assign new_n25466_ = ~new_n24820_ & ~new_n25465_;
  assign new_n25467_ = \b[48]  & ~new_n24809_;
  assign new_n25468_ = ~new_n24807_ & new_n25467_;
  assign new_n25469_ = ~new_n24811_ & ~new_n25468_;
  assign new_n25470_ = ~new_n25466_ & new_n25469_;
  assign new_n25471_ = ~new_n24811_ & ~new_n25470_;
  assign new_n25472_ = \b[49]  & ~new_n24800_;
  assign new_n25473_ = ~new_n24798_ & new_n25472_;
  assign new_n25474_ = ~new_n24802_ & ~new_n25473_;
  assign new_n25475_ = ~new_n25471_ & new_n25474_;
  assign new_n25476_ = ~new_n24802_ & ~new_n25475_;
  assign new_n25477_ = \b[50]  & ~new_n24791_;
  assign new_n25478_ = ~new_n24789_ & new_n25477_;
  assign new_n25479_ = ~new_n24793_ & ~new_n25478_;
  assign new_n25480_ = ~new_n25476_ & new_n25479_;
  assign new_n25481_ = ~new_n24793_ & ~new_n25480_;
  assign new_n25482_ = \b[51]  & ~new_n24782_;
  assign new_n25483_ = ~new_n24780_ & new_n25482_;
  assign new_n25484_ = ~new_n24784_ & ~new_n25483_;
  assign new_n25485_ = ~new_n25481_ & new_n25484_;
  assign new_n25486_ = ~new_n24784_ & ~new_n25485_;
  assign new_n25487_ = \b[52]  & ~new_n24773_;
  assign new_n25488_ = ~new_n24771_ & new_n25487_;
  assign new_n25489_ = ~new_n24775_ & ~new_n25488_;
  assign new_n25490_ = ~new_n25486_ & new_n25489_;
  assign new_n25491_ = ~new_n24775_ & ~new_n25490_;
  assign new_n25492_ = \b[53]  & ~new_n24764_;
  assign new_n25493_ = ~new_n24762_ & new_n25492_;
  assign new_n25494_ = ~new_n24766_ & ~new_n25493_;
  assign new_n25495_ = ~new_n25491_ & new_n25494_;
  assign new_n25496_ = ~new_n24766_ & ~new_n25495_;
  assign new_n25497_ = \b[54]  & ~new_n24755_;
  assign new_n25498_ = ~new_n24753_ & new_n25497_;
  assign new_n25499_ = ~new_n24757_ & ~new_n25498_;
  assign new_n25500_ = ~new_n25496_ & new_n25499_;
  assign new_n25501_ = ~new_n24757_ & ~new_n25500_;
  assign new_n25502_ = \b[55]  & ~new_n24746_;
  assign new_n25503_ = ~new_n24744_ & new_n25502_;
  assign new_n25504_ = ~new_n24748_ & ~new_n25503_;
  assign new_n25505_ = ~new_n25501_ & new_n25504_;
  assign new_n25506_ = ~new_n24748_ & ~new_n25505_;
  assign new_n25507_ = \b[56]  & ~new_n24737_;
  assign new_n25508_ = ~new_n24735_ & new_n25507_;
  assign new_n25509_ = ~new_n24739_ & ~new_n25508_;
  assign new_n25510_ = ~new_n25506_ & new_n25509_;
  assign new_n25511_ = ~new_n24739_ & ~new_n25510_;
  assign new_n25512_ = \b[57]  & ~new_n24728_;
  assign new_n25513_ = ~new_n24726_ & new_n25512_;
  assign new_n25514_ = ~new_n24730_ & ~new_n25513_;
  assign new_n25515_ = ~new_n25511_ & new_n25514_;
  assign new_n25516_ = ~new_n24730_ & ~new_n25515_;
  assign new_n25517_ = \b[58]  & ~new_n24719_;
  assign new_n25518_ = ~new_n24717_ & new_n25517_;
  assign new_n25519_ = ~new_n24721_ & ~new_n25518_;
  assign new_n25520_ = ~new_n25516_ & new_n25519_;
  assign new_n25521_ = ~new_n24721_ & ~new_n25520_;
  assign new_n25522_ = ~new_n23905_ & ~new_n24706_;
  assign new_n25523_ = ~new_n24704_ & new_n25522_;
  assign new_n25524_ = ~new_n24695_ & new_n25523_;
  assign new_n25525_ = ~new_n24704_ & ~new_n24706_;
  assign new_n25526_ = ~new_n24696_ & ~new_n25525_;
  assign new_n25527_ = ~new_n25524_ & ~new_n25526_;
  assign new_n25528_ = \quotient[5]  & ~new_n25527_;
  assign new_n25529_ = ~new_n24703_ & ~new_n24711_;
  assign new_n25530_ = ~new_n24710_ & new_n25529_;
  assign new_n25531_ = ~new_n25528_ & ~new_n25530_;
  assign new_n25532_ = ~\b[59]  & ~new_n25531_;
  assign new_n25533_ = \b[59]  & ~new_n25530_;
  assign new_n25534_ = ~new_n25528_ & new_n25533_;
  assign new_n25535_ = new_n280_ & ~new_n25534_;
  assign new_n25536_ = ~new_n25532_ & new_n25535_;
  assign new_n25537_ = ~new_n25521_ & new_n25536_;
  assign new_n25538_ = new_n24707_ & ~new_n25531_;
  assign \quotient[4]  = new_n25537_ | new_n25538_;
  assign new_n25540_ = ~new_n24730_ & new_n25519_;
  assign new_n25541_ = ~new_n25515_ & new_n25540_;
  assign new_n25542_ = ~new_n25516_ & ~new_n25519_;
  assign new_n25543_ = ~new_n25541_ & ~new_n25542_;
  assign new_n25544_ = \quotient[4]  & ~new_n25543_;
  assign new_n25545_ = ~new_n24720_ & ~new_n25538_;
  assign new_n25546_ = ~new_n25537_ & new_n25545_;
  assign new_n25547_ = ~new_n25544_ & ~new_n25546_;
  assign new_n25548_ = ~\b[59]  & ~new_n25547_;
  assign new_n25549_ = ~new_n24739_ & new_n25514_;
  assign new_n25550_ = ~new_n25510_ & new_n25549_;
  assign new_n25551_ = ~new_n25511_ & ~new_n25514_;
  assign new_n25552_ = ~new_n25550_ & ~new_n25551_;
  assign new_n25553_ = \quotient[4]  & ~new_n25552_;
  assign new_n25554_ = ~new_n24729_ & ~new_n25538_;
  assign new_n25555_ = ~new_n25537_ & new_n25554_;
  assign new_n25556_ = ~new_n25553_ & ~new_n25555_;
  assign new_n25557_ = ~\b[58]  & ~new_n25556_;
  assign new_n25558_ = ~new_n24748_ & new_n25509_;
  assign new_n25559_ = ~new_n25505_ & new_n25558_;
  assign new_n25560_ = ~new_n25506_ & ~new_n25509_;
  assign new_n25561_ = ~new_n25559_ & ~new_n25560_;
  assign new_n25562_ = \quotient[4]  & ~new_n25561_;
  assign new_n25563_ = ~new_n24738_ & ~new_n25538_;
  assign new_n25564_ = ~new_n25537_ & new_n25563_;
  assign new_n25565_ = ~new_n25562_ & ~new_n25564_;
  assign new_n25566_ = ~\b[57]  & ~new_n25565_;
  assign new_n25567_ = ~new_n24757_ & new_n25504_;
  assign new_n25568_ = ~new_n25500_ & new_n25567_;
  assign new_n25569_ = ~new_n25501_ & ~new_n25504_;
  assign new_n25570_ = ~new_n25568_ & ~new_n25569_;
  assign new_n25571_ = \quotient[4]  & ~new_n25570_;
  assign new_n25572_ = ~new_n24747_ & ~new_n25538_;
  assign new_n25573_ = ~new_n25537_ & new_n25572_;
  assign new_n25574_ = ~new_n25571_ & ~new_n25573_;
  assign new_n25575_ = ~\b[56]  & ~new_n25574_;
  assign new_n25576_ = ~new_n24766_ & new_n25499_;
  assign new_n25577_ = ~new_n25495_ & new_n25576_;
  assign new_n25578_ = ~new_n25496_ & ~new_n25499_;
  assign new_n25579_ = ~new_n25577_ & ~new_n25578_;
  assign new_n25580_ = \quotient[4]  & ~new_n25579_;
  assign new_n25581_ = ~new_n24756_ & ~new_n25538_;
  assign new_n25582_ = ~new_n25537_ & new_n25581_;
  assign new_n25583_ = ~new_n25580_ & ~new_n25582_;
  assign new_n25584_ = ~\b[55]  & ~new_n25583_;
  assign new_n25585_ = ~new_n24775_ & new_n25494_;
  assign new_n25586_ = ~new_n25490_ & new_n25585_;
  assign new_n25587_ = ~new_n25491_ & ~new_n25494_;
  assign new_n25588_ = ~new_n25586_ & ~new_n25587_;
  assign new_n25589_ = \quotient[4]  & ~new_n25588_;
  assign new_n25590_ = ~new_n24765_ & ~new_n25538_;
  assign new_n25591_ = ~new_n25537_ & new_n25590_;
  assign new_n25592_ = ~new_n25589_ & ~new_n25591_;
  assign new_n25593_ = ~\b[54]  & ~new_n25592_;
  assign new_n25594_ = ~new_n24784_ & new_n25489_;
  assign new_n25595_ = ~new_n25485_ & new_n25594_;
  assign new_n25596_ = ~new_n25486_ & ~new_n25489_;
  assign new_n25597_ = ~new_n25595_ & ~new_n25596_;
  assign new_n25598_ = \quotient[4]  & ~new_n25597_;
  assign new_n25599_ = ~new_n24774_ & ~new_n25538_;
  assign new_n25600_ = ~new_n25537_ & new_n25599_;
  assign new_n25601_ = ~new_n25598_ & ~new_n25600_;
  assign new_n25602_ = ~\b[53]  & ~new_n25601_;
  assign new_n25603_ = ~new_n24793_ & new_n25484_;
  assign new_n25604_ = ~new_n25480_ & new_n25603_;
  assign new_n25605_ = ~new_n25481_ & ~new_n25484_;
  assign new_n25606_ = ~new_n25604_ & ~new_n25605_;
  assign new_n25607_ = \quotient[4]  & ~new_n25606_;
  assign new_n25608_ = ~new_n24783_ & ~new_n25538_;
  assign new_n25609_ = ~new_n25537_ & new_n25608_;
  assign new_n25610_ = ~new_n25607_ & ~new_n25609_;
  assign new_n25611_ = ~\b[52]  & ~new_n25610_;
  assign new_n25612_ = ~new_n24802_ & new_n25479_;
  assign new_n25613_ = ~new_n25475_ & new_n25612_;
  assign new_n25614_ = ~new_n25476_ & ~new_n25479_;
  assign new_n25615_ = ~new_n25613_ & ~new_n25614_;
  assign new_n25616_ = \quotient[4]  & ~new_n25615_;
  assign new_n25617_ = ~new_n24792_ & ~new_n25538_;
  assign new_n25618_ = ~new_n25537_ & new_n25617_;
  assign new_n25619_ = ~new_n25616_ & ~new_n25618_;
  assign new_n25620_ = ~\b[51]  & ~new_n25619_;
  assign new_n25621_ = ~new_n24811_ & new_n25474_;
  assign new_n25622_ = ~new_n25470_ & new_n25621_;
  assign new_n25623_ = ~new_n25471_ & ~new_n25474_;
  assign new_n25624_ = ~new_n25622_ & ~new_n25623_;
  assign new_n25625_ = \quotient[4]  & ~new_n25624_;
  assign new_n25626_ = ~new_n24801_ & ~new_n25538_;
  assign new_n25627_ = ~new_n25537_ & new_n25626_;
  assign new_n25628_ = ~new_n25625_ & ~new_n25627_;
  assign new_n25629_ = ~\b[50]  & ~new_n25628_;
  assign new_n25630_ = ~new_n24820_ & new_n25469_;
  assign new_n25631_ = ~new_n25465_ & new_n25630_;
  assign new_n25632_ = ~new_n25466_ & ~new_n25469_;
  assign new_n25633_ = ~new_n25631_ & ~new_n25632_;
  assign new_n25634_ = \quotient[4]  & ~new_n25633_;
  assign new_n25635_ = ~new_n24810_ & ~new_n25538_;
  assign new_n25636_ = ~new_n25537_ & new_n25635_;
  assign new_n25637_ = ~new_n25634_ & ~new_n25636_;
  assign new_n25638_ = ~\b[49]  & ~new_n25637_;
  assign new_n25639_ = ~new_n24829_ & new_n25464_;
  assign new_n25640_ = ~new_n25460_ & new_n25639_;
  assign new_n25641_ = ~new_n25461_ & ~new_n25464_;
  assign new_n25642_ = ~new_n25640_ & ~new_n25641_;
  assign new_n25643_ = \quotient[4]  & ~new_n25642_;
  assign new_n25644_ = ~new_n24819_ & ~new_n25538_;
  assign new_n25645_ = ~new_n25537_ & new_n25644_;
  assign new_n25646_ = ~new_n25643_ & ~new_n25645_;
  assign new_n25647_ = ~\b[48]  & ~new_n25646_;
  assign new_n25648_ = ~new_n24838_ & new_n25459_;
  assign new_n25649_ = ~new_n25455_ & new_n25648_;
  assign new_n25650_ = ~new_n25456_ & ~new_n25459_;
  assign new_n25651_ = ~new_n25649_ & ~new_n25650_;
  assign new_n25652_ = \quotient[4]  & ~new_n25651_;
  assign new_n25653_ = ~new_n24828_ & ~new_n25538_;
  assign new_n25654_ = ~new_n25537_ & new_n25653_;
  assign new_n25655_ = ~new_n25652_ & ~new_n25654_;
  assign new_n25656_ = ~\b[47]  & ~new_n25655_;
  assign new_n25657_ = ~new_n24847_ & new_n25454_;
  assign new_n25658_ = ~new_n25450_ & new_n25657_;
  assign new_n25659_ = ~new_n25451_ & ~new_n25454_;
  assign new_n25660_ = ~new_n25658_ & ~new_n25659_;
  assign new_n25661_ = \quotient[4]  & ~new_n25660_;
  assign new_n25662_ = ~new_n24837_ & ~new_n25538_;
  assign new_n25663_ = ~new_n25537_ & new_n25662_;
  assign new_n25664_ = ~new_n25661_ & ~new_n25663_;
  assign new_n25665_ = ~\b[46]  & ~new_n25664_;
  assign new_n25666_ = ~new_n24856_ & new_n25449_;
  assign new_n25667_ = ~new_n25445_ & new_n25666_;
  assign new_n25668_ = ~new_n25446_ & ~new_n25449_;
  assign new_n25669_ = ~new_n25667_ & ~new_n25668_;
  assign new_n25670_ = \quotient[4]  & ~new_n25669_;
  assign new_n25671_ = ~new_n24846_ & ~new_n25538_;
  assign new_n25672_ = ~new_n25537_ & new_n25671_;
  assign new_n25673_ = ~new_n25670_ & ~new_n25672_;
  assign new_n25674_ = ~\b[45]  & ~new_n25673_;
  assign new_n25675_ = ~new_n24865_ & new_n25444_;
  assign new_n25676_ = ~new_n25440_ & new_n25675_;
  assign new_n25677_ = ~new_n25441_ & ~new_n25444_;
  assign new_n25678_ = ~new_n25676_ & ~new_n25677_;
  assign new_n25679_ = \quotient[4]  & ~new_n25678_;
  assign new_n25680_ = ~new_n24855_ & ~new_n25538_;
  assign new_n25681_ = ~new_n25537_ & new_n25680_;
  assign new_n25682_ = ~new_n25679_ & ~new_n25681_;
  assign new_n25683_ = ~\b[44]  & ~new_n25682_;
  assign new_n25684_ = ~new_n24874_ & new_n25439_;
  assign new_n25685_ = ~new_n25435_ & new_n25684_;
  assign new_n25686_ = ~new_n25436_ & ~new_n25439_;
  assign new_n25687_ = ~new_n25685_ & ~new_n25686_;
  assign new_n25688_ = \quotient[4]  & ~new_n25687_;
  assign new_n25689_ = ~new_n24864_ & ~new_n25538_;
  assign new_n25690_ = ~new_n25537_ & new_n25689_;
  assign new_n25691_ = ~new_n25688_ & ~new_n25690_;
  assign new_n25692_ = ~\b[43]  & ~new_n25691_;
  assign new_n25693_ = ~new_n24883_ & new_n25434_;
  assign new_n25694_ = ~new_n25430_ & new_n25693_;
  assign new_n25695_ = ~new_n25431_ & ~new_n25434_;
  assign new_n25696_ = ~new_n25694_ & ~new_n25695_;
  assign new_n25697_ = \quotient[4]  & ~new_n25696_;
  assign new_n25698_ = ~new_n24873_ & ~new_n25538_;
  assign new_n25699_ = ~new_n25537_ & new_n25698_;
  assign new_n25700_ = ~new_n25697_ & ~new_n25699_;
  assign new_n25701_ = ~\b[42]  & ~new_n25700_;
  assign new_n25702_ = ~new_n24892_ & new_n25429_;
  assign new_n25703_ = ~new_n25425_ & new_n25702_;
  assign new_n25704_ = ~new_n25426_ & ~new_n25429_;
  assign new_n25705_ = ~new_n25703_ & ~new_n25704_;
  assign new_n25706_ = \quotient[4]  & ~new_n25705_;
  assign new_n25707_ = ~new_n24882_ & ~new_n25538_;
  assign new_n25708_ = ~new_n25537_ & new_n25707_;
  assign new_n25709_ = ~new_n25706_ & ~new_n25708_;
  assign new_n25710_ = ~\b[41]  & ~new_n25709_;
  assign new_n25711_ = ~new_n24901_ & new_n25424_;
  assign new_n25712_ = ~new_n25420_ & new_n25711_;
  assign new_n25713_ = ~new_n25421_ & ~new_n25424_;
  assign new_n25714_ = ~new_n25712_ & ~new_n25713_;
  assign new_n25715_ = \quotient[4]  & ~new_n25714_;
  assign new_n25716_ = ~new_n24891_ & ~new_n25538_;
  assign new_n25717_ = ~new_n25537_ & new_n25716_;
  assign new_n25718_ = ~new_n25715_ & ~new_n25717_;
  assign new_n25719_ = ~\b[40]  & ~new_n25718_;
  assign new_n25720_ = ~new_n24910_ & new_n25419_;
  assign new_n25721_ = ~new_n25415_ & new_n25720_;
  assign new_n25722_ = ~new_n25416_ & ~new_n25419_;
  assign new_n25723_ = ~new_n25721_ & ~new_n25722_;
  assign new_n25724_ = \quotient[4]  & ~new_n25723_;
  assign new_n25725_ = ~new_n24900_ & ~new_n25538_;
  assign new_n25726_ = ~new_n25537_ & new_n25725_;
  assign new_n25727_ = ~new_n25724_ & ~new_n25726_;
  assign new_n25728_ = ~\b[39]  & ~new_n25727_;
  assign new_n25729_ = ~new_n24919_ & new_n25414_;
  assign new_n25730_ = ~new_n25410_ & new_n25729_;
  assign new_n25731_ = ~new_n25411_ & ~new_n25414_;
  assign new_n25732_ = ~new_n25730_ & ~new_n25731_;
  assign new_n25733_ = \quotient[4]  & ~new_n25732_;
  assign new_n25734_ = ~new_n24909_ & ~new_n25538_;
  assign new_n25735_ = ~new_n25537_ & new_n25734_;
  assign new_n25736_ = ~new_n25733_ & ~new_n25735_;
  assign new_n25737_ = ~\b[38]  & ~new_n25736_;
  assign new_n25738_ = ~new_n24928_ & new_n25409_;
  assign new_n25739_ = ~new_n25405_ & new_n25738_;
  assign new_n25740_ = ~new_n25406_ & ~new_n25409_;
  assign new_n25741_ = ~new_n25739_ & ~new_n25740_;
  assign new_n25742_ = \quotient[4]  & ~new_n25741_;
  assign new_n25743_ = ~new_n24918_ & ~new_n25538_;
  assign new_n25744_ = ~new_n25537_ & new_n25743_;
  assign new_n25745_ = ~new_n25742_ & ~new_n25744_;
  assign new_n25746_ = ~\b[37]  & ~new_n25745_;
  assign new_n25747_ = ~new_n24937_ & new_n25404_;
  assign new_n25748_ = ~new_n25400_ & new_n25747_;
  assign new_n25749_ = ~new_n25401_ & ~new_n25404_;
  assign new_n25750_ = ~new_n25748_ & ~new_n25749_;
  assign new_n25751_ = \quotient[4]  & ~new_n25750_;
  assign new_n25752_ = ~new_n24927_ & ~new_n25538_;
  assign new_n25753_ = ~new_n25537_ & new_n25752_;
  assign new_n25754_ = ~new_n25751_ & ~new_n25753_;
  assign new_n25755_ = ~\b[36]  & ~new_n25754_;
  assign new_n25756_ = ~new_n24946_ & new_n25399_;
  assign new_n25757_ = ~new_n25395_ & new_n25756_;
  assign new_n25758_ = ~new_n25396_ & ~new_n25399_;
  assign new_n25759_ = ~new_n25757_ & ~new_n25758_;
  assign new_n25760_ = \quotient[4]  & ~new_n25759_;
  assign new_n25761_ = ~new_n24936_ & ~new_n25538_;
  assign new_n25762_ = ~new_n25537_ & new_n25761_;
  assign new_n25763_ = ~new_n25760_ & ~new_n25762_;
  assign new_n25764_ = ~\b[35]  & ~new_n25763_;
  assign new_n25765_ = ~new_n24955_ & new_n25394_;
  assign new_n25766_ = ~new_n25390_ & new_n25765_;
  assign new_n25767_ = ~new_n25391_ & ~new_n25394_;
  assign new_n25768_ = ~new_n25766_ & ~new_n25767_;
  assign new_n25769_ = \quotient[4]  & ~new_n25768_;
  assign new_n25770_ = ~new_n24945_ & ~new_n25538_;
  assign new_n25771_ = ~new_n25537_ & new_n25770_;
  assign new_n25772_ = ~new_n25769_ & ~new_n25771_;
  assign new_n25773_ = ~\b[34]  & ~new_n25772_;
  assign new_n25774_ = ~new_n24964_ & new_n25389_;
  assign new_n25775_ = ~new_n25385_ & new_n25774_;
  assign new_n25776_ = ~new_n25386_ & ~new_n25389_;
  assign new_n25777_ = ~new_n25775_ & ~new_n25776_;
  assign new_n25778_ = \quotient[4]  & ~new_n25777_;
  assign new_n25779_ = ~new_n24954_ & ~new_n25538_;
  assign new_n25780_ = ~new_n25537_ & new_n25779_;
  assign new_n25781_ = ~new_n25778_ & ~new_n25780_;
  assign new_n25782_ = ~\b[33]  & ~new_n25781_;
  assign new_n25783_ = ~new_n24973_ & new_n25384_;
  assign new_n25784_ = ~new_n25380_ & new_n25783_;
  assign new_n25785_ = ~new_n25381_ & ~new_n25384_;
  assign new_n25786_ = ~new_n25784_ & ~new_n25785_;
  assign new_n25787_ = \quotient[4]  & ~new_n25786_;
  assign new_n25788_ = ~new_n24963_ & ~new_n25538_;
  assign new_n25789_ = ~new_n25537_ & new_n25788_;
  assign new_n25790_ = ~new_n25787_ & ~new_n25789_;
  assign new_n25791_ = ~\b[32]  & ~new_n25790_;
  assign new_n25792_ = ~new_n24982_ & new_n25379_;
  assign new_n25793_ = ~new_n25375_ & new_n25792_;
  assign new_n25794_ = ~new_n25376_ & ~new_n25379_;
  assign new_n25795_ = ~new_n25793_ & ~new_n25794_;
  assign new_n25796_ = \quotient[4]  & ~new_n25795_;
  assign new_n25797_ = ~new_n24972_ & ~new_n25538_;
  assign new_n25798_ = ~new_n25537_ & new_n25797_;
  assign new_n25799_ = ~new_n25796_ & ~new_n25798_;
  assign new_n25800_ = ~\b[31]  & ~new_n25799_;
  assign new_n25801_ = ~new_n24991_ & new_n25374_;
  assign new_n25802_ = ~new_n25370_ & new_n25801_;
  assign new_n25803_ = ~new_n25371_ & ~new_n25374_;
  assign new_n25804_ = ~new_n25802_ & ~new_n25803_;
  assign new_n25805_ = \quotient[4]  & ~new_n25804_;
  assign new_n25806_ = ~new_n24981_ & ~new_n25538_;
  assign new_n25807_ = ~new_n25537_ & new_n25806_;
  assign new_n25808_ = ~new_n25805_ & ~new_n25807_;
  assign new_n25809_ = ~\b[30]  & ~new_n25808_;
  assign new_n25810_ = ~new_n25000_ & new_n25369_;
  assign new_n25811_ = ~new_n25365_ & new_n25810_;
  assign new_n25812_ = ~new_n25366_ & ~new_n25369_;
  assign new_n25813_ = ~new_n25811_ & ~new_n25812_;
  assign new_n25814_ = \quotient[4]  & ~new_n25813_;
  assign new_n25815_ = ~new_n24990_ & ~new_n25538_;
  assign new_n25816_ = ~new_n25537_ & new_n25815_;
  assign new_n25817_ = ~new_n25814_ & ~new_n25816_;
  assign new_n25818_ = ~\b[29]  & ~new_n25817_;
  assign new_n25819_ = ~new_n25009_ & new_n25364_;
  assign new_n25820_ = ~new_n25360_ & new_n25819_;
  assign new_n25821_ = ~new_n25361_ & ~new_n25364_;
  assign new_n25822_ = ~new_n25820_ & ~new_n25821_;
  assign new_n25823_ = \quotient[4]  & ~new_n25822_;
  assign new_n25824_ = ~new_n24999_ & ~new_n25538_;
  assign new_n25825_ = ~new_n25537_ & new_n25824_;
  assign new_n25826_ = ~new_n25823_ & ~new_n25825_;
  assign new_n25827_ = ~\b[28]  & ~new_n25826_;
  assign new_n25828_ = ~new_n25018_ & new_n25359_;
  assign new_n25829_ = ~new_n25355_ & new_n25828_;
  assign new_n25830_ = ~new_n25356_ & ~new_n25359_;
  assign new_n25831_ = ~new_n25829_ & ~new_n25830_;
  assign new_n25832_ = \quotient[4]  & ~new_n25831_;
  assign new_n25833_ = ~new_n25008_ & ~new_n25538_;
  assign new_n25834_ = ~new_n25537_ & new_n25833_;
  assign new_n25835_ = ~new_n25832_ & ~new_n25834_;
  assign new_n25836_ = ~\b[27]  & ~new_n25835_;
  assign new_n25837_ = ~new_n25027_ & new_n25354_;
  assign new_n25838_ = ~new_n25350_ & new_n25837_;
  assign new_n25839_ = ~new_n25351_ & ~new_n25354_;
  assign new_n25840_ = ~new_n25838_ & ~new_n25839_;
  assign new_n25841_ = \quotient[4]  & ~new_n25840_;
  assign new_n25842_ = ~new_n25017_ & ~new_n25538_;
  assign new_n25843_ = ~new_n25537_ & new_n25842_;
  assign new_n25844_ = ~new_n25841_ & ~new_n25843_;
  assign new_n25845_ = ~\b[26]  & ~new_n25844_;
  assign new_n25846_ = ~new_n25036_ & new_n25349_;
  assign new_n25847_ = ~new_n25345_ & new_n25846_;
  assign new_n25848_ = ~new_n25346_ & ~new_n25349_;
  assign new_n25849_ = ~new_n25847_ & ~new_n25848_;
  assign new_n25850_ = \quotient[4]  & ~new_n25849_;
  assign new_n25851_ = ~new_n25026_ & ~new_n25538_;
  assign new_n25852_ = ~new_n25537_ & new_n25851_;
  assign new_n25853_ = ~new_n25850_ & ~new_n25852_;
  assign new_n25854_ = ~\b[25]  & ~new_n25853_;
  assign new_n25855_ = ~new_n25045_ & new_n25344_;
  assign new_n25856_ = ~new_n25340_ & new_n25855_;
  assign new_n25857_ = ~new_n25341_ & ~new_n25344_;
  assign new_n25858_ = ~new_n25856_ & ~new_n25857_;
  assign new_n25859_ = \quotient[4]  & ~new_n25858_;
  assign new_n25860_ = ~new_n25035_ & ~new_n25538_;
  assign new_n25861_ = ~new_n25537_ & new_n25860_;
  assign new_n25862_ = ~new_n25859_ & ~new_n25861_;
  assign new_n25863_ = ~\b[24]  & ~new_n25862_;
  assign new_n25864_ = ~new_n25054_ & new_n25339_;
  assign new_n25865_ = ~new_n25335_ & new_n25864_;
  assign new_n25866_ = ~new_n25336_ & ~new_n25339_;
  assign new_n25867_ = ~new_n25865_ & ~new_n25866_;
  assign new_n25868_ = \quotient[4]  & ~new_n25867_;
  assign new_n25869_ = ~new_n25044_ & ~new_n25538_;
  assign new_n25870_ = ~new_n25537_ & new_n25869_;
  assign new_n25871_ = ~new_n25868_ & ~new_n25870_;
  assign new_n25872_ = ~\b[23]  & ~new_n25871_;
  assign new_n25873_ = ~new_n25063_ & new_n25334_;
  assign new_n25874_ = ~new_n25330_ & new_n25873_;
  assign new_n25875_ = ~new_n25331_ & ~new_n25334_;
  assign new_n25876_ = ~new_n25874_ & ~new_n25875_;
  assign new_n25877_ = \quotient[4]  & ~new_n25876_;
  assign new_n25878_ = ~new_n25053_ & ~new_n25538_;
  assign new_n25879_ = ~new_n25537_ & new_n25878_;
  assign new_n25880_ = ~new_n25877_ & ~new_n25879_;
  assign new_n25881_ = ~\b[22]  & ~new_n25880_;
  assign new_n25882_ = ~new_n25072_ & new_n25329_;
  assign new_n25883_ = ~new_n25325_ & new_n25882_;
  assign new_n25884_ = ~new_n25326_ & ~new_n25329_;
  assign new_n25885_ = ~new_n25883_ & ~new_n25884_;
  assign new_n25886_ = \quotient[4]  & ~new_n25885_;
  assign new_n25887_ = ~new_n25062_ & ~new_n25538_;
  assign new_n25888_ = ~new_n25537_ & new_n25887_;
  assign new_n25889_ = ~new_n25886_ & ~new_n25888_;
  assign new_n25890_ = ~\b[21]  & ~new_n25889_;
  assign new_n25891_ = ~new_n25081_ & new_n25324_;
  assign new_n25892_ = ~new_n25320_ & new_n25891_;
  assign new_n25893_ = ~new_n25321_ & ~new_n25324_;
  assign new_n25894_ = ~new_n25892_ & ~new_n25893_;
  assign new_n25895_ = \quotient[4]  & ~new_n25894_;
  assign new_n25896_ = ~new_n25071_ & ~new_n25538_;
  assign new_n25897_ = ~new_n25537_ & new_n25896_;
  assign new_n25898_ = ~new_n25895_ & ~new_n25897_;
  assign new_n25899_ = ~\b[20]  & ~new_n25898_;
  assign new_n25900_ = ~new_n25090_ & new_n25319_;
  assign new_n25901_ = ~new_n25315_ & new_n25900_;
  assign new_n25902_ = ~new_n25316_ & ~new_n25319_;
  assign new_n25903_ = ~new_n25901_ & ~new_n25902_;
  assign new_n25904_ = \quotient[4]  & ~new_n25903_;
  assign new_n25905_ = ~new_n25080_ & ~new_n25538_;
  assign new_n25906_ = ~new_n25537_ & new_n25905_;
  assign new_n25907_ = ~new_n25904_ & ~new_n25906_;
  assign new_n25908_ = ~\b[19]  & ~new_n25907_;
  assign new_n25909_ = ~new_n25099_ & new_n25314_;
  assign new_n25910_ = ~new_n25310_ & new_n25909_;
  assign new_n25911_ = ~new_n25311_ & ~new_n25314_;
  assign new_n25912_ = ~new_n25910_ & ~new_n25911_;
  assign new_n25913_ = \quotient[4]  & ~new_n25912_;
  assign new_n25914_ = ~new_n25089_ & ~new_n25538_;
  assign new_n25915_ = ~new_n25537_ & new_n25914_;
  assign new_n25916_ = ~new_n25913_ & ~new_n25915_;
  assign new_n25917_ = ~\b[18]  & ~new_n25916_;
  assign new_n25918_ = ~new_n25108_ & new_n25309_;
  assign new_n25919_ = ~new_n25305_ & new_n25918_;
  assign new_n25920_ = ~new_n25306_ & ~new_n25309_;
  assign new_n25921_ = ~new_n25919_ & ~new_n25920_;
  assign new_n25922_ = \quotient[4]  & ~new_n25921_;
  assign new_n25923_ = ~new_n25098_ & ~new_n25538_;
  assign new_n25924_ = ~new_n25537_ & new_n25923_;
  assign new_n25925_ = ~new_n25922_ & ~new_n25924_;
  assign new_n25926_ = ~\b[17]  & ~new_n25925_;
  assign new_n25927_ = ~new_n25117_ & new_n25304_;
  assign new_n25928_ = ~new_n25300_ & new_n25927_;
  assign new_n25929_ = ~new_n25301_ & ~new_n25304_;
  assign new_n25930_ = ~new_n25928_ & ~new_n25929_;
  assign new_n25931_ = \quotient[4]  & ~new_n25930_;
  assign new_n25932_ = ~new_n25107_ & ~new_n25538_;
  assign new_n25933_ = ~new_n25537_ & new_n25932_;
  assign new_n25934_ = ~new_n25931_ & ~new_n25933_;
  assign new_n25935_ = ~\b[16]  & ~new_n25934_;
  assign new_n25936_ = ~new_n25126_ & new_n25299_;
  assign new_n25937_ = ~new_n25295_ & new_n25936_;
  assign new_n25938_ = ~new_n25296_ & ~new_n25299_;
  assign new_n25939_ = ~new_n25937_ & ~new_n25938_;
  assign new_n25940_ = \quotient[4]  & ~new_n25939_;
  assign new_n25941_ = ~new_n25116_ & ~new_n25538_;
  assign new_n25942_ = ~new_n25537_ & new_n25941_;
  assign new_n25943_ = ~new_n25940_ & ~new_n25942_;
  assign new_n25944_ = ~\b[15]  & ~new_n25943_;
  assign new_n25945_ = ~new_n25135_ & new_n25294_;
  assign new_n25946_ = ~new_n25290_ & new_n25945_;
  assign new_n25947_ = ~new_n25291_ & ~new_n25294_;
  assign new_n25948_ = ~new_n25946_ & ~new_n25947_;
  assign new_n25949_ = \quotient[4]  & ~new_n25948_;
  assign new_n25950_ = ~new_n25125_ & ~new_n25538_;
  assign new_n25951_ = ~new_n25537_ & new_n25950_;
  assign new_n25952_ = ~new_n25949_ & ~new_n25951_;
  assign new_n25953_ = ~\b[14]  & ~new_n25952_;
  assign new_n25954_ = ~new_n25144_ & new_n25289_;
  assign new_n25955_ = ~new_n25285_ & new_n25954_;
  assign new_n25956_ = ~new_n25286_ & ~new_n25289_;
  assign new_n25957_ = ~new_n25955_ & ~new_n25956_;
  assign new_n25958_ = \quotient[4]  & ~new_n25957_;
  assign new_n25959_ = ~new_n25134_ & ~new_n25538_;
  assign new_n25960_ = ~new_n25537_ & new_n25959_;
  assign new_n25961_ = ~new_n25958_ & ~new_n25960_;
  assign new_n25962_ = ~\b[13]  & ~new_n25961_;
  assign new_n25963_ = ~new_n25153_ & new_n25284_;
  assign new_n25964_ = ~new_n25280_ & new_n25963_;
  assign new_n25965_ = ~new_n25281_ & ~new_n25284_;
  assign new_n25966_ = ~new_n25964_ & ~new_n25965_;
  assign new_n25967_ = \quotient[4]  & ~new_n25966_;
  assign new_n25968_ = ~new_n25143_ & ~new_n25538_;
  assign new_n25969_ = ~new_n25537_ & new_n25968_;
  assign new_n25970_ = ~new_n25967_ & ~new_n25969_;
  assign new_n25971_ = ~\b[12]  & ~new_n25970_;
  assign new_n25972_ = ~new_n25162_ & new_n25279_;
  assign new_n25973_ = ~new_n25275_ & new_n25972_;
  assign new_n25974_ = ~new_n25276_ & ~new_n25279_;
  assign new_n25975_ = ~new_n25973_ & ~new_n25974_;
  assign new_n25976_ = \quotient[4]  & ~new_n25975_;
  assign new_n25977_ = ~new_n25152_ & ~new_n25538_;
  assign new_n25978_ = ~new_n25537_ & new_n25977_;
  assign new_n25979_ = ~new_n25976_ & ~new_n25978_;
  assign new_n25980_ = ~\b[11]  & ~new_n25979_;
  assign new_n25981_ = ~new_n25171_ & new_n25274_;
  assign new_n25982_ = ~new_n25270_ & new_n25981_;
  assign new_n25983_ = ~new_n25271_ & ~new_n25274_;
  assign new_n25984_ = ~new_n25982_ & ~new_n25983_;
  assign new_n25985_ = \quotient[4]  & ~new_n25984_;
  assign new_n25986_ = ~new_n25161_ & ~new_n25538_;
  assign new_n25987_ = ~new_n25537_ & new_n25986_;
  assign new_n25988_ = ~new_n25985_ & ~new_n25987_;
  assign new_n25989_ = ~\b[10]  & ~new_n25988_;
  assign new_n25990_ = ~new_n25180_ & new_n25269_;
  assign new_n25991_ = ~new_n25265_ & new_n25990_;
  assign new_n25992_ = ~new_n25266_ & ~new_n25269_;
  assign new_n25993_ = ~new_n25991_ & ~new_n25992_;
  assign new_n25994_ = \quotient[4]  & ~new_n25993_;
  assign new_n25995_ = ~new_n25170_ & ~new_n25538_;
  assign new_n25996_ = ~new_n25537_ & new_n25995_;
  assign new_n25997_ = ~new_n25994_ & ~new_n25996_;
  assign new_n25998_ = ~\b[9]  & ~new_n25997_;
  assign new_n25999_ = ~new_n25189_ & new_n25264_;
  assign new_n26000_ = ~new_n25260_ & new_n25999_;
  assign new_n26001_ = ~new_n25261_ & ~new_n25264_;
  assign new_n26002_ = ~new_n26000_ & ~new_n26001_;
  assign new_n26003_ = \quotient[4]  & ~new_n26002_;
  assign new_n26004_ = ~new_n25179_ & ~new_n25538_;
  assign new_n26005_ = ~new_n25537_ & new_n26004_;
  assign new_n26006_ = ~new_n26003_ & ~new_n26005_;
  assign new_n26007_ = ~\b[8]  & ~new_n26006_;
  assign new_n26008_ = ~new_n25198_ & new_n25259_;
  assign new_n26009_ = ~new_n25255_ & new_n26008_;
  assign new_n26010_ = ~new_n25256_ & ~new_n25259_;
  assign new_n26011_ = ~new_n26009_ & ~new_n26010_;
  assign new_n26012_ = \quotient[4]  & ~new_n26011_;
  assign new_n26013_ = ~new_n25188_ & ~new_n25538_;
  assign new_n26014_ = ~new_n25537_ & new_n26013_;
  assign new_n26015_ = ~new_n26012_ & ~new_n26014_;
  assign new_n26016_ = ~\b[7]  & ~new_n26015_;
  assign new_n26017_ = ~new_n25207_ & new_n25254_;
  assign new_n26018_ = ~new_n25250_ & new_n26017_;
  assign new_n26019_ = ~new_n25251_ & ~new_n25254_;
  assign new_n26020_ = ~new_n26018_ & ~new_n26019_;
  assign new_n26021_ = \quotient[4]  & ~new_n26020_;
  assign new_n26022_ = ~new_n25197_ & ~new_n25538_;
  assign new_n26023_ = ~new_n25537_ & new_n26022_;
  assign new_n26024_ = ~new_n26021_ & ~new_n26023_;
  assign new_n26025_ = ~\b[6]  & ~new_n26024_;
  assign new_n26026_ = ~new_n25216_ & new_n25249_;
  assign new_n26027_ = ~new_n25245_ & new_n26026_;
  assign new_n26028_ = ~new_n25246_ & ~new_n25249_;
  assign new_n26029_ = ~new_n26027_ & ~new_n26028_;
  assign new_n26030_ = \quotient[4]  & ~new_n26029_;
  assign new_n26031_ = ~new_n25206_ & ~new_n25538_;
  assign new_n26032_ = ~new_n25537_ & new_n26031_;
  assign new_n26033_ = ~new_n26030_ & ~new_n26032_;
  assign new_n26034_ = ~\b[5]  & ~new_n26033_;
  assign new_n26035_ = ~new_n25224_ & new_n25244_;
  assign new_n26036_ = ~new_n25240_ & new_n26035_;
  assign new_n26037_ = ~new_n25241_ & ~new_n25244_;
  assign new_n26038_ = ~new_n26036_ & ~new_n26037_;
  assign new_n26039_ = \quotient[4]  & ~new_n26038_;
  assign new_n26040_ = ~new_n25215_ & ~new_n25538_;
  assign new_n26041_ = ~new_n25537_ & new_n26040_;
  assign new_n26042_ = ~new_n26039_ & ~new_n26041_;
  assign new_n26043_ = ~\b[4]  & ~new_n26042_;
  assign new_n26044_ = ~new_n25235_ & new_n25239_;
  assign new_n26045_ = ~new_n25234_ & new_n26044_;
  assign new_n26046_ = ~new_n25236_ & ~new_n25239_;
  assign new_n26047_ = ~new_n26045_ & ~new_n26046_;
  assign new_n26048_ = \quotient[4]  & ~new_n26047_;
  assign new_n26049_ = ~new_n25223_ & ~new_n25538_;
  assign new_n26050_ = ~new_n25537_ & new_n26049_;
  assign new_n26051_ = ~new_n26048_ & ~new_n26050_;
  assign new_n26052_ = ~\b[3]  & ~new_n26051_;
  assign new_n26053_ = ~new_n25231_ & new_n25233_;
  assign new_n26054_ = ~new_n25229_ & new_n26053_;
  assign new_n26055_ = ~new_n25234_ & ~new_n26054_;
  assign new_n26056_ = \quotient[4]  & new_n26055_;
  assign new_n26057_ = ~new_n25228_ & ~new_n25538_;
  assign new_n26058_ = ~new_n25537_ & new_n26057_;
  assign new_n26059_ = ~new_n26056_ & ~new_n26058_;
  assign new_n26060_ = ~\b[2]  & ~new_n26059_;
  assign new_n26061_ = \b[0]  & \quotient[4] ;
  assign new_n26062_ = \a[4]  & ~new_n26061_;
  assign new_n26063_ = new_n25233_ & \quotient[4] ;
  assign new_n26064_ = ~new_n26062_ & ~new_n26063_;
  assign new_n26065_ = \b[1]  & ~new_n26064_;
  assign new_n26066_ = ~\b[1]  & ~new_n26063_;
  assign new_n26067_ = ~new_n26062_ & new_n26066_;
  assign new_n26068_ = ~new_n26065_ & ~new_n26067_;
  assign new_n26069_ = ~\a[3]  & \b[0] ;
  assign new_n26070_ = ~new_n26068_ & ~new_n26069_;
  assign new_n26071_ = ~\b[1]  & ~new_n26064_;
  assign new_n26072_ = ~new_n26070_ & ~new_n26071_;
  assign new_n26073_ = \b[2]  & ~new_n26058_;
  assign new_n26074_ = ~new_n26056_ & new_n26073_;
  assign new_n26075_ = ~new_n26060_ & ~new_n26074_;
  assign new_n26076_ = ~new_n26072_ & new_n26075_;
  assign new_n26077_ = ~new_n26060_ & ~new_n26076_;
  assign new_n26078_ = \b[3]  & ~new_n26050_;
  assign new_n26079_ = ~new_n26048_ & new_n26078_;
  assign new_n26080_ = ~new_n26052_ & ~new_n26079_;
  assign new_n26081_ = ~new_n26077_ & new_n26080_;
  assign new_n26082_ = ~new_n26052_ & ~new_n26081_;
  assign new_n26083_ = \b[4]  & ~new_n26041_;
  assign new_n26084_ = ~new_n26039_ & new_n26083_;
  assign new_n26085_ = ~new_n26043_ & ~new_n26084_;
  assign new_n26086_ = ~new_n26082_ & new_n26085_;
  assign new_n26087_ = ~new_n26043_ & ~new_n26086_;
  assign new_n26088_ = \b[5]  & ~new_n26032_;
  assign new_n26089_ = ~new_n26030_ & new_n26088_;
  assign new_n26090_ = ~new_n26034_ & ~new_n26089_;
  assign new_n26091_ = ~new_n26087_ & new_n26090_;
  assign new_n26092_ = ~new_n26034_ & ~new_n26091_;
  assign new_n26093_ = \b[6]  & ~new_n26023_;
  assign new_n26094_ = ~new_n26021_ & new_n26093_;
  assign new_n26095_ = ~new_n26025_ & ~new_n26094_;
  assign new_n26096_ = ~new_n26092_ & new_n26095_;
  assign new_n26097_ = ~new_n26025_ & ~new_n26096_;
  assign new_n26098_ = \b[7]  & ~new_n26014_;
  assign new_n26099_ = ~new_n26012_ & new_n26098_;
  assign new_n26100_ = ~new_n26016_ & ~new_n26099_;
  assign new_n26101_ = ~new_n26097_ & new_n26100_;
  assign new_n26102_ = ~new_n26016_ & ~new_n26101_;
  assign new_n26103_ = \b[8]  & ~new_n26005_;
  assign new_n26104_ = ~new_n26003_ & new_n26103_;
  assign new_n26105_ = ~new_n26007_ & ~new_n26104_;
  assign new_n26106_ = ~new_n26102_ & new_n26105_;
  assign new_n26107_ = ~new_n26007_ & ~new_n26106_;
  assign new_n26108_ = \b[9]  & ~new_n25996_;
  assign new_n26109_ = ~new_n25994_ & new_n26108_;
  assign new_n26110_ = ~new_n25998_ & ~new_n26109_;
  assign new_n26111_ = ~new_n26107_ & new_n26110_;
  assign new_n26112_ = ~new_n25998_ & ~new_n26111_;
  assign new_n26113_ = \b[10]  & ~new_n25987_;
  assign new_n26114_ = ~new_n25985_ & new_n26113_;
  assign new_n26115_ = ~new_n25989_ & ~new_n26114_;
  assign new_n26116_ = ~new_n26112_ & new_n26115_;
  assign new_n26117_ = ~new_n25989_ & ~new_n26116_;
  assign new_n26118_ = \b[11]  & ~new_n25978_;
  assign new_n26119_ = ~new_n25976_ & new_n26118_;
  assign new_n26120_ = ~new_n25980_ & ~new_n26119_;
  assign new_n26121_ = ~new_n26117_ & new_n26120_;
  assign new_n26122_ = ~new_n25980_ & ~new_n26121_;
  assign new_n26123_ = \b[12]  & ~new_n25969_;
  assign new_n26124_ = ~new_n25967_ & new_n26123_;
  assign new_n26125_ = ~new_n25971_ & ~new_n26124_;
  assign new_n26126_ = ~new_n26122_ & new_n26125_;
  assign new_n26127_ = ~new_n25971_ & ~new_n26126_;
  assign new_n26128_ = \b[13]  & ~new_n25960_;
  assign new_n26129_ = ~new_n25958_ & new_n26128_;
  assign new_n26130_ = ~new_n25962_ & ~new_n26129_;
  assign new_n26131_ = ~new_n26127_ & new_n26130_;
  assign new_n26132_ = ~new_n25962_ & ~new_n26131_;
  assign new_n26133_ = \b[14]  & ~new_n25951_;
  assign new_n26134_ = ~new_n25949_ & new_n26133_;
  assign new_n26135_ = ~new_n25953_ & ~new_n26134_;
  assign new_n26136_ = ~new_n26132_ & new_n26135_;
  assign new_n26137_ = ~new_n25953_ & ~new_n26136_;
  assign new_n26138_ = \b[15]  & ~new_n25942_;
  assign new_n26139_ = ~new_n25940_ & new_n26138_;
  assign new_n26140_ = ~new_n25944_ & ~new_n26139_;
  assign new_n26141_ = ~new_n26137_ & new_n26140_;
  assign new_n26142_ = ~new_n25944_ & ~new_n26141_;
  assign new_n26143_ = \b[16]  & ~new_n25933_;
  assign new_n26144_ = ~new_n25931_ & new_n26143_;
  assign new_n26145_ = ~new_n25935_ & ~new_n26144_;
  assign new_n26146_ = ~new_n26142_ & new_n26145_;
  assign new_n26147_ = ~new_n25935_ & ~new_n26146_;
  assign new_n26148_ = \b[17]  & ~new_n25924_;
  assign new_n26149_ = ~new_n25922_ & new_n26148_;
  assign new_n26150_ = ~new_n25926_ & ~new_n26149_;
  assign new_n26151_ = ~new_n26147_ & new_n26150_;
  assign new_n26152_ = ~new_n25926_ & ~new_n26151_;
  assign new_n26153_ = \b[18]  & ~new_n25915_;
  assign new_n26154_ = ~new_n25913_ & new_n26153_;
  assign new_n26155_ = ~new_n25917_ & ~new_n26154_;
  assign new_n26156_ = ~new_n26152_ & new_n26155_;
  assign new_n26157_ = ~new_n25917_ & ~new_n26156_;
  assign new_n26158_ = \b[19]  & ~new_n25906_;
  assign new_n26159_ = ~new_n25904_ & new_n26158_;
  assign new_n26160_ = ~new_n25908_ & ~new_n26159_;
  assign new_n26161_ = ~new_n26157_ & new_n26160_;
  assign new_n26162_ = ~new_n25908_ & ~new_n26161_;
  assign new_n26163_ = \b[20]  & ~new_n25897_;
  assign new_n26164_ = ~new_n25895_ & new_n26163_;
  assign new_n26165_ = ~new_n25899_ & ~new_n26164_;
  assign new_n26166_ = ~new_n26162_ & new_n26165_;
  assign new_n26167_ = ~new_n25899_ & ~new_n26166_;
  assign new_n26168_ = \b[21]  & ~new_n25888_;
  assign new_n26169_ = ~new_n25886_ & new_n26168_;
  assign new_n26170_ = ~new_n25890_ & ~new_n26169_;
  assign new_n26171_ = ~new_n26167_ & new_n26170_;
  assign new_n26172_ = ~new_n25890_ & ~new_n26171_;
  assign new_n26173_ = \b[22]  & ~new_n25879_;
  assign new_n26174_ = ~new_n25877_ & new_n26173_;
  assign new_n26175_ = ~new_n25881_ & ~new_n26174_;
  assign new_n26176_ = ~new_n26172_ & new_n26175_;
  assign new_n26177_ = ~new_n25881_ & ~new_n26176_;
  assign new_n26178_ = \b[23]  & ~new_n25870_;
  assign new_n26179_ = ~new_n25868_ & new_n26178_;
  assign new_n26180_ = ~new_n25872_ & ~new_n26179_;
  assign new_n26181_ = ~new_n26177_ & new_n26180_;
  assign new_n26182_ = ~new_n25872_ & ~new_n26181_;
  assign new_n26183_ = \b[24]  & ~new_n25861_;
  assign new_n26184_ = ~new_n25859_ & new_n26183_;
  assign new_n26185_ = ~new_n25863_ & ~new_n26184_;
  assign new_n26186_ = ~new_n26182_ & new_n26185_;
  assign new_n26187_ = ~new_n25863_ & ~new_n26186_;
  assign new_n26188_ = \b[25]  & ~new_n25852_;
  assign new_n26189_ = ~new_n25850_ & new_n26188_;
  assign new_n26190_ = ~new_n25854_ & ~new_n26189_;
  assign new_n26191_ = ~new_n26187_ & new_n26190_;
  assign new_n26192_ = ~new_n25854_ & ~new_n26191_;
  assign new_n26193_ = \b[26]  & ~new_n25843_;
  assign new_n26194_ = ~new_n25841_ & new_n26193_;
  assign new_n26195_ = ~new_n25845_ & ~new_n26194_;
  assign new_n26196_ = ~new_n26192_ & new_n26195_;
  assign new_n26197_ = ~new_n25845_ & ~new_n26196_;
  assign new_n26198_ = \b[27]  & ~new_n25834_;
  assign new_n26199_ = ~new_n25832_ & new_n26198_;
  assign new_n26200_ = ~new_n25836_ & ~new_n26199_;
  assign new_n26201_ = ~new_n26197_ & new_n26200_;
  assign new_n26202_ = ~new_n25836_ & ~new_n26201_;
  assign new_n26203_ = \b[28]  & ~new_n25825_;
  assign new_n26204_ = ~new_n25823_ & new_n26203_;
  assign new_n26205_ = ~new_n25827_ & ~new_n26204_;
  assign new_n26206_ = ~new_n26202_ & new_n26205_;
  assign new_n26207_ = ~new_n25827_ & ~new_n26206_;
  assign new_n26208_ = \b[29]  & ~new_n25816_;
  assign new_n26209_ = ~new_n25814_ & new_n26208_;
  assign new_n26210_ = ~new_n25818_ & ~new_n26209_;
  assign new_n26211_ = ~new_n26207_ & new_n26210_;
  assign new_n26212_ = ~new_n25818_ & ~new_n26211_;
  assign new_n26213_ = \b[30]  & ~new_n25807_;
  assign new_n26214_ = ~new_n25805_ & new_n26213_;
  assign new_n26215_ = ~new_n25809_ & ~new_n26214_;
  assign new_n26216_ = ~new_n26212_ & new_n26215_;
  assign new_n26217_ = ~new_n25809_ & ~new_n26216_;
  assign new_n26218_ = \b[31]  & ~new_n25798_;
  assign new_n26219_ = ~new_n25796_ & new_n26218_;
  assign new_n26220_ = ~new_n25800_ & ~new_n26219_;
  assign new_n26221_ = ~new_n26217_ & new_n26220_;
  assign new_n26222_ = ~new_n25800_ & ~new_n26221_;
  assign new_n26223_ = \b[32]  & ~new_n25789_;
  assign new_n26224_ = ~new_n25787_ & new_n26223_;
  assign new_n26225_ = ~new_n25791_ & ~new_n26224_;
  assign new_n26226_ = ~new_n26222_ & new_n26225_;
  assign new_n26227_ = ~new_n25791_ & ~new_n26226_;
  assign new_n26228_ = \b[33]  & ~new_n25780_;
  assign new_n26229_ = ~new_n25778_ & new_n26228_;
  assign new_n26230_ = ~new_n25782_ & ~new_n26229_;
  assign new_n26231_ = ~new_n26227_ & new_n26230_;
  assign new_n26232_ = ~new_n25782_ & ~new_n26231_;
  assign new_n26233_ = \b[34]  & ~new_n25771_;
  assign new_n26234_ = ~new_n25769_ & new_n26233_;
  assign new_n26235_ = ~new_n25773_ & ~new_n26234_;
  assign new_n26236_ = ~new_n26232_ & new_n26235_;
  assign new_n26237_ = ~new_n25773_ & ~new_n26236_;
  assign new_n26238_ = \b[35]  & ~new_n25762_;
  assign new_n26239_ = ~new_n25760_ & new_n26238_;
  assign new_n26240_ = ~new_n25764_ & ~new_n26239_;
  assign new_n26241_ = ~new_n26237_ & new_n26240_;
  assign new_n26242_ = ~new_n25764_ & ~new_n26241_;
  assign new_n26243_ = \b[36]  & ~new_n25753_;
  assign new_n26244_ = ~new_n25751_ & new_n26243_;
  assign new_n26245_ = ~new_n25755_ & ~new_n26244_;
  assign new_n26246_ = ~new_n26242_ & new_n26245_;
  assign new_n26247_ = ~new_n25755_ & ~new_n26246_;
  assign new_n26248_ = \b[37]  & ~new_n25744_;
  assign new_n26249_ = ~new_n25742_ & new_n26248_;
  assign new_n26250_ = ~new_n25746_ & ~new_n26249_;
  assign new_n26251_ = ~new_n26247_ & new_n26250_;
  assign new_n26252_ = ~new_n25746_ & ~new_n26251_;
  assign new_n26253_ = \b[38]  & ~new_n25735_;
  assign new_n26254_ = ~new_n25733_ & new_n26253_;
  assign new_n26255_ = ~new_n25737_ & ~new_n26254_;
  assign new_n26256_ = ~new_n26252_ & new_n26255_;
  assign new_n26257_ = ~new_n25737_ & ~new_n26256_;
  assign new_n26258_ = \b[39]  & ~new_n25726_;
  assign new_n26259_ = ~new_n25724_ & new_n26258_;
  assign new_n26260_ = ~new_n25728_ & ~new_n26259_;
  assign new_n26261_ = ~new_n26257_ & new_n26260_;
  assign new_n26262_ = ~new_n25728_ & ~new_n26261_;
  assign new_n26263_ = \b[40]  & ~new_n25717_;
  assign new_n26264_ = ~new_n25715_ & new_n26263_;
  assign new_n26265_ = ~new_n25719_ & ~new_n26264_;
  assign new_n26266_ = ~new_n26262_ & new_n26265_;
  assign new_n26267_ = ~new_n25719_ & ~new_n26266_;
  assign new_n26268_ = \b[41]  & ~new_n25708_;
  assign new_n26269_ = ~new_n25706_ & new_n26268_;
  assign new_n26270_ = ~new_n25710_ & ~new_n26269_;
  assign new_n26271_ = ~new_n26267_ & new_n26270_;
  assign new_n26272_ = ~new_n25710_ & ~new_n26271_;
  assign new_n26273_ = \b[42]  & ~new_n25699_;
  assign new_n26274_ = ~new_n25697_ & new_n26273_;
  assign new_n26275_ = ~new_n25701_ & ~new_n26274_;
  assign new_n26276_ = ~new_n26272_ & new_n26275_;
  assign new_n26277_ = ~new_n25701_ & ~new_n26276_;
  assign new_n26278_ = \b[43]  & ~new_n25690_;
  assign new_n26279_ = ~new_n25688_ & new_n26278_;
  assign new_n26280_ = ~new_n25692_ & ~new_n26279_;
  assign new_n26281_ = ~new_n26277_ & new_n26280_;
  assign new_n26282_ = ~new_n25692_ & ~new_n26281_;
  assign new_n26283_ = \b[44]  & ~new_n25681_;
  assign new_n26284_ = ~new_n25679_ & new_n26283_;
  assign new_n26285_ = ~new_n25683_ & ~new_n26284_;
  assign new_n26286_ = ~new_n26282_ & new_n26285_;
  assign new_n26287_ = ~new_n25683_ & ~new_n26286_;
  assign new_n26288_ = \b[45]  & ~new_n25672_;
  assign new_n26289_ = ~new_n25670_ & new_n26288_;
  assign new_n26290_ = ~new_n25674_ & ~new_n26289_;
  assign new_n26291_ = ~new_n26287_ & new_n26290_;
  assign new_n26292_ = ~new_n25674_ & ~new_n26291_;
  assign new_n26293_ = \b[46]  & ~new_n25663_;
  assign new_n26294_ = ~new_n25661_ & new_n26293_;
  assign new_n26295_ = ~new_n25665_ & ~new_n26294_;
  assign new_n26296_ = ~new_n26292_ & new_n26295_;
  assign new_n26297_ = ~new_n25665_ & ~new_n26296_;
  assign new_n26298_ = \b[47]  & ~new_n25654_;
  assign new_n26299_ = ~new_n25652_ & new_n26298_;
  assign new_n26300_ = ~new_n25656_ & ~new_n26299_;
  assign new_n26301_ = ~new_n26297_ & new_n26300_;
  assign new_n26302_ = ~new_n25656_ & ~new_n26301_;
  assign new_n26303_ = \b[48]  & ~new_n25645_;
  assign new_n26304_ = ~new_n25643_ & new_n26303_;
  assign new_n26305_ = ~new_n25647_ & ~new_n26304_;
  assign new_n26306_ = ~new_n26302_ & new_n26305_;
  assign new_n26307_ = ~new_n25647_ & ~new_n26306_;
  assign new_n26308_ = \b[49]  & ~new_n25636_;
  assign new_n26309_ = ~new_n25634_ & new_n26308_;
  assign new_n26310_ = ~new_n25638_ & ~new_n26309_;
  assign new_n26311_ = ~new_n26307_ & new_n26310_;
  assign new_n26312_ = ~new_n25638_ & ~new_n26311_;
  assign new_n26313_ = \b[50]  & ~new_n25627_;
  assign new_n26314_ = ~new_n25625_ & new_n26313_;
  assign new_n26315_ = ~new_n25629_ & ~new_n26314_;
  assign new_n26316_ = ~new_n26312_ & new_n26315_;
  assign new_n26317_ = ~new_n25629_ & ~new_n26316_;
  assign new_n26318_ = \b[51]  & ~new_n25618_;
  assign new_n26319_ = ~new_n25616_ & new_n26318_;
  assign new_n26320_ = ~new_n25620_ & ~new_n26319_;
  assign new_n26321_ = ~new_n26317_ & new_n26320_;
  assign new_n26322_ = ~new_n25620_ & ~new_n26321_;
  assign new_n26323_ = \b[52]  & ~new_n25609_;
  assign new_n26324_ = ~new_n25607_ & new_n26323_;
  assign new_n26325_ = ~new_n25611_ & ~new_n26324_;
  assign new_n26326_ = ~new_n26322_ & new_n26325_;
  assign new_n26327_ = ~new_n25611_ & ~new_n26326_;
  assign new_n26328_ = \b[53]  & ~new_n25600_;
  assign new_n26329_ = ~new_n25598_ & new_n26328_;
  assign new_n26330_ = ~new_n25602_ & ~new_n26329_;
  assign new_n26331_ = ~new_n26327_ & new_n26330_;
  assign new_n26332_ = ~new_n25602_ & ~new_n26331_;
  assign new_n26333_ = \b[54]  & ~new_n25591_;
  assign new_n26334_ = ~new_n25589_ & new_n26333_;
  assign new_n26335_ = ~new_n25593_ & ~new_n26334_;
  assign new_n26336_ = ~new_n26332_ & new_n26335_;
  assign new_n26337_ = ~new_n25593_ & ~new_n26336_;
  assign new_n26338_ = \b[55]  & ~new_n25582_;
  assign new_n26339_ = ~new_n25580_ & new_n26338_;
  assign new_n26340_ = ~new_n25584_ & ~new_n26339_;
  assign new_n26341_ = ~new_n26337_ & new_n26340_;
  assign new_n26342_ = ~new_n25584_ & ~new_n26341_;
  assign new_n26343_ = \b[56]  & ~new_n25573_;
  assign new_n26344_ = ~new_n25571_ & new_n26343_;
  assign new_n26345_ = ~new_n25575_ & ~new_n26344_;
  assign new_n26346_ = ~new_n26342_ & new_n26345_;
  assign new_n26347_ = ~new_n25575_ & ~new_n26346_;
  assign new_n26348_ = \b[57]  & ~new_n25564_;
  assign new_n26349_ = ~new_n25562_ & new_n26348_;
  assign new_n26350_ = ~new_n25566_ & ~new_n26349_;
  assign new_n26351_ = ~new_n26347_ & new_n26350_;
  assign new_n26352_ = ~new_n25566_ & ~new_n26351_;
  assign new_n26353_ = \b[58]  & ~new_n25555_;
  assign new_n26354_ = ~new_n25553_ & new_n26353_;
  assign new_n26355_ = ~new_n25557_ & ~new_n26354_;
  assign new_n26356_ = ~new_n26352_ & new_n26355_;
  assign new_n26357_ = ~new_n25557_ & ~new_n26356_;
  assign new_n26358_ = \b[59]  & ~new_n25546_;
  assign new_n26359_ = ~new_n25544_ & new_n26358_;
  assign new_n26360_ = ~new_n25548_ & ~new_n26359_;
  assign new_n26361_ = ~new_n26357_ & new_n26360_;
  assign new_n26362_ = ~new_n25548_ & ~new_n26361_;
  assign new_n26363_ = ~new_n24721_ & ~new_n25534_;
  assign new_n26364_ = ~new_n25532_ & new_n26363_;
  assign new_n26365_ = ~new_n25520_ & new_n26364_;
  assign new_n26366_ = ~new_n25532_ & ~new_n25534_;
  assign new_n26367_ = ~new_n25521_ & ~new_n26366_;
  assign new_n26368_ = ~new_n26365_ & ~new_n26367_;
  assign new_n26369_ = \quotient[4]  & ~new_n26368_;
  assign new_n26370_ = ~new_n25531_ & ~new_n25538_;
  assign new_n26371_ = ~new_n25537_ & new_n26370_;
  assign new_n26372_ = ~new_n26369_ & ~new_n26371_;
  assign new_n26373_ = ~\b[60]  & ~new_n26372_;
  assign new_n26374_ = \b[60]  & ~new_n26371_;
  assign new_n26375_ = ~new_n26369_ & new_n26374_;
  assign new_n26376_ = new_n403_ & ~new_n26375_;
  assign new_n26377_ = ~new_n26373_ & new_n26376_;
  assign new_n26378_ = ~new_n26362_ & new_n26377_;
  assign new_n26379_ = new_n280_ & ~new_n26372_;
  assign \quotient[3]  = new_n26378_ | new_n26379_;
  assign new_n26381_ = ~new_n25557_ & new_n26360_;
  assign new_n26382_ = ~new_n26356_ & new_n26381_;
  assign new_n26383_ = ~new_n26357_ & ~new_n26360_;
  assign new_n26384_ = ~new_n26382_ & ~new_n26383_;
  assign new_n26385_ = \quotient[3]  & ~new_n26384_;
  assign new_n26386_ = ~new_n25547_ & ~new_n26379_;
  assign new_n26387_ = ~new_n26378_ & new_n26386_;
  assign new_n26388_ = ~new_n26385_ & ~new_n26387_;
  assign new_n26389_ = ~\b[60]  & ~new_n26388_;
  assign new_n26390_ = ~new_n25566_ & new_n26355_;
  assign new_n26391_ = ~new_n26351_ & new_n26390_;
  assign new_n26392_ = ~new_n26352_ & ~new_n26355_;
  assign new_n26393_ = ~new_n26391_ & ~new_n26392_;
  assign new_n26394_ = \quotient[3]  & ~new_n26393_;
  assign new_n26395_ = ~new_n25556_ & ~new_n26379_;
  assign new_n26396_ = ~new_n26378_ & new_n26395_;
  assign new_n26397_ = ~new_n26394_ & ~new_n26396_;
  assign new_n26398_ = ~\b[59]  & ~new_n26397_;
  assign new_n26399_ = ~new_n25575_ & new_n26350_;
  assign new_n26400_ = ~new_n26346_ & new_n26399_;
  assign new_n26401_ = ~new_n26347_ & ~new_n26350_;
  assign new_n26402_ = ~new_n26400_ & ~new_n26401_;
  assign new_n26403_ = \quotient[3]  & ~new_n26402_;
  assign new_n26404_ = ~new_n25565_ & ~new_n26379_;
  assign new_n26405_ = ~new_n26378_ & new_n26404_;
  assign new_n26406_ = ~new_n26403_ & ~new_n26405_;
  assign new_n26407_ = ~\b[58]  & ~new_n26406_;
  assign new_n26408_ = ~new_n25584_ & new_n26345_;
  assign new_n26409_ = ~new_n26341_ & new_n26408_;
  assign new_n26410_ = ~new_n26342_ & ~new_n26345_;
  assign new_n26411_ = ~new_n26409_ & ~new_n26410_;
  assign new_n26412_ = \quotient[3]  & ~new_n26411_;
  assign new_n26413_ = ~new_n25574_ & ~new_n26379_;
  assign new_n26414_ = ~new_n26378_ & new_n26413_;
  assign new_n26415_ = ~new_n26412_ & ~new_n26414_;
  assign new_n26416_ = ~\b[57]  & ~new_n26415_;
  assign new_n26417_ = ~new_n25593_ & new_n26340_;
  assign new_n26418_ = ~new_n26336_ & new_n26417_;
  assign new_n26419_ = ~new_n26337_ & ~new_n26340_;
  assign new_n26420_ = ~new_n26418_ & ~new_n26419_;
  assign new_n26421_ = \quotient[3]  & ~new_n26420_;
  assign new_n26422_ = ~new_n25583_ & ~new_n26379_;
  assign new_n26423_ = ~new_n26378_ & new_n26422_;
  assign new_n26424_ = ~new_n26421_ & ~new_n26423_;
  assign new_n26425_ = ~\b[56]  & ~new_n26424_;
  assign new_n26426_ = ~new_n25602_ & new_n26335_;
  assign new_n26427_ = ~new_n26331_ & new_n26426_;
  assign new_n26428_ = ~new_n26332_ & ~new_n26335_;
  assign new_n26429_ = ~new_n26427_ & ~new_n26428_;
  assign new_n26430_ = \quotient[3]  & ~new_n26429_;
  assign new_n26431_ = ~new_n25592_ & ~new_n26379_;
  assign new_n26432_ = ~new_n26378_ & new_n26431_;
  assign new_n26433_ = ~new_n26430_ & ~new_n26432_;
  assign new_n26434_ = ~\b[55]  & ~new_n26433_;
  assign new_n26435_ = ~new_n25611_ & new_n26330_;
  assign new_n26436_ = ~new_n26326_ & new_n26435_;
  assign new_n26437_ = ~new_n26327_ & ~new_n26330_;
  assign new_n26438_ = ~new_n26436_ & ~new_n26437_;
  assign new_n26439_ = \quotient[3]  & ~new_n26438_;
  assign new_n26440_ = ~new_n25601_ & ~new_n26379_;
  assign new_n26441_ = ~new_n26378_ & new_n26440_;
  assign new_n26442_ = ~new_n26439_ & ~new_n26441_;
  assign new_n26443_ = ~\b[54]  & ~new_n26442_;
  assign new_n26444_ = ~new_n25620_ & new_n26325_;
  assign new_n26445_ = ~new_n26321_ & new_n26444_;
  assign new_n26446_ = ~new_n26322_ & ~new_n26325_;
  assign new_n26447_ = ~new_n26445_ & ~new_n26446_;
  assign new_n26448_ = \quotient[3]  & ~new_n26447_;
  assign new_n26449_ = ~new_n25610_ & ~new_n26379_;
  assign new_n26450_ = ~new_n26378_ & new_n26449_;
  assign new_n26451_ = ~new_n26448_ & ~new_n26450_;
  assign new_n26452_ = ~\b[53]  & ~new_n26451_;
  assign new_n26453_ = ~new_n25629_ & new_n26320_;
  assign new_n26454_ = ~new_n26316_ & new_n26453_;
  assign new_n26455_ = ~new_n26317_ & ~new_n26320_;
  assign new_n26456_ = ~new_n26454_ & ~new_n26455_;
  assign new_n26457_ = \quotient[3]  & ~new_n26456_;
  assign new_n26458_ = ~new_n25619_ & ~new_n26379_;
  assign new_n26459_ = ~new_n26378_ & new_n26458_;
  assign new_n26460_ = ~new_n26457_ & ~new_n26459_;
  assign new_n26461_ = ~\b[52]  & ~new_n26460_;
  assign new_n26462_ = ~new_n25638_ & new_n26315_;
  assign new_n26463_ = ~new_n26311_ & new_n26462_;
  assign new_n26464_ = ~new_n26312_ & ~new_n26315_;
  assign new_n26465_ = ~new_n26463_ & ~new_n26464_;
  assign new_n26466_ = \quotient[3]  & ~new_n26465_;
  assign new_n26467_ = ~new_n25628_ & ~new_n26379_;
  assign new_n26468_ = ~new_n26378_ & new_n26467_;
  assign new_n26469_ = ~new_n26466_ & ~new_n26468_;
  assign new_n26470_ = ~\b[51]  & ~new_n26469_;
  assign new_n26471_ = ~new_n25647_ & new_n26310_;
  assign new_n26472_ = ~new_n26306_ & new_n26471_;
  assign new_n26473_ = ~new_n26307_ & ~new_n26310_;
  assign new_n26474_ = ~new_n26472_ & ~new_n26473_;
  assign new_n26475_ = \quotient[3]  & ~new_n26474_;
  assign new_n26476_ = ~new_n25637_ & ~new_n26379_;
  assign new_n26477_ = ~new_n26378_ & new_n26476_;
  assign new_n26478_ = ~new_n26475_ & ~new_n26477_;
  assign new_n26479_ = ~\b[50]  & ~new_n26478_;
  assign new_n26480_ = ~new_n25656_ & new_n26305_;
  assign new_n26481_ = ~new_n26301_ & new_n26480_;
  assign new_n26482_ = ~new_n26302_ & ~new_n26305_;
  assign new_n26483_ = ~new_n26481_ & ~new_n26482_;
  assign new_n26484_ = \quotient[3]  & ~new_n26483_;
  assign new_n26485_ = ~new_n25646_ & ~new_n26379_;
  assign new_n26486_ = ~new_n26378_ & new_n26485_;
  assign new_n26487_ = ~new_n26484_ & ~new_n26486_;
  assign new_n26488_ = ~\b[49]  & ~new_n26487_;
  assign new_n26489_ = ~new_n25665_ & new_n26300_;
  assign new_n26490_ = ~new_n26296_ & new_n26489_;
  assign new_n26491_ = ~new_n26297_ & ~new_n26300_;
  assign new_n26492_ = ~new_n26490_ & ~new_n26491_;
  assign new_n26493_ = \quotient[3]  & ~new_n26492_;
  assign new_n26494_ = ~new_n25655_ & ~new_n26379_;
  assign new_n26495_ = ~new_n26378_ & new_n26494_;
  assign new_n26496_ = ~new_n26493_ & ~new_n26495_;
  assign new_n26497_ = ~\b[48]  & ~new_n26496_;
  assign new_n26498_ = ~new_n25674_ & new_n26295_;
  assign new_n26499_ = ~new_n26291_ & new_n26498_;
  assign new_n26500_ = ~new_n26292_ & ~new_n26295_;
  assign new_n26501_ = ~new_n26499_ & ~new_n26500_;
  assign new_n26502_ = \quotient[3]  & ~new_n26501_;
  assign new_n26503_ = ~new_n25664_ & ~new_n26379_;
  assign new_n26504_ = ~new_n26378_ & new_n26503_;
  assign new_n26505_ = ~new_n26502_ & ~new_n26504_;
  assign new_n26506_ = ~\b[47]  & ~new_n26505_;
  assign new_n26507_ = ~new_n25683_ & new_n26290_;
  assign new_n26508_ = ~new_n26286_ & new_n26507_;
  assign new_n26509_ = ~new_n26287_ & ~new_n26290_;
  assign new_n26510_ = ~new_n26508_ & ~new_n26509_;
  assign new_n26511_ = \quotient[3]  & ~new_n26510_;
  assign new_n26512_ = ~new_n25673_ & ~new_n26379_;
  assign new_n26513_ = ~new_n26378_ & new_n26512_;
  assign new_n26514_ = ~new_n26511_ & ~new_n26513_;
  assign new_n26515_ = ~\b[46]  & ~new_n26514_;
  assign new_n26516_ = ~new_n25692_ & new_n26285_;
  assign new_n26517_ = ~new_n26281_ & new_n26516_;
  assign new_n26518_ = ~new_n26282_ & ~new_n26285_;
  assign new_n26519_ = ~new_n26517_ & ~new_n26518_;
  assign new_n26520_ = \quotient[3]  & ~new_n26519_;
  assign new_n26521_ = ~new_n25682_ & ~new_n26379_;
  assign new_n26522_ = ~new_n26378_ & new_n26521_;
  assign new_n26523_ = ~new_n26520_ & ~new_n26522_;
  assign new_n26524_ = ~\b[45]  & ~new_n26523_;
  assign new_n26525_ = ~new_n25701_ & new_n26280_;
  assign new_n26526_ = ~new_n26276_ & new_n26525_;
  assign new_n26527_ = ~new_n26277_ & ~new_n26280_;
  assign new_n26528_ = ~new_n26526_ & ~new_n26527_;
  assign new_n26529_ = \quotient[3]  & ~new_n26528_;
  assign new_n26530_ = ~new_n25691_ & ~new_n26379_;
  assign new_n26531_ = ~new_n26378_ & new_n26530_;
  assign new_n26532_ = ~new_n26529_ & ~new_n26531_;
  assign new_n26533_ = ~\b[44]  & ~new_n26532_;
  assign new_n26534_ = ~new_n25710_ & new_n26275_;
  assign new_n26535_ = ~new_n26271_ & new_n26534_;
  assign new_n26536_ = ~new_n26272_ & ~new_n26275_;
  assign new_n26537_ = ~new_n26535_ & ~new_n26536_;
  assign new_n26538_ = \quotient[3]  & ~new_n26537_;
  assign new_n26539_ = ~new_n25700_ & ~new_n26379_;
  assign new_n26540_ = ~new_n26378_ & new_n26539_;
  assign new_n26541_ = ~new_n26538_ & ~new_n26540_;
  assign new_n26542_ = ~\b[43]  & ~new_n26541_;
  assign new_n26543_ = ~new_n25719_ & new_n26270_;
  assign new_n26544_ = ~new_n26266_ & new_n26543_;
  assign new_n26545_ = ~new_n26267_ & ~new_n26270_;
  assign new_n26546_ = ~new_n26544_ & ~new_n26545_;
  assign new_n26547_ = \quotient[3]  & ~new_n26546_;
  assign new_n26548_ = ~new_n25709_ & ~new_n26379_;
  assign new_n26549_ = ~new_n26378_ & new_n26548_;
  assign new_n26550_ = ~new_n26547_ & ~new_n26549_;
  assign new_n26551_ = ~\b[42]  & ~new_n26550_;
  assign new_n26552_ = ~new_n25728_ & new_n26265_;
  assign new_n26553_ = ~new_n26261_ & new_n26552_;
  assign new_n26554_ = ~new_n26262_ & ~new_n26265_;
  assign new_n26555_ = ~new_n26553_ & ~new_n26554_;
  assign new_n26556_ = \quotient[3]  & ~new_n26555_;
  assign new_n26557_ = ~new_n25718_ & ~new_n26379_;
  assign new_n26558_ = ~new_n26378_ & new_n26557_;
  assign new_n26559_ = ~new_n26556_ & ~new_n26558_;
  assign new_n26560_ = ~\b[41]  & ~new_n26559_;
  assign new_n26561_ = ~new_n25737_ & new_n26260_;
  assign new_n26562_ = ~new_n26256_ & new_n26561_;
  assign new_n26563_ = ~new_n26257_ & ~new_n26260_;
  assign new_n26564_ = ~new_n26562_ & ~new_n26563_;
  assign new_n26565_ = \quotient[3]  & ~new_n26564_;
  assign new_n26566_ = ~new_n25727_ & ~new_n26379_;
  assign new_n26567_ = ~new_n26378_ & new_n26566_;
  assign new_n26568_ = ~new_n26565_ & ~new_n26567_;
  assign new_n26569_ = ~\b[40]  & ~new_n26568_;
  assign new_n26570_ = ~new_n25746_ & new_n26255_;
  assign new_n26571_ = ~new_n26251_ & new_n26570_;
  assign new_n26572_ = ~new_n26252_ & ~new_n26255_;
  assign new_n26573_ = ~new_n26571_ & ~new_n26572_;
  assign new_n26574_ = \quotient[3]  & ~new_n26573_;
  assign new_n26575_ = ~new_n25736_ & ~new_n26379_;
  assign new_n26576_ = ~new_n26378_ & new_n26575_;
  assign new_n26577_ = ~new_n26574_ & ~new_n26576_;
  assign new_n26578_ = ~\b[39]  & ~new_n26577_;
  assign new_n26579_ = ~new_n25755_ & new_n26250_;
  assign new_n26580_ = ~new_n26246_ & new_n26579_;
  assign new_n26581_ = ~new_n26247_ & ~new_n26250_;
  assign new_n26582_ = ~new_n26580_ & ~new_n26581_;
  assign new_n26583_ = \quotient[3]  & ~new_n26582_;
  assign new_n26584_ = ~new_n25745_ & ~new_n26379_;
  assign new_n26585_ = ~new_n26378_ & new_n26584_;
  assign new_n26586_ = ~new_n26583_ & ~new_n26585_;
  assign new_n26587_ = ~\b[38]  & ~new_n26586_;
  assign new_n26588_ = ~new_n25764_ & new_n26245_;
  assign new_n26589_ = ~new_n26241_ & new_n26588_;
  assign new_n26590_ = ~new_n26242_ & ~new_n26245_;
  assign new_n26591_ = ~new_n26589_ & ~new_n26590_;
  assign new_n26592_ = \quotient[3]  & ~new_n26591_;
  assign new_n26593_ = ~new_n25754_ & ~new_n26379_;
  assign new_n26594_ = ~new_n26378_ & new_n26593_;
  assign new_n26595_ = ~new_n26592_ & ~new_n26594_;
  assign new_n26596_ = ~\b[37]  & ~new_n26595_;
  assign new_n26597_ = ~new_n25773_ & new_n26240_;
  assign new_n26598_ = ~new_n26236_ & new_n26597_;
  assign new_n26599_ = ~new_n26237_ & ~new_n26240_;
  assign new_n26600_ = ~new_n26598_ & ~new_n26599_;
  assign new_n26601_ = \quotient[3]  & ~new_n26600_;
  assign new_n26602_ = ~new_n25763_ & ~new_n26379_;
  assign new_n26603_ = ~new_n26378_ & new_n26602_;
  assign new_n26604_ = ~new_n26601_ & ~new_n26603_;
  assign new_n26605_ = ~\b[36]  & ~new_n26604_;
  assign new_n26606_ = ~new_n25782_ & new_n26235_;
  assign new_n26607_ = ~new_n26231_ & new_n26606_;
  assign new_n26608_ = ~new_n26232_ & ~new_n26235_;
  assign new_n26609_ = ~new_n26607_ & ~new_n26608_;
  assign new_n26610_ = \quotient[3]  & ~new_n26609_;
  assign new_n26611_ = ~new_n25772_ & ~new_n26379_;
  assign new_n26612_ = ~new_n26378_ & new_n26611_;
  assign new_n26613_ = ~new_n26610_ & ~new_n26612_;
  assign new_n26614_ = ~\b[35]  & ~new_n26613_;
  assign new_n26615_ = ~new_n25791_ & new_n26230_;
  assign new_n26616_ = ~new_n26226_ & new_n26615_;
  assign new_n26617_ = ~new_n26227_ & ~new_n26230_;
  assign new_n26618_ = ~new_n26616_ & ~new_n26617_;
  assign new_n26619_ = \quotient[3]  & ~new_n26618_;
  assign new_n26620_ = ~new_n25781_ & ~new_n26379_;
  assign new_n26621_ = ~new_n26378_ & new_n26620_;
  assign new_n26622_ = ~new_n26619_ & ~new_n26621_;
  assign new_n26623_ = ~\b[34]  & ~new_n26622_;
  assign new_n26624_ = ~new_n25800_ & new_n26225_;
  assign new_n26625_ = ~new_n26221_ & new_n26624_;
  assign new_n26626_ = ~new_n26222_ & ~new_n26225_;
  assign new_n26627_ = ~new_n26625_ & ~new_n26626_;
  assign new_n26628_ = \quotient[3]  & ~new_n26627_;
  assign new_n26629_ = ~new_n25790_ & ~new_n26379_;
  assign new_n26630_ = ~new_n26378_ & new_n26629_;
  assign new_n26631_ = ~new_n26628_ & ~new_n26630_;
  assign new_n26632_ = ~\b[33]  & ~new_n26631_;
  assign new_n26633_ = ~new_n25809_ & new_n26220_;
  assign new_n26634_ = ~new_n26216_ & new_n26633_;
  assign new_n26635_ = ~new_n26217_ & ~new_n26220_;
  assign new_n26636_ = ~new_n26634_ & ~new_n26635_;
  assign new_n26637_ = \quotient[3]  & ~new_n26636_;
  assign new_n26638_ = ~new_n25799_ & ~new_n26379_;
  assign new_n26639_ = ~new_n26378_ & new_n26638_;
  assign new_n26640_ = ~new_n26637_ & ~new_n26639_;
  assign new_n26641_ = ~\b[32]  & ~new_n26640_;
  assign new_n26642_ = ~new_n25818_ & new_n26215_;
  assign new_n26643_ = ~new_n26211_ & new_n26642_;
  assign new_n26644_ = ~new_n26212_ & ~new_n26215_;
  assign new_n26645_ = ~new_n26643_ & ~new_n26644_;
  assign new_n26646_ = \quotient[3]  & ~new_n26645_;
  assign new_n26647_ = ~new_n25808_ & ~new_n26379_;
  assign new_n26648_ = ~new_n26378_ & new_n26647_;
  assign new_n26649_ = ~new_n26646_ & ~new_n26648_;
  assign new_n26650_ = ~\b[31]  & ~new_n26649_;
  assign new_n26651_ = ~new_n25827_ & new_n26210_;
  assign new_n26652_ = ~new_n26206_ & new_n26651_;
  assign new_n26653_ = ~new_n26207_ & ~new_n26210_;
  assign new_n26654_ = ~new_n26652_ & ~new_n26653_;
  assign new_n26655_ = \quotient[3]  & ~new_n26654_;
  assign new_n26656_ = ~new_n25817_ & ~new_n26379_;
  assign new_n26657_ = ~new_n26378_ & new_n26656_;
  assign new_n26658_ = ~new_n26655_ & ~new_n26657_;
  assign new_n26659_ = ~\b[30]  & ~new_n26658_;
  assign new_n26660_ = ~new_n25836_ & new_n26205_;
  assign new_n26661_ = ~new_n26201_ & new_n26660_;
  assign new_n26662_ = ~new_n26202_ & ~new_n26205_;
  assign new_n26663_ = ~new_n26661_ & ~new_n26662_;
  assign new_n26664_ = \quotient[3]  & ~new_n26663_;
  assign new_n26665_ = ~new_n25826_ & ~new_n26379_;
  assign new_n26666_ = ~new_n26378_ & new_n26665_;
  assign new_n26667_ = ~new_n26664_ & ~new_n26666_;
  assign new_n26668_ = ~\b[29]  & ~new_n26667_;
  assign new_n26669_ = ~new_n25845_ & new_n26200_;
  assign new_n26670_ = ~new_n26196_ & new_n26669_;
  assign new_n26671_ = ~new_n26197_ & ~new_n26200_;
  assign new_n26672_ = ~new_n26670_ & ~new_n26671_;
  assign new_n26673_ = \quotient[3]  & ~new_n26672_;
  assign new_n26674_ = ~new_n25835_ & ~new_n26379_;
  assign new_n26675_ = ~new_n26378_ & new_n26674_;
  assign new_n26676_ = ~new_n26673_ & ~new_n26675_;
  assign new_n26677_ = ~\b[28]  & ~new_n26676_;
  assign new_n26678_ = ~new_n25854_ & new_n26195_;
  assign new_n26679_ = ~new_n26191_ & new_n26678_;
  assign new_n26680_ = ~new_n26192_ & ~new_n26195_;
  assign new_n26681_ = ~new_n26679_ & ~new_n26680_;
  assign new_n26682_ = \quotient[3]  & ~new_n26681_;
  assign new_n26683_ = ~new_n25844_ & ~new_n26379_;
  assign new_n26684_ = ~new_n26378_ & new_n26683_;
  assign new_n26685_ = ~new_n26682_ & ~new_n26684_;
  assign new_n26686_ = ~\b[27]  & ~new_n26685_;
  assign new_n26687_ = ~new_n25863_ & new_n26190_;
  assign new_n26688_ = ~new_n26186_ & new_n26687_;
  assign new_n26689_ = ~new_n26187_ & ~new_n26190_;
  assign new_n26690_ = ~new_n26688_ & ~new_n26689_;
  assign new_n26691_ = \quotient[3]  & ~new_n26690_;
  assign new_n26692_ = ~new_n25853_ & ~new_n26379_;
  assign new_n26693_ = ~new_n26378_ & new_n26692_;
  assign new_n26694_ = ~new_n26691_ & ~new_n26693_;
  assign new_n26695_ = ~\b[26]  & ~new_n26694_;
  assign new_n26696_ = ~new_n25872_ & new_n26185_;
  assign new_n26697_ = ~new_n26181_ & new_n26696_;
  assign new_n26698_ = ~new_n26182_ & ~new_n26185_;
  assign new_n26699_ = ~new_n26697_ & ~new_n26698_;
  assign new_n26700_ = \quotient[3]  & ~new_n26699_;
  assign new_n26701_ = ~new_n25862_ & ~new_n26379_;
  assign new_n26702_ = ~new_n26378_ & new_n26701_;
  assign new_n26703_ = ~new_n26700_ & ~new_n26702_;
  assign new_n26704_ = ~\b[25]  & ~new_n26703_;
  assign new_n26705_ = ~new_n25881_ & new_n26180_;
  assign new_n26706_ = ~new_n26176_ & new_n26705_;
  assign new_n26707_ = ~new_n26177_ & ~new_n26180_;
  assign new_n26708_ = ~new_n26706_ & ~new_n26707_;
  assign new_n26709_ = \quotient[3]  & ~new_n26708_;
  assign new_n26710_ = ~new_n25871_ & ~new_n26379_;
  assign new_n26711_ = ~new_n26378_ & new_n26710_;
  assign new_n26712_ = ~new_n26709_ & ~new_n26711_;
  assign new_n26713_ = ~\b[24]  & ~new_n26712_;
  assign new_n26714_ = ~new_n25890_ & new_n26175_;
  assign new_n26715_ = ~new_n26171_ & new_n26714_;
  assign new_n26716_ = ~new_n26172_ & ~new_n26175_;
  assign new_n26717_ = ~new_n26715_ & ~new_n26716_;
  assign new_n26718_ = \quotient[3]  & ~new_n26717_;
  assign new_n26719_ = ~new_n25880_ & ~new_n26379_;
  assign new_n26720_ = ~new_n26378_ & new_n26719_;
  assign new_n26721_ = ~new_n26718_ & ~new_n26720_;
  assign new_n26722_ = ~\b[23]  & ~new_n26721_;
  assign new_n26723_ = ~new_n25899_ & new_n26170_;
  assign new_n26724_ = ~new_n26166_ & new_n26723_;
  assign new_n26725_ = ~new_n26167_ & ~new_n26170_;
  assign new_n26726_ = ~new_n26724_ & ~new_n26725_;
  assign new_n26727_ = \quotient[3]  & ~new_n26726_;
  assign new_n26728_ = ~new_n25889_ & ~new_n26379_;
  assign new_n26729_ = ~new_n26378_ & new_n26728_;
  assign new_n26730_ = ~new_n26727_ & ~new_n26729_;
  assign new_n26731_ = ~\b[22]  & ~new_n26730_;
  assign new_n26732_ = ~new_n25908_ & new_n26165_;
  assign new_n26733_ = ~new_n26161_ & new_n26732_;
  assign new_n26734_ = ~new_n26162_ & ~new_n26165_;
  assign new_n26735_ = ~new_n26733_ & ~new_n26734_;
  assign new_n26736_ = \quotient[3]  & ~new_n26735_;
  assign new_n26737_ = ~new_n25898_ & ~new_n26379_;
  assign new_n26738_ = ~new_n26378_ & new_n26737_;
  assign new_n26739_ = ~new_n26736_ & ~new_n26738_;
  assign new_n26740_ = ~\b[21]  & ~new_n26739_;
  assign new_n26741_ = ~new_n25917_ & new_n26160_;
  assign new_n26742_ = ~new_n26156_ & new_n26741_;
  assign new_n26743_ = ~new_n26157_ & ~new_n26160_;
  assign new_n26744_ = ~new_n26742_ & ~new_n26743_;
  assign new_n26745_ = \quotient[3]  & ~new_n26744_;
  assign new_n26746_ = ~new_n25907_ & ~new_n26379_;
  assign new_n26747_ = ~new_n26378_ & new_n26746_;
  assign new_n26748_ = ~new_n26745_ & ~new_n26747_;
  assign new_n26749_ = ~\b[20]  & ~new_n26748_;
  assign new_n26750_ = ~new_n25926_ & new_n26155_;
  assign new_n26751_ = ~new_n26151_ & new_n26750_;
  assign new_n26752_ = ~new_n26152_ & ~new_n26155_;
  assign new_n26753_ = ~new_n26751_ & ~new_n26752_;
  assign new_n26754_ = \quotient[3]  & ~new_n26753_;
  assign new_n26755_ = ~new_n25916_ & ~new_n26379_;
  assign new_n26756_ = ~new_n26378_ & new_n26755_;
  assign new_n26757_ = ~new_n26754_ & ~new_n26756_;
  assign new_n26758_ = ~\b[19]  & ~new_n26757_;
  assign new_n26759_ = ~new_n25935_ & new_n26150_;
  assign new_n26760_ = ~new_n26146_ & new_n26759_;
  assign new_n26761_ = ~new_n26147_ & ~new_n26150_;
  assign new_n26762_ = ~new_n26760_ & ~new_n26761_;
  assign new_n26763_ = \quotient[3]  & ~new_n26762_;
  assign new_n26764_ = ~new_n25925_ & ~new_n26379_;
  assign new_n26765_ = ~new_n26378_ & new_n26764_;
  assign new_n26766_ = ~new_n26763_ & ~new_n26765_;
  assign new_n26767_ = ~\b[18]  & ~new_n26766_;
  assign new_n26768_ = ~new_n25944_ & new_n26145_;
  assign new_n26769_ = ~new_n26141_ & new_n26768_;
  assign new_n26770_ = ~new_n26142_ & ~new_n26145_;
  assign new_n26771_ = ~new_n26769_ & ~new_n26770_;
  assign new_n26772_ = \quotient[3]  & ~new_n26771_;
  assign new_n26773_ = ~new_n25934_ & ~new_n26379_;
  assign new_n26774_ = ~new_n26378_ & new_n26773_;
  assign new_n26775_ = ~new_n26772_ & ~new_n26774_;
  assign new_n26776_ = ~\b[17]  & ~new_n26775_;
  assign new_n26777_ = ~new_n25953_ & new_n26140_;
  assign new_n26778_ = ~new_n26136_ & new_n26777_;
  assign new_n26779_ = ~new_n26137_ & ~new_n26140_;
  assign new_n26780_ = ~new_n26778_ & ~new_n26779_;
  assign new_n26781_ = \quotient[3]  & ~new_n26780_;
  assign new_n26782_ = ~new_n25943_ & ~new_n26379_;
  assign new_n26783_ = ~new_n26378_ & new_n26782_;
  assign new_n26784_ = ~new_n26781_ & ~new_n26783_;
  assign new_n26785_ = ~\b[16]  & ~new_n26784_;
  assign new_n26786_ = ~new_n25962_ & new_n26135_;
  assign new_n26787_ = ~new_n26131_ & new_n26786_;
  assign new_n26788_ = ~new_n26132_ & ~new_n26135_;
  assign new_n26789_ = ~new_n26787_ & ~new_n26788_;
  assign new_n26790_ = \quotient[3]  & ~new_n26789_;
  assign new_n26791_ = ~new_n25952_ & ~new_n26379_;
  assign new_n26792_ = ~new_n26378_ & new_n26791_;
  assign new_n26793_ = ~new_n26790_ & ~new_n26792_;
  assign new_n26794_ = ~\b[15]  & ~new_n26793_;
  assign new_n26795_ = ~new_n25971_ & new_n26130_;
  assign new_n26796_ = ~new_n26126_ & new_n26795_;
  assign new_n26797_ = ~new_n26127_ & ~new_n26130_;
  assign new_n26798_ = ~new_n26796_ & ~new_n26797_;
  assign new_n26799_ = \quotient[3]  & ~new_n26798_;
  assign new_n26800_ = ~new_n25961_ & ~new_n26379_;
  assign new_n26801_ = ~new_n26378_ & new_n26800_;
  assign new_n26802_ = ~new_n26799_ & ~new_n26801_;
  assign new_n26803_ = ~\b[14]  & ~new_n26802_;
  assign new_n26804_ = ~new_n25980_ & new_n26125_;
  assign new_n26805_ = ~new_n26121_ & new_n26804_;
  assign new_n26806_ = ~new_n26122_ & ~new_n26125_;
  assign new_n26807_ = ~new_n26805_ & ~new_n26806_;
  assign new_n26808_ = \quotient[3]  & ~new_n26807_;
  assign new_n26809_ = ~new_n25970_ & ~new_n26379_;
  assign new_n26810_ = ~new_n26378_ & new_n26809_;
  assign new_n26811_ = ~new_n26808_ & ~new_n26810_;
  assign new_n26812_ = ~\b[13]  & ~new_n26811_;
  assign new_n26813_ = ~new_n25989_ & new_n26120_;
  assign new_n26814_ = ~new_n26116_ & new_n26813_;
  assign new_n26815_ = ~new_n26117_ & ~new_n26120_;
  assign new_n26816_ = ~new_n26814_ & ~new_n26815_;
  assign new_n26817_ = \quotient[3]  & ~new_n26816_;
  assign new_n26818_ = ~new_n25979_ & ~new_n26379_;
  assign new_n26819_ = ~new_n26378_ & new_n26818_;
  assign new_n26820_ = ~new_n26817_ & ~new_n26819_;
  assign new_n26821_ = ~\b[12]  & ~new_n26820_;
  assign new_n26822_ = ~new_n25998_ & new_n26115_;
  assign new_n26823_ = ~new_n26111_ & new_n26822_;
  assign new_n26824_ = ~new_n26112_ & ~new_n26115_;
  assign new_n26825_ = ~new_n26823_ & ~new_n26824_;
  assign new_n26826_ = \quotient[3]  & ~new_n26825_;
  assign new_n26827_ = ~new_n25988_ & ~new_n26379_;
  assign new_n26828_ = ~new_n26378_ & new_n26827_;
  assign new_n26829_ = ~new_n26826_ & ~new_n26828_;
  assign new_n26830_ = ~\b[11]  & ~new_n26829_;
  assign new_n26831_ = ~new_n26007_ & new_n26110_;
  assign new_n26832_ = ~new_n26106_ & new_n26831_;
  assign new_n26833_ = ~new_n26107_ & ~new_n26110_;
  assign new_n26834_ = ~new_n26832_ & ~new_n26833_;
  assign new_n26835_ = \quotient[3]  & ~new_n26834_;
  assign new_n26836_ = ~new_n25997_ & ~new_n26379_;
  assign new_n26837_ = ~new_n26378_ & new_n26836_;
  assign new_n26838_ = ~new_n26835_ & ~new_n26837_;
  assign new_n26839_ = ~\b[10]  & ~new_n26838_;
  assign new_n26840_ = ~new_n26016_ & new_n26105_;
  assign new_n26841_ = ~new_n26101_ & new_n26840_;
  assign new_n26842_ = ~new_n26102_ & ~new_n26105_;
  assign new_n26843_ = ~new_n26841_ & ~new_n26842_;
  assign new_n26844_ = \quotient[3]  & ~new_n26843_;
  assign new_n26845_ = ~new_n26006_ & ~new_n26379_;
  assign new_n26846_ = ~new_n26378_ & new_n26845_;
  assign new_n26847_ = ~new_n26844_ & ~new_n26846_;
  assign new_n26848_ = ~\b[9]  & ~new_n26847_;
  assign new_n26849_ = ~new_n26025_ & new_n26100_;
  assign new_n26850_ = ~new_n26096_ & new_n26849_;
  assign new_n26851_ = ~new_n26097_ & ~new_n26100_;
  assign new_n26852_ = ~new_n26850_ & ~new_n26851_;
  assign new_n26853_ = \quotient[3]  & ~new_n26852_;
  assign new_n26854_ = ~new_n26015_ & ~new_n26379_;
  assign new_n26855_ = ~new_n26378_ & new_n26854_;
  assign new_n26856_ = ~new_n26853_ & ~new_n26855_;
  assign new_n26857_ = ~\b[8]  & ~new_n26856_;
  assign new_n26858_ = ~new_n26034_ & new_n26095_;
  assign new_n26859_ = ~new_n26091_ & new_n26858_;
  assign new_n26860_ = ~new_n26092_ & ~new_n26095_;
  assign new_n26861_ = ~new_n26859_ & ~new_n26860_;
  assign new_n26862_ = \quotient[3]  & ~new_n26861_;
  assign new_n26863_ = ~new_n26024_ & ~new_n26379_;
  assign new_n26864_ = ~new_n26378_ & new_n26863_;
  assign new_n26865_ = ~new_n26862_ & ~new_n26864_;
  assign new_n26866_ = ~\b[7]  & ~new_n26865_;
  assign new_n26867_ = ~new_n26043_ & new_n26090_;
  assign new_n26868_ = ~new_n26086_ & new_n26867_;
  assign new_n26869_ = ~new_n26087_ & ~new_n26090_;
  assign new_n26870_ = ~new_n26868_ & ~new_n26869_;
  assign new_n26871_ = \quotient[3]  & ~new_n26870_;
  assign new_n26872_ = ~new_n26033_ & ~new_n26379_;
  assign new_n26873_ = ~new_n26378_ & new_n26872_;
  assign new_n26874_ = ~new_n26871_ & ~new_n26873_;
  assign new_n26875_ = ~\b[6]  & ~new_n26874_;
  assign new_n26876_ = ~new_n26052_ & new_n26085_;
  assign new_n26877_ = ~new_n26081_ & new_n26876_;
  assign new_n26878_ = ~new_n26082_ & ~new_n26085_;
  assign new_n26879_ = ~new_n26877_ & ~new_n26878_;
  assign new_n26880_ = \quotient[3]  & ~new_n26879_;
  assign new_n26881_ = ~new_n26042_ & ~new_n26379_;
  assign new_n26882_ = ~new_n26378_ & new_n26881_;
  assign new_n26883_ = ~new_n26880_ & ~new_n26882_;
  assign new_n26884_ = ~\b[5]  & ~new_n26883_;
  assign new_n26885_ = ~new_n26060_ & new_n26080_;
  assign new_n26886_ = ~new_n26076_ & new_n26885_;
  assign new_n26887_ = ~new_n26077_ & ~new_n26080_;
  assign new_n26888_ = ~new_n26886_ & ~new_n26887_;
  assign new_n26889_ = \quotient[3]  & ~new_n26888_;
  assign new_n26890_ = ~new_n26051_ & ~new_n26379_;
  assign new_n26891_ = ~new_n26378_ & new_n26890_;
  assign new_n26892_ = ~new_n26889_ & ~new_n26891_;
  assign new_n26893_ = ~\b[4]  & ~new_n26892_;
  assign new_n26894_ = ~new_n26071_ & new_n26075_;
  assign new_n26895_ = ~new_n26070_ & new_n26894_;
  assign new_n26896_ = ~new_n26072_ & ~new_n26075_;
  assign new_n26897_ = ~new_n26895_ & ~new_n26896_;
  assign new_n26898_ = \quotient[3]  & ~new_n26897_;
  assign new_n26899_ = ~new_n26059_ & ~new_n26379_;
  assign new_n26900_ = ~new_n26378_ & new_n26899_;
  assign new_n26901_ = ~new_n26898_ & ~new_n26900_;
  assign new_n26902_ = ~\b[3]  & ~new_n26901_;
  assign new_n26903_ = ~new_n26067_ & new_n26069_;
  assign new_n26904_ = ~new_n26065_ & new_n26903_;
  assign new_n26905_ = ~new_n26070_ & ~new_n26904_;
  assign new_n26906_ = \quotient[3]  & new_n26905_;
  assign new_n26907_ = ~new_n26064_ & ~new_n26379_;
  assign new_n26908_ = ~new_n26378_ & new_n26907_;
  assign new_n26909_ = ~new_n26906_ & ~new_n26908_;
  assign new_n26910_ = ~\b[2]  & ~new_n26909_;
  assign new_n26911_ = \b[0]  & \quotient[3] ;
  assign new_n26912_ = \a[3]  & ~new_n26911_;
  assign new_n26913_ = new_n26069_ & \quotient[3] ;
  assign new_n26914_ = ~new_n26912_ & ~new_n26913_;
  assign new_n26915_ = \b[1]  & ~new_n26914_;
  assign new_n26916_ = ~\b[1]  & ~new_n26913_;
  assign new_n26917_ = ~new_n26912_ & new_n26916_;
  assign new_n26918_ = ~new_n26915_ & ~new_n26917_;
  assign new_n26919_ = ~\a[2]  & \b[0] ;
  assign new_n26920_ = ~new_n26918_ & ~new_n26919_;
  assign new_n26921_ = ~\b[1]  & ~new_n26914_;
  assign new_n26922_ = ~new_n26920_ & ~new_n26921_;
  assign new_n26923_ = \b[2]  & ~new_n26908_;
  assign new_n26924_ = ~new_n26906_ & new_n26923_;
  assign new_n26925_ = ~new_n26910_ & ~new_n26924_;
  assign new_n26926_ = ~new_n26922_ & new_n26925_;
  assign new_n26927_ = ~new_n26910_ & ~new_n26926_;
  assign new_n26928_ = \b[3]  & ~new_n26900_;
  assign new_n26929_ = ~new_n26898_ & new_n26928_;
  assign new_n26930_ = ~new_n26902_ & ~new_n26929_;
  assign new_n26931_ = ~new_n26927_ & new_n26930_;
  assign new_n26932_ = ~new_n26902_ & ~new_n26931_;
  assign new_n26933_ = \b[4]  & ~new_n26891_;
  assign new_n26934_ = ~new_n26889_ & new_n26933_;
  assign new_n26935_ = ~new_n26893_ & ~new_n26934_;
  assign new_n26936_ = ~new_n26932_ & new_n26935_;
  assign new_n26937_ = ~new_n26893_ & ~new_n26936_;
  assign new_n26938_ = \b[5]  & ~new_n26882_;
  assign new_n26939_ = ~new_n26880_ & new_n26938_;
  assign new_n26940_ = ~new_n26884_ & ~new_n26939_;
  assign new_n26941_ = ~new_n26937_ & new_n26940_;
  assign new_n26942_ = ~new_n26884_ & ~new_n26941_;
  assign new_n26943_ = \b[6]  & ~new_n26873_;
  assign new_n26944_ = ~new_n26871_ & new_n26943_;
  assign new_n26945_ = ~new_n26875_ & ~new_n26944_;
  assign new_n26946_ = ~new_n26942_ & new_n26945_;
  assign new_n26947_ = ~new_n26875_ & ~new_n26946_;
  assign new_n26948_ = \b[7]  & ~new_n26864_;
  assign new_n26949_ = ~new_n26862_ & new_n26948_;
  assign new_n26950_ = ~new_n26866_ & ~new_n26949_;
  assign new_n26951_ = ~new_n26947_ & new_n26950_;
  assign new_n26952_ = ~new_n26866_ & ~new_n26951_;
  assign new_n26953_ = \b[8]  & ~new_n26855_;
  assign new_n26954_ = ~new_n26853_ & new_n26953_;
  assign new_n26955_ = ~new_n26857_ & ~new_n26954_;
  assign new_n26956_ = ~new_n26952_ & new_n26955_;
  assign new_n26957_ = ~new_n26857_ & ~new_n26956_;
  assign new_n26958_ = \b[9]  & ~new_n26846_;
  assign new_n26959_ = ~new_n26844_ & new_n26958_;
  assign new_n26960_ = ~new_n26848_ & ~new_n26959_;
  assign new_n26961_ = ~new_n26957_ & new_n26960_;
  assign new_n26962_ = ~new_n26848_ & ~new_n26961_;
  assign new_n26963_ = \b[10]  & ~new_n26837_;
  assign new_n26964_ = ~new_n26835_ & new_n26963_;
  assign new_n26965_ = ~new_n26839_ & ~new_n26964_;
  assign new_n26966_ = ~new_n26962_ & new_n26965_;
  assign new_n26967_ = ~new_n26839_ & ~new_n26966_;
  assign new_n26968_ = \b[11]  & ~new_n26828_;
  assign new_n26969_ = ~new_n26826_ & new_n26968_;
  assign new_n26970_ = ~new_n26830_ & ~new_n26969_;
  assign new_n26971_ = ~new_n26967_ & new_n26970_;
  assign new_n26972_ = ~new_n26830_ & ~new_n26971_;
  assign new_n26973_ = \b[12]  & ~new_n26819_;
  assign new_n26974_ = ~new_n26817_ & new_n26973_;
  assign new_n26975_ = ~new_n26821_ & ~new_n26974_;
  assign new_n26976_ = ~new_n26972_ & new_n26975_;
  assign new_n26977_ = ~new_n26821_ & ~new_n26976_;
  assign new_n26978_ = \b[13]  & ~new_n26810_;
  assign new_n26979_ = ~new_n26808_ & new_n26978_;
  assign new_n26980_ = ~new_n26812_ & ~new_n26979_;
  assign new_n26981_ = ~new_n26977_ & new_n26980_;
  assign new_n26982_ = ~new_n26812_ & ~new_n26981_;
  assign new_n26983_ = \b[14]  & ~new_n26801_;
  assign new_n26984_ = ~new_n26799_ & new_n26983_;
  assign new_n26985_ = ~new_n26803_ & ~new_n26984_;
  assign new_n26986_ = ~new_n26982_ & new_n26985_;
  assign new_n26987_ = ~new_n26803_ & ~new_n26986_;
  assign new_n26988_ = \b[15]  & ~new_n26792_;
  assign new_n26989_ = ~new_n26790_ & new_n26988_;
  assign new_n26990_ = ~new_n26794_ & ~new_n26989_;
  assign new_n26991_ = ~new_n26987_ & new_n26990_;
  assign new_n26992_ = ~new_n26794_ & ~new_n26991_;
  assign new_n26993_ = \b[16]  & ~new_n26783_;
  assign new_n26994_ = ~new_n26781_ & new_n26993_;
  assign new_n26995_ = ~new_n26785_ & ~new_n26994_;
  assign new_n26996_ = ~new_n26992_ & new_n26995_;
  assign new_n26997_ = ~new_n26785_ & ~new_n26996_;
  assign new_n26998_ = \b[17]  & ~new_n26774_;
  assign new_n26999_ = ~new_n26772_ & new_n26998_;
  assign new_n27000_ = ~new_n26776_ & ~new_n26999_;
  assign new_n27001_ = ~new_n26997_ & new_n27000_;
  assign new_n27002_ = ~new_n26776_ & ~new_n27001_;
  assign new_n27003_ = \b[18]  & ~new_n26765_;
  assign new_n27004_ = ~new_n26763_ & new_n27003_;
  assign new_n27005_ = ~new_n26767_ & ~new_n27004_;
  assign new_n27006_ = ~new_n27002_ & new_n27005_;
  assign new_n27007_ = ~new_n26767_ & ~new_n27006_;
  assign new_n27008_ = \b[19]  & ~new_n26756_;
  assign new_n27009_ = ~new_n26754_ & new_n27008_;
  assign new_n27010_ = ~new_n26758_ & ~new_n27009_;
  assign new_n27011_ = ~new_n27007_ & new_n27010_;
  assign new_n27012_ = ~new_n26758_ & ~new_n27011_;
  assign new_n27013_ = \b[20]  & ~new_n26747_;
  assign new_n27014_ = ~new_n26745_ & new_n27013_;
  assign new_n27015_ = ~new_n26749_ & ~new_n27014_;
  assign new_n27016_ = ~new_n27012_ & new_n27015_;
  assign new_n27017_ = ~new_n26749_ & ~new_n27016_;
  assign new_n27018_ = \b[21]  & ~new_n26738_;
  assign new_n27019_ = ~new_n26736_ & new_n27018_;
  assign new_n27020_ = ~new_n26740_ & ~new_n27019_;
  assign new_n27021_ = ~new_n27017_ & new_n27020_;
  assign new_n27022_ = ~new_n26740_ & ~new_n27021_;
  assign new_n27023_ = \b[22]  & ~new_n26729_;
  assign new_n27024_ = ~new_n26727_ & new_n27023_;
  assign new_n27025_ = ~new_n26731_ & ~new_n27024_;
  assign new_n27026_ = ~new_n27022_ & new_n27025_;
  assign new_n27027_ = ~new_n26731_ & ~new_n27026_;
  assign new_n27028_ = \b[23]  & ~new_n26720_;
  assign new_n27029_ = ~new_n26718_ & new_n27028_;
  assign new_n27030_ = ~new_n26722_ & ~new_n27029_;
  assign new_n27031_ = ~new_n27027_ & new_n27030_;
  assign new_n27032_ = ~new_n26722_ & ~new_n27031_;
  assign new_n27033_ = \b[24]  & ~new_n26711_;
  assign new_n27034_ = ~new_n26709_ & new_n27033_;
  assign new_n27035_ = ~new_n26713_ & ~new_n27034_;
  assign new_n27036_ = ~new_n27032_ & new_n27035_;
  assign new_n27037_ = ~new_n26713_ & ~new_n27036_;
  assign new_n27038_ = \b[25]  & ~new_n26702_;
  assign new_n27039_ = ~new_n26700_ & new_n27038_;
  assign new_n27040_ = ~new_n26704_ & ~new_n27039_;
  assign new_n27041_ = ~new_n27037_ & new_n27040_;
  assign new_n27042_ = ~new_n26704_ & ~new_n27041_;
  assign new_n27043_ = \b[26]  & ~new_n26693_;
  assign new_n27044_ = ~new_n26691_ & new_n27043_;
  assign new_n27045_ = ~new_n26695_ & ~new_n27044_;
  assign new_n27046_ = ~new_n27042_ & new_n27045_;
  assign new_n27047_ = ~new_n26695_ & ~new_n27046_;
  assign new_n27048_ = \b[27]  & ~new_n26684_;
  assign new_n27049_ = ~new_n26682_ & new_n27048_;
  assign new_n27050_ = ~new_n26686_ & ~new_n27049_;
  assign new_n27051_ = ~new_n27047_ & new_n27050_;
  assign new_n27052_ = ~new_n26686_ & ~new_n27051_;
  assign new_n27053_ = \b[28]  & ~new_n26675_;
  assign new_n27054_ = ~new_n26673_ & new_n27053_;
  assign new_n27055_ = ~new_n26677_ & ~new_n27054_;
  assign new_n27056_ = ~new_n27052_ & new_n27055_;
  assign new_n27057_ = ~new_n26677_ & ~new_n27056_;
  assign new_n27058_ = \b[29]  & ~new_n26666_;
  assign new_n27059_ = ~new_n26664_ & new_n27058_;
  assign new_n27060_ = ~new_n26668_ & ~new_n27059_;
  assign new_n27061_ = ~new_n27057_ & new_n27060_;
  assign new_n27062_ = ~new_n26668_ & ~new_n27061_;
  assign new_n27063_ = \b[30]  & ~new_n26657_;
  assign new_n27064_ = ~new_n26655_ & new_n27063_;
  assign new_n27065_ = ~new_n26659_ & ~new_n27064_;
  assign new_n27066_ = ~new_n27062_ & new_n27065_;
  assign new_n27067_ = ~new_n26659_ & ~new_n27066_;
  assign new_n27068_ = \b[31]  & ~new_n26648_;
  assign new_n27069_ = ~new_n26646_ & new_n27068_;
  assign new_n27070_ = ~new_n26650_ & ~new_n27069_;
  assign new_n27071_ = ~new_n27067_ & new_n27070_;
  assign new_n27072_ = ~new_n26650_ & ~new_n27071_;
  assign new_n27073_ = \b[32]  & ~new_n26639_;
  assign new_n27074_ = ~new_n26637_ & new_n27073_;
  assign new_n27075_ = ~new_n26641_ & ~new_n27074_;
  assign new_n27076_ = ~new_n27072_ & new_n27075_;
  assign new_n27077_ = ~new_n26641_ & ~new_n27076_;
  assign new_n27078_ = \b[33]  & ~new_n26630_;
  assign new_n27079_ = ~new_n26628_ & new_n27078_;
  assign new_n27080_ = ~new_n26632_ & ~new_n27079_;
  assign new_n27081_ = ~new_n27077_ & new_n27080_;
  assign new_n27082_ = ~new_n26632_ & ~new_n27081_;
  assign new_n27083_ = \b[34]  & ~new_n26621_;
  assign new_n27084_ = ~new_n26619_ & new_n27083_;
  assign new_n27085_ = ~new_n26623_ & ~new_n27084_;
  assign new_n27086_ = ~new_n27082_ & new_n27085_;
  assign new_n27087_ = ~new_n26623_ & ~new_n27086_;
  assign new_n27088_ = \b[35]  & ~new_n26612_;
  assign new_n27089_ = ~new_n26610_ & new_n27088_;
  assign new_n27090_ = ~new_n26614_ & ~new_n27089_;
  assign new_n27091_ = ~new_n27087_ & new_n27090_;
  assign new_n27092_ = ~new_n26614_ & ~new_n27091_;
  assign new_n27093_ = \b[36]  & ~new_n26603_;
  assign new_n27094_ = ~new_n26601_ & new_n27093_;
  assign new_n27095_ = ~new_n26605_ & ~new_n27094_;
  assign new_n27096_ = ~new_n27092_ & new_n27095_;
  assign new_n27097_ = ~new_n26605_ & ~new_n27096_;
  assign new_n27098_ = \b[37]  & ~new_n26594_;
  assign new_n27099_ = ~new_n26592_ & new_n27098_;
  assign new_n27100_ = ~new_n26596_ & ~new_n27099_;
  assign new_n27101_ = ~new_n27097_ & new_n27100_;
  assign new_n27102_ = ~new_n26596_ & ~new_n27101_;
  assign new_n27103_ = \b[38]  & ~new_n26585_;
  assign new_n27104_ = ~new_n26583_ & new_n27103_;
  assign new_n27105_ = ~new_n26587_ & ~new_n27104_;
  assign new_n27106_ = ~new_n27102_ & new_n27105_;
  assign new_n27107_ = ~new_n26587_ & ~new_n27106_;
  assign new_n27108_ = \b[39]  & ~new_n26576_;
  assign new_n27109_ = ~new_n26574_ & new_n27108_;
  assign new_n27110_ = ~new_n26578_ & ~new_n27109_;
  assign new_n27111_ = ~new_n27107_ & new_n27110_;
  assign new_n27112_ = ~new_n26578_ & ~new_n27111_;
  assign new_n27113_ = \b[40]  & ~new_n26567_;
  assign new_n27114_ = ~new_n26565_ & new_n27113_;
  assign new_n27115_ = ~new_n26569_ & ~new_n27114_;
  assign new_n27116_ = ~new_n27112_ & new_n27115_;
  assign new_n27117_ = ~new_n26569_ & ~new_n27116_;
  assign new_n27118_ = \b[41]  & ~new_n26558_;
  assign new_n27119_ = ~new_n26556_ & new_n27118_;
  assign new_n27120_ = ~new_n26560_ & ~new_n27119_;
  assign new_n27121_ = ~new_n27117_ & new_n27120_;
  assign new_n27122_ = ~new_n26560_ & ~new_n27121_;
  assign new_n27123_ = \b[42]  & ~new_n26549_;
  assign new_n27124_ = ~new_n26547_ & new_n27123_;
  assign new_n27125_ = ~new_n26551_ & ~new_n27124_;
  assign new_n27126_ = ~new_n27122_ & new_n27125_;
  assign new_n27127_ = ~new_n26551_ & ~new_n27126_;
  assign new_n27128_ = \b[43]  & ~new_n26540_;
  assign new_n27129_ = ~new_n26538_ & new_n27128_;
  assign new_n27130_ = ~new_n26542_ & ~new_n27129_;
  assign new_n27131_ = ~new_n27127_ & new_n27130_;
  assign new_n27132_ = ~new_n26542_ & ~new_n27131_;
  assign new_n27133_ = \b[44]  & ~new_n26531_;
  assign new_n27134_ = ~new_n26529_ & new_n27133_;
  assign new_n27135_ = ~new_n26533_ & ~new_n27134_;
  assign new_n27136_ = ~new_n27132_ & new_n27135_;
  assign new_n27137_ = ~new_n26533_ & ~new_n27136_;
  assign new_n27138_ = \b[45]  & ~new_n26522_;
  assign new_n27139_ = ~new_n26520_ & new_n27138_;
  assign new_n27140_ = ~new_n26524_ & ~new_n27139_;
  assign new_n27141_ = ~new_n27137_ & new_n27140_;
  assign new_n27142_ = ~new_n26524_ & ~new_n27141_;
  assign new_n27143_ = \b[46]  & ~new_n26513_;
  assign new_n27144_ = ~new_n26511_ & new_n27143_;
  assign new_n27145_ = ~new_n26515_ & ~new_n27144_;
  assign new_n27146_ = ~new_n27142_ & new_n27145_;
  assign new_n27147_ = ~new_n26515_ & ~new_n27146_;
  assign new_n27148_ = \b[47]  & ~new_n26504_;
  assign new_n27149_ = ~new_n26502_ & new_n27148_;
  assign new_n27150_ = ~new_n26506_ & ~new_n27149_;
  assign new_n27151_ = ~new_n27147_ & new_n27150_;
  assign new_n27152_ = ~new_n26506_ & ~new_n27151_;
  assign new_n27153_ = \b[48]  & ~new_n26495_;
  assign new_n27154_ = ~new_n26493_ & new_n27153_;
  assign new_n27155_ = ~new_n26497_ & ~new_n27154_;
  assign new_n27156_ = ~new_n27152_ & new_n27155_;
  assign new_n27157_ = ~new_n26497_ & ~new_n27156_;
  assign new_n27158_ = \b[49]  & ~new_n26486_;
  assign new_n27159_ = ~new_n26484_ & new_n27158_;
  assign new_n27160_ = ~new_n26488_ & ~new_n27159_;
  assign new_n27161_ = ~new_n27157_ & new_n27160_;
  assign new_n27162_ = ~new_n26488_ & ~new_n27161_;
  assign new_n27163_ = \b[50]  & ~new_n26477_;
  assign new_n27164_ = ~new_n26475_ & new_n27163_;
  assign new_n27165_ = ~new_n26479_ & ~new_n27164_;
  assign new_n27166_ = ~new_n27162_ & new_n27165_;
  assign new_n27167_ = ~new_n26479_ & ~new_n27166_;
  assign new_n27168_ = \b[51]  & ~new_n26468_;
  assign new_n27169_ = ~new_n26466_ & new_n27168_;
  assign new_n27170_ = ~new_n26470_ & ~new_n27169_;
  assign new_n27171_ = ~new_n27167_ & new_n27170_;
  assign new_n27172_ = ~new_n26470_ & ~new_n27171_;
  assign new_n27173_ = \b[52]  & ~new_n26459_;
  assign new_n27174_ = ~new_n26457_ & new_n27173_;
  assign new_n27175_ = ~new_n26461_ & ~new_n27174_;
  assign new_n27176_ = ~new_n27172_ & new_n27175_;
  assign new_n27177_ = ~new_n26461_ & ~new_n27176_;
  assign new_n27178_ = \b[53]  & ~new_n26450_;
  assign new_n27179_ = ~new_n26448_ & new_n27178_;
  assign new_n27180_ = ~new_n26452_ & ~new_n27179_;
  assign new_n27181_ = ~new_n27177_ & new_n27180_;
  assign new_n27182_ = ~new_n26452_ & ~new_n27181_;
  assign new_n27183_ = \b[54]  & ~new_n26441_;
  assign new_n27184_ = ~new_n26439_ & new_n27183_;
  assign new_n27185_ = ~new_n26443_ & ~new_n27184_;
  assign new_n27186_ = ~new_n27182_ & new_n27185_;
  assign new_n27187_ = ~new_n26443_ & ~new_n27186_;
  assign new_n27188_ = \b[55]  & ~new_n26432_;
  assign new_n27189_ = ~new_n26430_ & new_n27188_;
  assign new_n27190_ = ~new_n26434_ & ~new_n27189_;
  assign new_n27191_ = ~new_n27187_ & new_n27190_;
  assign new_n27192_ = ~new_n26434_ & ~new_n27191_;
  assign new_n27193_ = \b[56]  & ~new_n26423_;
  assign new_n27194_ = ~new_n26421_ & new_n27193_;
  assign new_n27195_ = ~new_n26425_ & ~new_n27194_;
  assign new_n27196_ = ~new_n27192_ & new_n27195_;
  assign new_n27197_ = ~new_n26425_ & ~new_n27196_;
  assign new_n27198_ = \b[57]  & ~new_n26414_;
  assign new_n27199_ = ~new_n26412_ & new_n27198_;
  assign new_n27200_ = ~new_n26416_ & ~new_n27199_;
  assign new_n27201_ = ~new_n27197_ & new_n27200_;
  assign new_n27202_ = ~new_n26416_ & ~new_n27201_;
  assign new_n27203_ = \b[58]  & ~new_n26405_;
  assign new_n27204_ = ~new_n26403_ & new_n27203_;
  assign new_n27205_ = ~new_n26407_ & ~new_n27204_;
  assign new_n27206_ = ~new_n27202_ & new_n27205_;
  assign new_n27207_ = ~new_n26407_ & ~new_n27206_;
  assign new_n27208_ = \b[59]  & ~new_n26396_;
  assign new_n27209_ = ~new_n26394_ & new_n27208_;
  assign new_n27210_ = ~new_n26398_ & ~new_n27209_;
  assign new_n27211_ = ~new_n27207_ & new_n27210_;
  assign new_n27212_ = ~new_n26398_ & ~new_n27211_;
  assign new_n27213_ = \b[60]  & ~new_n26387_;
  assign new_n27214_ = ~new_n26385_ & new_n27213_;
  assign new_n27215_ = ~new_n26389_ & ~new_n27214_;
  assign new_n27216_ = ~new_n27212_ & new_n27215_;
  assign new_n27217_ = ~new_n26389_ & ~new_n27216_;
  assign new_n27218_ = ~new_n25548_ & ~new_n26375_;
  assign new_n27219_ = ~new_n26373_ & new_n27218_;
  assign new_n27220_ = ~new_n26361_ & new_n27219_;
  assign new_n27221_ = ~new_n26373_ & ~new_n26375_;
  assign new_n27222_ = ~new_n26362_ & ~new_n27221_;
  assign new_n27223_ = ~new_n27220_ & ~new_n27222_;
  assign new_n27224_ = \quotient[3]  & ~new_n27223_;
  assign new_n27225_ = ~new_n26372_ & ~new_n26379_;
  assign new_n27226_ = ~new_n26378_ & new_n27225_;
  assign new_n27227_ = ~new_n27224_ & ~new_n27226_;
  assign new_n27228_ = ~\b[61]  & ~new_n27227_;
  assign new_n27229_ = \b[61]  & ~new_n27226_;
  assign new_n27230_ = ~new_n27224_ & new_n27229_;
  assign new_n27231_ = new_n279_ & ~new_n27230_;
  assign new_n27232_ = ~new_n27228_ & new_n27231_;
  assign new_n27233_ = ~new_n27217_ & new_n27232_;
  assign new_n27234_ = new_n403_ & ~new_n27227_;
  assign \quotient[2]  = new_n27233_ | new_n27234_;
  assign new_n27236_ = ~new_n26398_ & new_n27215_;
  assign new_n27237_ = ~new_n27211_ & new_n27236_;
  assign new_n27238_ = ~new_n27212_ & ~new_n27215_;
  assign new_n27239_ = ~new_n27237_ & ~new_n27238_;
  assign new_n27240_ = \quotient[2]  & ~new_n27239_;
  assign new_n27241_ = ~new_n26388_ & ~new_n27234_;
  assign new_n27242_ = ~new_n27233_ & new_n27241_;
  assign new_n27243_ = ~new_n27240_ & ~new_n27242_;
  assign new_n27244_ = ~\b[61]  & ~new_n27243_;
  assign new_n27245_ = ~new_n26407_ & new_n27210_;
  assign new_n27246_ = ~new_n27206_ & new_n27245_;
  assign new_n27247_ = ~new_n27207_ & ~new_n27210_;
  assign new_n27248_ = ~new_n27246_ & ~new_n27247_;
  assign new_n27249_ = \quotient[2]  & ~new_n27248_;
  assign new_n27250_ = ~new_n26397_ & ~new_n27234_;
  assign new_n27251_ = ~new_n27233_ & new_n27250_;
  assign new_n27252_ = ~new_n27249_ & ~new_n27251_;
  assign new_n27253_ = ~\b[60]  & ~new_n27252_;
  assign new_n27254_ = ~new_n26416_ & new_n27205_;
  assign new_n27255_ = ~new_n27201_ & new_n27254_;
  assign new_n27256_ = ~new_n27202_ & ~new_n27205_;
  assign new_n27257_ = ~new_n27255_ & ~new_n27256_;
  assign new_n27258_ = \quotient[2]  & ~new_n27257_;
  assign new_n27259_ = ~new_n26406_ & ~new_n27234_;
  assign new_n27260_ = ~new_n27233_ & new_n27259_;
  assign new_n27261_ = ~new_n27258_ & ~new_n27260_;
  assign new_n27262_ = ~\b[59]  & ~new_n27261_;
  assign new_n27263_ = ~new_n26425_ & new_n27200_;
  assign new_n27264_ = ~new_n27196_ & new_n27263_;
  assign new_n27265_ = ~new_n27197_ & ~new_n27200_;
  assign new_n27266_ = ~new_n27264_ & ~new_n27265_;
  assign new_n27267_ = \quotient[2]  & ~new_n27266_;
  assign new_n27268_ = ~new_n26415_ & ~new_n27234_;
  assign new_n27269_ = ~new_n27233_ & new_n27268_;
  assign new_n27270_ = ~new_n27267_ & ~new_n27269_;
  assign new_n27271_ = ~\b[58]  & ~new_n27270_;
  assign new_n27272_ = ~new_n26434_ & new_n27195_;
  assign new_n27273_ = ~new_n27191_ & new_n27272_;
  assign new_n27274_ = ~new_n27192_ & ~new_n27195_;
  assign new_n27275_ = ~new_n27273_ & ~new_n27274_;
  assign new_n27276_ = \quotient[2]  & ~new_n27275_;
  assign new_n27277_ = ~new_n26424_ & ~new_n27234_;
  assign new_n27278_ = ~new_n27233_ & new_n27277_;
  assign new_n27279_ = ~new_n27276_ & ~new_n27278_;
  assign new_n27280_ = ~\b[57]  & ~new_n27279_;
  assign new_n27281_ = ~new_n26443_ & new_n27190_;
  assign new_n27282_ = ~new_n27186_ & new_n27281_;
  assign new_n27283_ = ~new_n27187_ & ~new_n27190_;
  assign new_n27284_ = ~new_n27282_ & ~new_n27283_;
  assign new_n27285_ = \quotient[2]  & ~new_n27284_;
  assign new_n27286_ = ~new_n26433_ & ~new_n27234_;
  assign new_n27287_ = ~new_n27233_ & new_n27286_;
  assign new_n27288_ = ~new_n27285_ & ~new_n27287_;
  assign new_n27289_ = ~\b[56]  & ~new_n27288_;
  assign new_n27290_ = ~new_n26452_ & new_n27185_;
  assign new_n27291_ = ~new_n27181_ & new_n27290_;
  assign new_n27292_ = ~new_n27182_ & ~new_n27185_;
  assign new_n27293_ = ~new_n27291_ & ~new_n27292_;
  assign new_n27294_ = \quotient[2]  & ~new_n27293_;
  assign new_n27295_ = ~new_n26442_ & ~new_n27234_;
  assign new_n27296_ = ~new_n27233_ & new_n27295_;
  assign new_n27297_ = ~new_n27294_ & ~new_n27296_;
  assign new_n27298_ = ~\b[55]  & ~new_n27297_;
  assign new_n27299_ = ~new_n26461_ & new_n27180_;
  assign new_n27300_ = ~new_n27176_ & new_n27299_;
  assign new_n27301_ = ~new_n27177_ & ~new_n27180_;
  assign new_n27302_ = ~new_n27300_ & ~new_n27301_;
  assign new_n27303_ = \quotient[2]  & ~new_n27302_;
  assign new_n27304_ = ~new_n26451_ & ~new_n27234_;
  assign new_n27305_ = ~new_n27233_ & new_n27304_;
  assign new_n27306_ = ~new_n27303_ & ~new_n27305_;
  assign new_n27307_ = ~\b[54]  & ~new_n27306_;
  assign new_n27308_ = ~new_n26470_ & new_n27175_;
  assign new_n27309_ = ~new_n27171_ & new_n27308_;
  assign new_n27310_ = ~new_n27172_ & ~new_n27175_;
  assign new_n27311_ = ~new_n27309_ & ~new_n27310_;
  assign new_n27312_ = \quotient[2]  & ~new_n27311_;
  assign new_n27313_ = ~new_n26460_ & ~new_n27234_;
  assign new_n27314_ = ~new_n27233_ & new_n27313_;
  assign new_n27315_ = ~new_n27312_ & ~new_n27314_;
  assign new_n27316_ = ~\b[53]  & ~new_n27315_;
  assign new_n27317_ = ~new_n26479_ & new_n27170_;
  assign new_n27318_ = ~new_n27166_ & new_n27317_;
  assign new_n27319_ = ~new_n27167_ & ~new_n27170_;
  assign new_n27320_ = ~new_n27318_ & ~new_n27319_;
  assign new_n27321_ = \quotient[2]  & ~new_n27320_;
  assign new_n27322_ = ~new_n26469_ & ~new_n27234_;
  assign new_n27323_ = ~new_n27233_ & new_n27322_;
  assign new_n27324_ = ~new_n27321_ & ~new_n27323_;
  assign new_n27325_ = ~\b[52]  & ~new_n27324_;
  assign new_n27326_ = ~new_n26488_ & new_n27165_;
  assign new_n27327_ = ~new_n27161_ & new_n27326_;
  assign new_n27328_ = ~new_n27162_ & ~new_n27165_;
  assign new_n27329_ = ~new_n27327_ & ~new_n27328_;
  assign new_n27330_ = \quotient[2]  & ~new_n27329_;
  assign new_n27331_ = ~new_n26478_ & ~new_n27234_;
  assign new_n27332_ = ~new_n27233_ & new_n27331_;
  assign new_n27333_ = ~new_n27330_ & ~new_n27332_;
  assign new_n27334_ = ~\b[51]  & ~new_n27333_;
  assign new_n27335_ = ~new_n26497_ & new_n27160_;
  assign new_n27336_ = ~new_n27156_ & new_n27335_;
  assign new_n27337_ = ~new_n27157_ & ~new_n27160_;
  assign new_n27338_ = ~new_n27336_ & ~new_n27337_;
  assign new_n27339_ = \quotient[2]  & ~new_n27338_;
  assign new_n27340_ = ~new_n26487_ & ~new_n27234_;
  assign new_n27341_ = ~new_n27233_ & new_n27340_;
  assign new_n27342_ = ~new_n27339_ & ~new_n27341_;
  assign new_n27343_ = ~\b[50]  & ~new_n27342_;
  assign new_n27344_ = ~new_n26506_ & new_n27155_;
  assign new_n27345_ = ~new_n27151_ & new_n27344_;
  assign new_n27346_ = ~new_n27152_ & ~new_n27155_;
  assign new_n27347_ = ~new_n27345_ & ~new_n27346_;
  assign new_n27348_ = \quotient[2]  & ~new_n27347_;
  assign new_n27349_ = ~new_n26496_ & ~new_n27234_;
  assign new_n27350_ = ~new_n27233_ & new_n27349_;
  assign new_n27351_ = ~new_n27348_ & ~new_n27350_;
  assign new_n27352_ = ~\b[49]  & ~new_n27351_;
  assign new_n27353_ = ~new_n26515_ & new_n27150_;
  assign new_n27354_ = ~new_n27146_ & new_n27353_;
  assign new_n27355_ = ~new_n27147_ & ~new_n27150_;
  assign new_n27356_ = ~new_n27354_ & ~new_n27355_;
  assign new_n27357_ = \quotient[2]  & ~new_n27356_;
  assign new_n27358_ = ~new_n26505_ & ~new_n27234_;
  assign new_n27359_ = ~new_n27233_ & new_n27358_;
  assign new_n27360_ = ~new_n27357_ & ~new_n27359_;
  assign new_n27361_ = ~\b[48]  & ~new_n27360_;
  assign new_n27362_ = ~new_n26524_ & new_n27145_;
  assign new_n27363_ = ~new_n27141_ & new_n27362_;
  assign new_n27364_ = ~new_n27142_ & ~new_n27145_;
  assign new_n27365_ = ~new_n27363_ & ~new_n27364_;
  assign new_n27366_ = \quotient[2]  & ~new_n27365_;
  assign new_n27367_ = ~new_n26514_ & ~new_n27234_;
  assign new_n27368_ = ~new_n27233_ & new_n27367_;
  assign new_n27369_ = ~new_n27366_ & ~new_n27368_;
  assign new_n27370_ = ~\b[47]  & ~new_n27369_;
  assign new_n27371_ = ~new_n26533_ & new_n27140_;
  assign new_n27372_ = ~new_n27136_ & new_n27371_;
  assign new_n27373_ = ~new_n27137_ & ~new_n27140_;
  assign new_n27374_ = ~new_n27372_ & ~new_n27373_;
  assign new_n27375_ = \quotient[2]  & ~new_n27374_;
  assign new_n27376_ = ~new_n26523_ & ~new_n27234_;
  assign new_n27377_ = ~new_n27233_ & new_n27376_;
  assign new_n27378_ = ~new_n27375_ & ~new_n27377_;
  assign new_n27379_ = ~\b[46]  & ~new_n27378_;
  assign new_n27380_ = ~new_n26542_ & new_n27135_;
  assign new_n27381_ = ~new_n27131_ & new_n27380_;
  assign new_n27382_ = ~new_n27132_ & ~new_n27135_;
  assign new_n27383_ = ~new_n27381_ & ~new_n27382_;
  assign new_n27384_ = \quotient[2]  & ~new_n27383_;
  assign new_n27385_ = ~new_n26532_ & ~new_n27234_;
  assign new_n27386_ = ~new_n27233_ & new_n27385_;
  assign new_n27387_ = ~new_n27384_ & ~new_n27386_;
  assign new_n27388_ = ~\b[45]  & ~new_n27387_;
  assign new_n27389_ = ~new_n26551_ & new_n27130_;
  assign new_n27390_ = ~new_n27126_ & new_n27389_;
  assign new_n27391_ = ~new_n27127_ & ~new_n27130_;
  assign new_n27392_ = ~new_n27390_ & ~new_n27391_;
  assign new_n27393_ = \quotient[2]  & ~new_n27392_;
  assign new_n27394_ = ~new_n26541_ & ~new_n27234_;
  assign new_n27395_ = ~new_n27233_ & new_n27394_;
  assign new_n27396_ = ~new_n27393_ & ~new_n27395_;
  assign new_n27397_ = ~\b[44]  & ~new_n27396_;
  assign new_n27398_ = ~new_n26560_ & new_n27125_;
  assign new_n27399_ = ~new_n27121_ & new_n27398_;
  assign new_n27400_ = ~new_n27122_ & ~new_n27125_;
  assign new_n27401_ = ~new_n27399_ & ~new_n27400_;
  assign new_n27402_ = \quotient[2]  & ~new_n27401_;
  assign new_n27403_ = ~new_n26550_ & ~new_n27234_;
  assign new_n27404_ = ~new_n27233_ & new_n27403_;
  assign new_n27405_ = ~new_n27402_ & ~new_n27404_;
  assign new_n27406_ = ~\b[43]  & ~new_n27405_;
  assign new_n27407_ = ~new_n26569_ & new_n27120_;
  assign new_n27408_ = ~new_n27116_ & new_n27407_;
  assign new_n27409_ = ~new_n27117_ & ~new_n27120_;
  assign new_n27410_ = ~new_n27408_ & ~new_n27409_;
  assign new_n27411_ = \quotient[2]  & ~new_n27410_;
  assign new_n27412_ = ~new_n26559_ & ~new_n27234_;
  assign new_n27413_ = ~new_n27233_ & new_n27412_;
  assign new_n27414_ = ~new_n27411_ & ~new_n27413_;
  assign new_n27415_ = ~\b[42]  & ~new_n27414_;
  assign new_n27416_ = ~new_n26578_ & new_n27115_;
  assign new_n27417_ = ~new_n27111_ & new_n27416_;
  assign new_n27418_ = ~new_n27112_ & ~new_n27115_;
  assign new_n27419_ = ~new_n27417_ & ~new_n27418_;
  assign new_n27420_ = \quotient[2]  & ~new_n27419_;
  assign new_n27421_ = ~new_n26568_ & ~new_n27234_;
  assign new_n27422_ = ~new_n27233_ & new_n27421_;
  assign new_n27423_ = ~new_n27420_ & ~new_n27422_;
  assign new_n27424_ = ~\b[41]  & ~new_n27423_;
  assign new_n27425_ = ~new_n26587_ & new_n27110_;
  assign new_n27426_ = ~new_n27106_ & new_n27425_;
  assign new_n27427_ = ~new_n27107_ & ~new_n27110_;
  assign new_n27428_ = ~new_n27426_ & ~new_n27427_;
  assign new_n27429_ = \quotient[2]  & ~new_n27428_;
  assign new_n27430_ = ~new_n26577_ & ~new_n27234_;
  assign new_n27431_ = ~new_n27233_ & new_n27430_;
  assign new_n27432_ = ~new_n27429_ & ~new_n27431_;
  assign new_n27433_ = ~\b[40]  & ~new_n27432_;
  assign new_n27434_ = ~new_n26596_ & new_n27105_;
  assign new_n27435_ = ~new_n27101_ & new_n27434_;
  assign new_n27436_ = ~new_n27102_ & ~new_n27105_;
  assign new_n27437_ = ~new_n27435_ & ~new_n27436_;
  assign new_n27438_ = \quotient[2]  & ~new_n27437_;
  assign new_n27439_ = ~new_n26586_ & ~new_n27234_;
  assign new_n27440_ = ~new_n27233_ & new_n27439_;
  assign new_n27441_ = ~new_n27438_ & ~new_n27440_;
  assign new_n27442_ = ~\b[39]  & ~new_n27441_;
  assign new_n27443_ = ~new_n26605_ & new_n27100_;
  assign new_n27444_ = ~new_n27096_ & new_n27443_;
  assign new_n27445_ = ~new_n27097_ & ~new_n27100_;
  assign new_n27446_ = ~new_n27444_ & ~new_n27445_;
  assign new_n27447_ = \quotient[2]  & ~new_n27446_;
  assign new_n27448_ = ~new_n26595_ & ~new_n27234_;
  assign new_n27449_ = ~new_n27233_ & new_n27448_;
  assign new_n27450_ = ~new_n27447_ & ~new_n27449_;
  assign new_n27451_ = ~\b[38]  & ~new_n27450_;
  assign new_n27452_ = ~new_n26614_ & new_n27095_;
  assign new_n27453_ = ~new_n27091_ & new_n27452_;
  assign new_n27454_ = ~new_n27092_ & ~new_n27095_;
  assign new_n27455_ = ~new_n27453_ & ~new_n27454_;
  assign new_n27456_ = \quotient[2]  & ~new_n27455_;
  assign new_n27457_ = ~new_n26604_ & ~new_n27234_;
  assign new_n27458_ = ~new_n27233_ & new_n27457_;
  assign new_n27459_ = ~new_n27456_ & ~new_n27458_;
  assign new_n27460_ = ~\b[37]  & ~new_n27459_;
  assign new_n27461_ = ~new_n26623_ & new_n27090_;
  assign new_n27462_ = ~new_n27086_ & new_n27461_;
  assign new_n27463_ = ~new_n27087_ & ~new_n27090_;
  assign new_n27464_ = ~new_n27462_ & ~new_n27463_;
  assign new_n27465_ = \quotient[2]  & ~new_n27464_;
  assign new_n27466_ = ~new_n26613_ & ~new_n27234_;
  assign new_n27467_ = ~new_n27233_ & new_n27466_;
  assign new_n27468_ = ~new_n27465_ & ~new_n27467_;
  assign new_n27469_ = ~\b[36]  & ~new_n27468_;
  assign new_n27470_ = ~new_n26632_ & new_n27085_;
  assign new_n27471_ = ~new_n27081_ & new_n27470_;
  assign new_n27472_ = ~new_n27082_ & ~new_n27085_;
  assign new_n27473_ = ~new_n27471_ & ~new_n27472_;
  assign new_n27474_ = \quotient[2]  & ~new_n27473_;
  assign new_n27475_ = ~new_n26622_ & ~new_n27234_;
  assign new_n27476_ = ~new_n27233_ & new_n27475_;
  assign new_n27477_ = ~new_n27474_ & ~new_n27476_;
  assign new_n27478_ = ~\b[35]  & ~new_n27477_;
  assign new_n27479_ = ~new_n26641_ & new_n27080_;
  assign new_n27480_ = ~new_n27076_ & new_n27479_;
  assign new_n27481_ = ~new_n27077_ & ~new_n27080_;
  assign new_n27482_ = ~new_n27480_ & ~new_n27481_;
  assign new_n27483_ = \quotient[2]  & ~new_n27482_;
  assign new_n27484_ = ~new_n26631_ & ~new_n27234_;
  assign new_n27485_ = ~new_n27233_ & new_n27484_;
  assign new_n27486_ = ~new_n27483_ & ~new_n27485_;
  assign new_n27487_ = ~\b[34]  & ~new_n27486_;
  assign new_n27488_ = ~new_n26650_ & new_n27075_;
  assign new_n27489_ = ~new_n27071_ & new_n27488_;
  assign new_n27490_ = ~new_n27072_ & ~new_n27075_;
  assign new_n27491_ = ~new_n27489_ & ~new_n27490_;
  assign new_n27492_ = \quotient[2]  & ~new_n27491_;
  assign new_n27493_ = ~new_n26640_ & ~new_n27234_;
  assign new_n27494_ = ~new_n27233_ & new_n27493_;
  assign new_n27495_ = ~new_n27492_ & ~new_n27494_;
  assign new_n27496_ = ~\b[33]  & ~new_n27495_;
  assign new_n27497_ = ~new_n26659_ & new_n27070_;
  assign new_n27498_ = ~new_n27066_ & new_n27497_;
  assign new_n27499_ = ~new_n27067_ & ~new_n27070_;
  assign new_n27500_ = ~new_n27498_ & ~new_n27499_;
  assign new_n27501_ = \quotient[2]  & ~new_n27500_;
  assign new_n27502_ = ~new_n26649_ & ~new_n27234_;
  assign new_n27503_ = ~new_n27233_ & new_n27502_;
  assign new_n27504_ = ~new_n27501_ & ~new_n27503_;
  assign new_n27505_ = ~\b[32]  & ~new_n27504_;
  assign new_n27506_ = ~new_n26668_ & new_n27065_;
  assign new_n27507_ = ~new_n27061_ & new_n27506_;
  assign new_n27508_ = ~new_n27062_ & ~new_n27065_;
  assign new_n27509_ = ~new_n27507_ & ~new_n27508_;
  assign new_n27510_ = \quotient[2]  & ~new_n27509_;
  assign new_n27511_ = ~new_n26658_ & ~new_n27234_;
  assign new_n27512_ = ~new_n27233_ & new_n27511_;
  assign new_n27513_ = ~new_n27510_ & ~new_n27512_;
  assign new_n27514_ = ~\b[31]  & ~new_n27513_;
  assign new_n27515_ = ~new_n26677_ & new_n27060_;
  assign new_n27516_ = ~new_n27056_ & new_n27515_;
  assign new_n27517_ = ~new_n27057_ & ~new_n27060_;
  assign new_n27518_ = ~new_n27516_ & ~new_n27517_;
  assign new_n27519_ = \quotient[2]  & ~new_n27518_;
  assign new_n27520_ = ~new_n26667_ & ~new_n27234_;
  assign new_n27521_ = ~new_n27233_ & new_n27520_;
  assign new_n27522_ = ~new_n27519_ & ~new_n27521_;
  assign new_n27523_ = ~\b[30]  & ~new_n27522_;
  assign new_n27524_ = ~new_n26686_ & new_n27055_;
  assign new_n27525_ = ~new_n27051_ & new_n27524_;
  assign new_n27526_ = ~new_n27052_ & ~new_n27055_;
  assign new_n27527_ = ~new_n27525_ & ~new_n27526_;
  assign new_n27528_ = \quotient[2]  & ~new_n27527_;
  assign new_n27529_ = ~new_n26676_ & ~new_n27234_;
  assign new_n27530_ = ~new_n27233_ & new_n27529_;
  assign new_n27531_ = ~new_n27528_ & ~new_n27530_;
  assign new_n27532_ = ~\b[29]  & ~new_n27531_;
  assign new_n27533_ = ~new_n26695_ & new_n27050_;
  assign new_n27534_ = ~new_n27046_ & new_n27533_;
  assign new_n27535_ = ~new_n27047_ & ~new_n27050_;
  assign new_n27536_ = ~new_n27534_ & ~new_n27535_;
  assign new_n27537_ = \quotient[2]  & ~new_n27536_;
  assign new_n27538_ = ~new_n26685_ & ~new_n27234_;
  assign new_n27539_ = ~new_n27233_ & new_n27538_;
  assign new_n27540_ = ~new_n27537_ & ~new_n27539_;
  assign new_n27541_ = ~\b[28]  & ~new_n27540_;
  assign new_n27542_ = ~new_n26704_ & new_n27045_;
  assign new_n27543_ = ~new_n27041_ & new_n27542_;
  assign new_n27544_ = ~new_n27042_ & ~new_n27045_;
  assign new_n27545_ = ~new_n27543_ & ~new_n27544_;
  assign new_n27546_ = \quotient[2]  & ~new_n27545_;
  assign new_n27547_ = ~new_n26694_ & ~new_n27234_;
  assign new_n27548_ = ~new_n27233_ & new_n27547_;
  assign new_n27549_ = ~new_n27546_ & ~new_n27548_;
  assign new_n27550_ = ~\b[27]  & ~new_n27549_;
  assign new_n27551_ = ~new_n26713_ & new_n27040_;
  assign new_n27552_ = ~new_n27036_ & new_n27551_;
  assign new_n27553_ = ~new_n27037_ & ~new_n27040_;
  assign new_n27554_ = ~new_n27552_ & ~new_n27553_;
  assign new_n27555_ = \quotient[2]  & ~new_n27554_;
  assign new_n27556_ = ~new_n26703_ & ~new_n27234_;
  assign new_n27557_ = ~new_n27233_ & new_n27556_;
  assign new_n27558_ = ~new_n27555_ & ~new_n27557_;
  assign new_n27559_ = ~\b[26]  & ~new_n27558_;
  assign new_n27560_ = ~new_n26722_ & new_n27035_;
  assign new_n27561_ = ~new_n27031_ & new_n27560_;
  assign new_n27562_ = ~new_n27032_ & ~new_n27035_;
  assign new_n27563_ = ~new_n27561_ & ~new_n27562_;
  assign new_n27564_ = \quotient[2]  & ~new_n27563_;
  assign new_n27565_ = ~new_n26712_ & ~new_n27234_;
  assign new_n27566_ = ~new_n27233_ & new_n27565_;
  assign new_n27567_ = ~new_n27564_ & ~new_n27566_;
  assign new_n27568_ = ~\b[25]  & ~new_n27567_;
  assign new_n27569_ = ~new_n26731_ & new_n27030_;
  assign new_n27570_ = ~new_n27026_ & new_n27569_;
  assign new_n27571_ = ~new_n27027_ & ~new_n27030_;
  assign new_n27572_ = ~new_n27570_ & ~new_n27571_;
  assign new_n27573_ = \quotient[2]  & ~new_n27572_;
  assign new_n27574_ = ~new_n26721_ & ~new_n27234_;
  assign new_n27575_ = ~new_n27233_ & new_n27574_;
  assign new_n27576_ = ~new_n27573_ & ~new_n27575_;
  assign new_n27577_ = ~\b[24]  & ~new_n27576_;
  assign new_n27578_ = ~new_n26740_ & new_n27025_;
  assign new_n27579_ = ~new_n27021_ & new_n27578_;
  assign new_n27580_ = ~new_n27022_ & ~new_n27025_;
  assign new_n27581_ = ~new_n27579_ & ~new_n27580_;
  assign new_n27582_ = \quotient[2]  & ~new_n27581_;
  assign new_n27583_ = ~new_n26730_ & ~new_n27234_;
  assign new_n27584_ = ~new_n27233_ & new_n27583_;
  assign new_n27585_ = ~new_n27582_ & ~new_n27584_;
  assign new_n27586_ = ~\b[23]  & ~new_n27585_;
  assign new_n27587_ = ~new_n26749_ & new_n27020_;
  assign new_n27588_ = ~new_n27016_ & new_n27587_;
  assign new_n27589_ = ~new_n27017_ & ~new_n27020_;
  assign new_n27590_ = ~new_n27588_ & ~new_n27589_;
  assign new_n27591_ = \quotient[2]  & ~new_n27590_;
  assign new_n27592_ = ~new_n26739_ & ~new_n27234_;
  assign new_n27593_ = ~new_n27233_ & new_n27592_;
  assign new_n27594_ = ~new_n27591_ & ~new_n27593_;
  assign new_n27595_ = ~\b[22]  & ~new_n27594_;
  assign new_n27596_ = ~new_n26758_ & new_n27015_;
  assign new_n27597_ = ~new_n27011_ & new_n27596_;
  assign new_n27598_ = ~new_n27012_ & ~new_n27015_;
  assign new_n27599_ = ~new_n27597_ & ~new_n27598_;
  assign new_n27600_ = \quotient[2]  & ~new_n27599_;
  assign new_n27601_ = ~new_n26748_ & ~new_n27234_;
  assign new_n27602_ = ~new_n27233_ & new_n27601_;
  assign new_n27603_ = ~new_n27600_ & ~new_n27602_;
  assign new_n27604_ = ~\b[21]  & ~new_n27603_;
  assign new_n27605_ = ~new_n26767_ & new_n27010_;
  assign new_n27606_ = ~new_n27006_ & new_n27605_;
  assign new_n27607_ = ~new_n27007_ & ~new_n27010_;
  assign new_n27608_ = ~new_n27606_ & ~new_n27607_;
  assign new_n27609_ = \quotient[2]  & ~new_n27608_;
  assign new_n27610_ = ~new_n26757_ & ~new_n27234_;
  assign new_n27611_ = ~new_n27233_ & new_n27610_;
  assign new_n27612_ = ~new_n27609_ & ~new_n27611_;
  assign new_n27613_ = ~\b[20]  & ~new_n27612_;
  assign new_n27614_ = ~new_n26776_ & new_n27005_;
  assign new_n27615_ = ~new_n27001_ & new_n27614_;
  assign new_n27616_ = ~new_n27002_ & ~new_n27005_;
  assign new_n27617_ = ~new_n27615_ & ~new_n27616_;
  assign new_n27618_ = \quotient[2]  & ~new_n27617_;
  assign new_n27619_ = ~new_n26766_ & ~new_n27234_;
  assign new_n27620_ = ~new_n27233_ & new_n27619_;
  assign new_n27621_ = ~new_n27618_ & ~new_n27620_;
  assign new_n27622_ = ~\b[19]  & ~new_n27621_;
  assign new_n27623_ = ~new_n26785_ & new_n27000_;
  assign new_n27624_ = ~new_n26996_ & new_n27623_;
  assign new_n27625_ = ~new_n26997_ & ~new_n27000_;
  assign new_n27626_ = ~new_n27624_ & ~new_n27625_;
  assign new_n27627_ = \quotient[2]  & ~new_n27626_;
  assign new_n27628_ = ~new_n26775_ & ~new_n27234_;
  assign new_n27629_ = ~new_n27233_ & new_n27628_;
  assign new_n27630_ = ~new_n27627_ & ~new_n27629_;
  assign new_n27631_ = ~\b[18]  & ~new_n27630_;
  assign new_n27632_ = ~new_n26794_ & new_n26995_;
  assign new_n27633_ = ~new_n26991_ & new_n27632_;
  assign new_n27634_ = ~new_n26992_ & ~new_n26995_;
  assign new_n27635_ = ~new_n27633_ & ~new_n27634_;
  assign new_n27636_ = \quotient[2]  & ~new_n27635_;
  assign new_n27637_ = ~new_n26784_ & ~new_n27234_;
  assign new_n27638_ = ~new_n27233_ & new_n27637_;
  assign new_n27639_ = ~new_n27636_ & ~new_n27638_;
  assign new_n27640_ = ~\b[17]  & ~new_n27639_;
  assign new_n27641_ = ~new_n26803_ & new_n26990_;
  assign new_n27642_ = ~new_n26986_ & new_n27641_;
  assign new_n27643_ = ~new_n26987_ & ~new_n26990_;
  assign new_n27644_ = ~new_n27642_ & ~new_n27643_;
  assign new_n27645_ = \quotient[2]  & ~new_n27644_;
  assign new_n27646_ = ~new_n26793_ & ~new_n27234_;
  assign new_n27647_ = ~new_n27233_ & new_n27646_;
  assign new_n27648_ = ~new_n27645_ & ~new_n27647_;
  assign new_n27649_ = ~\b[16]  & ~new_n27648_;
  assign new_n27650_ = ~new_n26812_ & new_n26985_;
  assign new_n27651_ = ~new_n26981_ & new_n27650_;
  assign new_n27652_ = ~new_n26982_ & ~new_n26985_;
  assign new_n27653_ = ~new_n27651_ & ~new_n27652_;
  assign new_n27654_ = \quotient[2]  & ~new_n27653_;
  assign new_n27655_ = ~new_n26802_ & ~new_n27234_;
  assign new_n27656_ = ~new_n27233_ & new_n27655_;
  assign new_n27657_ = ~new_n27654_ & ~new_n27656_;
  assign new_n27658_ = ~\b[15]  & ~new_n27657_;
  assign new_n27659_ = ~new_n26821_ & new_n26980_;
  assign new_n27660_ = ~new_n26976_ & new_n27659_;
  assign new_n27661_ = ~new_n26977_ & ~new_n26980_;
  assign new_n27662_ = ~new_n27660_ & ~new_n27661_;
  assign new_n27663_ = \quotient[2]  & ~new_n27662_;
  assign new_n27664_ = ~new_n26811_ & ~new_n27234_;
  assign new_n27665_ = ~new_n27233_ & new_n27664_;
  assign new_n27666_ = ~new_n27663_ & ~new_n27665_;
  assign new_n27667_ = ~\b[14]  & ~new_n27666_;
  assign new_n27668_ = ~new_n26830_ & new_n26975_;
  assign new_n27669_ = ~new_n26971_ & new_n27668_;
  assign new_n27670_ = ~new_n26972_ & ~new_n26975_;
  assign new_n27671_ = ~new_n27669_ & ~new_n27670_;
  assign new_n27672_ = \quotient[2]  & ~new_n27671_;
  assign new_n27673_ = ~new_n26820_ & ~new_n27234_;
  assign new_n27674_ = ~new_n27233_ & new_n27673_;
  assign new_n27675_ = ~new_n27672_ & ~new_n27674_;
  assign new_n27676_ = ~\b[13]  & ~new_n27675_;
  assign new_n27677_ = ~new_n26839_ & new_n26970_;
  assign new_n27678_ = ~new_n26966_ & new_n27677_;
  assign new_n27679_ = ~new_n26967_ & ~new_n26970_;
  assign new_n27680_ = ~new_n27678_ & ~new_n27679_;
  assign new_n27681_ = \quotient[2]  & ~new_n27680_;
  assign new_n27682_ = ~new_n26829_ & ~new_n27234_;
  assign new_n27683_ = ~new_n27233_ & new_n27682_;
  assign new_n27684_ = ~new_n27681_ & ~new_n27683_;
  assign new_n27685_ = ~\b[12]  & ~new_n27684_;
  assign new_n27686_ = ~new_n26848_ & new_n26965_;
  assign new_n27687_ = ~new_n26961_ & new_n27686_;
  assign new_n27688_ = ~new_n26962_ & ~new_n26965_;
  assign new_n27689_ = ~new_n27687_ & ~new_n27688_;
  assign new_n27690_ = \quotient[2]  & ~new_n27689_;
  assign new_n27691_ = ~new_n26838_ & ~new_n27234_;
  assign new_n27692_ = ~new_n27233_ & new_n27691_;
  assign new_n27693_ = ~new_n27690_ & ~new_n27692_;
  assign new_n27694_ = ~\b[11]  & ~new_n27693_;
  assign new_n27695_ = ~new_n26857_ & new_n26960_;
  assign new_n27696_ = ~new_n26956_ & new_n27695_;
  assign new_n27697_ = ~new_n26957_ & ~new_n26960_;
  assign new_n27698_ = ~new_n27696_ & ~new_n27697_;
  assign new_n27699_ = \quotient[2]  & ~new_n27698_;
  assign new_n27700_ = ~new_n26847_ & ~new_n27234_;
  assign new_n27701_ = ~new_n27233_ & new_n27700_;
  assign new_n27702_ = ~new_n27699_ & ~new_n27701_;
  assign new_n27703_ = ~\b[10]  & ~new_n27702_;
  assign new_n27704_ = ~new_n26866_ & new_n26955_;
  assign new_n27705_ = ~new_n26951_ & new_n27704_;
  assign new_n27706_ = ~new_n26952_ & ~new_n26955_;
  assign new_n27707_ = ~new_n27705_ & ~new_n27706_;
  assign new_n27708_ = \quotient[2]  & ~new_n27707_;
  assign new_n27709_ = ~new_n26856_ & ~new_n27234_;
  assign new_n27710_ = ~new_n27233_ & new_n27709_;
  assign new_n27711_ = ~new_n27708_ & ~new_n27710_;
  assign new_n27712_ = ~\b[9]  & ~new_n27711_;
  assign new_n27713_ = ~new_n26875_ & new_n26950_;
  assign new_n27714_ = ~new_n26946_ & new_n27713_;
  assign new_n27715_ = ~new_n26947_ & ~new_n26950_;
  assign new_n27716_ = ~new_n27714_ & ~new_n27715_;
  assign new_n27717_ = \quotient[2]  & ~new_n27716_;
  assign new_n27718_ = ~new_n26865_ & ~new_n27234_;
  assign new_n27719_ = ~new_n27233_ & new_n27718_;
  assign new_n27720_ = ~new_n27717_ & ~new_n27719_;
  assign new_n27721_ = ~\b[8]  & ~new_n27720_;
  assign new_n27722_ = ~new_n26884_ & new_n26945_;
  assign new_n27723_ = ~new_n26941_ & new_n27722_;
  assign new_n27724_ = ~new_n26942_ & ~new_n26945_;
  assign new_n27725_ = ~new_n27723_ & ~new_n27724_;
  assign new_n27726_ = \quotient[2]  & ~new_n27725_;
  assign new_n27727_ = ~new_n26874_ & ~new_n27234_;
  assign new_n27728_ = ~new_n27233_ & new_n27727_;
  assign new_n27729_ = ~new_n27726_ & ~new_n27728_;
  assign new_n27730_ = ~\b[7]  & ~new_n27729_;
  assign new_n27731_ = ~new_n26893_ & new_n26940_;
  assign new_n27732_ = ~new_n26936_ & new_n27731_;
  assign new_n27733_ = ~new_n26937_ & ~new_n26940_;
  assign new_n27734_ = ~new_n27732_ & ~new_n27733_;
  assign new_n27735_ = \quotient[2]  & ~new_n27734_;
  assign new_n27736_ = ~new_n26883_ & ~new_n27234_;
  assign new_n27737_ = ~new_n27233_ & new_n27736_;
  assign new_n27738_ = ~new_n27735_ & ~new_n27737_;
  assign new_n27739_ = ~\b[6]  & ~new_n27738_;
  assign new_n27740_ = ~new_n26902_ & new_n26935_;
  assign new_n27741_ = ~new_n26931_ & new_n27740_;
  assign new_n27742_ = ~new_n26932_ & ~new_n26935_;
  assign new_n27743_ = ~new_n27741_ & ~new_n27742_;
  assign new_n27744_ = \quotient[2]  & ~new_n27743_;
  assign new_n27745_ = ~new_n26892_ & ~new_n27234_;
  assign new_n27746_ = ~new_n27233_ & new_n27745_;
  assign new_n27747_ = ~new_n27744_ & ~new_n27746_;
  assign new_n27748_ = ~\b[5]  & ~new_n27747_;
  assign new_n27749_ = ~new_n26910_ & new_n26930_;
  assign new_n27750_ = ~new_n26926_ & new_n27749_;
  assign new_n27751_ = ~new_n26927_ & ~new_n26930_;
  assign new_n27752_ = ~new_n27750_ & ~new_n27751_;
  assign new_n27753_ = \quotient[2]  & ~new_n27752_;
  assign new_n27754_ = ~new_n26901_ & ~new_n27234_;
  assign new_n27755_ = ~new_n27233_ & new_n27754_;
  assign new_n27756_ = ~new_n27753_ & ~new_n27755_;
  assign new_n27757_ = ~\b[4]  & ~new_n27756_;
  assign new_n27758_ = ~new_n26921_ & new_n26925_;
  assign new_n27759_ = ~new_n26920_ & new_n27758_;
  assign new_n27760_ = ~new_n26922_ & ~new_n26925_;
  assign new_n27761_ = ~new_n27759_ & ~new_n27760_;
  assign new_n27762_ = \quotient[2]  & ~new_n27761_;
  assign new_n27763_ = ~new_n26909_ & ~new_n27234_;
  assign new_n27764_ = ~new_n27233_ & new_n27763_;
  assign new_n27765_ = ~new_n27762_ & ~new_n27764_;
  assign new_n27766_ = ~\b[3]  & ~new_n27765_;
  assign new_n27767_ = ~new_n26917_ & new_n26919_;
  assign new_n27768_ = ~new_n26915_ & new_n27767_;
  assign new_n27769_ = ~new_n26920_ & ~new_n27768_;
  assign new_n27770_ = \quotient[2]  & new_n27769_;
  assign new_n27771_ = ~new_n26914_ & ~new_n27234_;
  assign new_n27772_ = ~new_n27233_ & new_n27771_;
  assign new_n27773_ = ~new_n27770_ & ~new_n27772_;
  assign new_n27774_ = ~\b[2]  & ~new_n27773_;
  assign new_n27775_ = \b[0]  & \quotient[2] ;
  assign new_n27776_ = \a[2]  & ~new_n27775_;
  assign new_n27777_ = new_n26919_ & \quotient[2] ;
  assign new_n27778_ = ~new_n27776_ & ~new_n27777_;
  assign new_n27779_ = \b[1]  & ~new_n27778_;
  assign new_n27780_ = ~\b[1]  & ~new_n27777_;
  assign new_n27781_ = ~new_n27776_ & new_n27780_;
  assign new_n27782_ = ~new_n27779_ & ~new_n27781_;
  assign new_n27783_ = ~\a[1]  & \b[0] ;
  assign new_n27784_ = ~new_n27782_ & ~new_n27783_;
  assign new_n27785_ = ~\b[1]  & ~new_n27778_;
  assign new_n27786_ = ~new_n27784_ & ~new_n27785_;
  assign new_n27787_ = \b[2]  & ~new_n27772_;
  assign new_n27788_ = ~new_n27770_ & new_n27787_;
  assign new_n27789_ = ~new_n27774_ & ~new_n27788_;
  assign new_n27790_ = ~new_n27786_ & new_n27789_;
  assign new_n27791_ = ~new_n27774_ & ~new_n27790_;
  assign new_n27792_ = \b[3]  & ~new_n27764_;
  assign new_n27793_ = ~new_n27762_ & new_n27792_;
  assign new_n27794_ = ~new_n27766_ & ~new_n27793_;
  assign new_n27795_ = ~new_n27791_ & new_n27794_;
  assign new_n27796_ = ~new_n27766_ & ~new_n27795_;
  assign new_n27797_ = \b[4]  & ~new_n27755_;
  assign new_n27798_ = ~new_n27753_ & new_n27797_;
  assign new_n27799_ = ~new_n27757_ & ~new_n27798_;
  assign new_n27800_ = ~new_n27796_ & new_n27799_;
  assign new_n27801_ = ~new_n27757_ & ~new_n27800_;
  assign new_n27802_ = \b[5]  & ~new_n27746_;
  assign new_n27803_ = ~new_n27744_ & new_n27802_;
  assign new_n27804_ = ~new_n27748_ & ~new_n27803_;
  assign new_n27805_ = ~new_n27801_ & new_n27804_;
  assign new_n27806_ = ~new_n27748_ & ~new_n27805_;
  assign new_n27807_ = \b[6]  & ~new_n27737_;
  assign new_n27808_ = ~new_n27735_ & new_n27807_;
  assign new_n27809_ = ~new_n27739_ & ~new_n27808_;
  assign new_n27810_ = ~new_n27806_ & new_n27809_;
  assign new_n27811_ = ~new_n27739_ & ~new_n27810_;
  assign new_n27812_ = \b[7]  & ~new_n27728_;
  assign new_n27813_ = ~new_n27726_ & new_n27812_;
  assign new_n27814_ = ~new_n27730_ & ~new_n27813_;
  assign new_n27815_ = ~new_n27811_ & new_n27814_;
  assign new_n27816_ = ~new_n27730_ & ~new_n27815_;
  assign new_n27817_ = \b[8]  & ~new_n27719_;
  assign new_n27818_ = ~new_n27717_ & new_n27817_;
  assign new_n27819_ = ~new_n27721_ & ~new_n27818_;
  assign new_n27820_ = ~new_n27816_ & new_n27819_;
  assign new_n27821_ = ~new_n27721_ & ~new_n27820_;
  assign new_n27822_ = \b[9]  & ~new_n27710_;
  assign new_n27823_ = ~new_n27708_ & new_n27822_;
  assign new_n27824_ = ~new_n27712_ & ~new_n27823_;
  assign new_n27825_ = ~new_n27821_ & new_n27824_;
  assign new_n27826_ = ~new_n27712_ & ~new_n27825_;
  assign new_n27827_ = \b[10]  & ~new_n27701_;
  assign new_n27828_ = ~new_n27699_ & new_n27827_;
  assign new_n27829_ = ~new_n27703_ & ~new_n27828_;
  assign new_n27830_ = ~new_n27826_ & new_n27829_;
  assign new_n27831_ = ~new_n27703_ & ~new_n27830_;
  assign new_n27832_ = \b[11]  & ~new_n27692_;
  assign new_n27833_ = ~new_n27690_ & new_n27832_;
  assign new_n27834_ = ~new_n27694_ & ~new_n27833_;
  assign new_n27835_ = ~new_n27831_ & new_n27834_;
  assign new_n27836_ = ~new_n27694_ & ~new_n27835_;
  assign new_n27837_ = \b[12]  & ~new_n27683_;
  assign new_n27838_ = ~new_n27681_ & new_n27837_;
  assign new_n27839_ = ~new_n27685_ & ~new_n27838_;
  assign new_n27840_ = ~new_n27836_ & new_n27839_;
  assign new_n27841_ = ~new_n27685_ & ~new_n27840_;
  assign new_n27842_ = \b[13]  & ~new_n27674_;
  assign new_n27843_ = ~new_n27672_ & new_n27842_;
  assign new_n27844_ = ~new_n27676_ & ~new_n27843_;
  assign new_n27845_ = ~new_n27841_ & new_n27844_;
  assign new_n27846_ = ~new_n27676_ & ~new_n27845_;
  assign new_n27847_ = \b[14]  & ~new_n27665_;
  assign new_n27848_ = ~new_n27663_ & new_n27847_;
  assign new_n27849_ = ~new_n27667_ & ~new_n27848_;
  assign new_n27850_ = ~new_n27846_ & new_n27849_;
  assign new_n27851_ = ~new_n27667_ & ~new_n27850_;
  assign new_n27852_ = \b[15]  & ~new_n27656_;
  assign new_n27853_ = ~new_n27654_ & new_n27852_;
  assign new_n27854_ = ~new_n27658_ & ~new_n27853_;
  assign new_n27855_ = ~new_n27851_ & new_n27854_;
  assign new_n27856_ = ~new_n27658_ & ~new_n27855_;
  assign new_n27857_ = \b[16]  & ~new_n27647_;
  assign new_n27858_ = ~new_n27645_ & new_n27857_;
  assign new_n27859_ = ~new_n27649_ & ~new_n27858_;
  assign new_n27860_ = ~new_n27856_ & new_n27859_;
  assign new_n27861_ = ~new_n27649_ & ~new_n27860_;
  assign new_n27862_ = \b[17]  & ~new_n27638_;
  assign new_n27863_ = ~new_n27636_ & new_n27862_;
  assign new_n27864_ = ~new_n27640_ & ~new_n27863_;
  assign new_n27865_ = ~new_n27861_ & new_n27864_;
  assign new_n27866_ = ~new_n27640_ & ~new_n27865_;
  assign new_n27867_ = \b[18]  & ~new_n27629_;
  assign new_n27868_ = ~new_n27627_ & new_n27867_;
  assign new_n27869_ = ~new_n27631_ & ~new_n27868_;
  assign new_n27870_ = ~new_n27866_ & new_n27869_;
  assign new_n27871_ = ~new_n27631_ & ~new_n27870_;
  assign new_n27872_ = \b[19]  & ~new_n27620_;
  assign new_n27873_ = ~new_n27618_ & new_n27872_;
  assign new_n27874_ = ~new_n27622_ & ~new_n27873_;
  assign new_n27875_ = ~new_n27871_ & new_n27874_;
  assign new_n27876_ = ~new_n27622_ & ~new_n27875_;
  assign new_n27877_ = \b[20]  & ~new_n27611_;
  assign new_n27878_ = ~new_n27609_ & new_n27877_;
  assign new_n27879_ = ~new_n27613_ & ~new_n27878_;
  assign new_n27880_ = ~new_n27876_ & new_n27879_;
  assign new_n27881_ = ~new_n27613_ & ~new_n27880_;
  assign new_n27882_ = \b[21]  & ~new_n27602_;
  assign new_n27883_ = ~new_n27600_ & new_n27882_;
  assign new_n27884_ = ~new_n27604_ & ~new_n27883_;
  assign new_n27885_ = ~new_n27881_ & new_n27884_;
  assign new_n27886_ = ~new_n27604_ & ~new_n27885_;
  assign new_n27887_ = \b[22]  & ~new_n27593_;
  assign new_n27888_ = ~new_n27591_ & new_n27887_;
  assign new_n27889_ = ~new_n27595_ & ~new_n27888_;
  assign new_n27890_ = ~new_n27886_ & new_n27889_;
  assign new_n27891_ = ~new_n27595_ & ~new_n27890_;
  assign new_n27892_ = \b[23]  & ~new_n27584_;
  assign new_n27893_ = ~new_n27582_ & new_n27892_;
  assign new_n27894_ = ~new_n27586_ & ~new_n27893_;
  assign new_n27895_ = ~new_n27891_ & new_n27894_;
  assign new_n27896_ = ~new_n27586_ & ~new_n27895_;
  assign new_n27897_ = \b[24]  & ~new_n27575_;
  assign new_n27898_ = ~new_n27573_ & new_n27897_;
  assign new_n27899_ = ~new_n27577_ & ~new_n27898_;
  assign new_n27900_ = ~new_n27896_ & new_n27899_;
  assign new_n27901_ = ~new_n27577_ & ~new_n27900_;
  assign new_n27902_ = \b[25]  & ~new_n27566_;
  assign new_n27903_ = ~new_n27564_ & new_n27902_;
  assign new_n27904_ = ~new_n27568_ & ~new_n27903_;
  assign new_n27905_ = ~new_n27901_ & new_n27904_;
  assign new_n27906_ = ~new_n27568_ & ~new_n27905_;
  assign new_n27907_ = \b[26]  & ~new_n27557_;
  assign new_n27908_ = ~new_n27555_ & new_n27907_;
  assign new_n27909_ = ~new_n27559_ & ~new_n27908_;
  assign new_n27910_ = ~new_n27906_ & new_n27909_;
  assign new_n27911_ = ~new_n27559_ & ~new_n27910_;
  assign new_n27912_ = \b[27]  & ~new_n27548_;
  assign new_n27913_ = ~new_n27546_ & new_n27912_;
  assign new_n27914_ = ~new_n27550_ & ~new_n27913_;
  assign new_n27915_ = ~new_n27911_ & new_n27914_;
  assign new_n27916_ = ~new_n27550_ & ~new_n27915_;
  assign new_n27917_ = \b[28]  & ~new_n27539_;
  assign new_n27918_ = ~new_n27537_ & new_n27917_;
  assign new_n27919_ = ~new_n27541_ & ~new_n27918_;
  assign new_n27920_ = ~new_n27916_ & new_n27919_;
  assign new_n27921_ = ~new_n27541_ & ~new_n27920_;
  assign new_n27922_ = \b[29]  & ~new_n27530_;
  assign new_n27923_ = ~new_n27528_ & new_n27922_;
  assign new_n27924_ = ~new_n27532_ & ~new_n27923_;
  assign new_n27925_ = ~new_n27921_ & new_n27924_;
  assign new_n27926_ = ~new_n27532_ & ~new_n27925_;
  assign new_n27927_ = \b[30]  & ~new_n27521_;
  assign new_n27928_ = ~new_n27519_ & new_n27927_;
  assign new_n27929_ = ~new_n27523_ & ~new_n27928_;
  assign new_n27930_ = ~new_n27926_ & new_n27929_;
  assign new_n27931_ = ~new_n27523_ & ~new_n27930_;
  assign new_n27932_ = \b[31]  & ~new_n27512_;
  assign new_n27933_ = ~new_n27510_ & new_n27932_;
  assign new_n27934_ = ~new_n27514_ & ~new_n27933_;
  assign new_n27935_ = ~new_n27931_ & new_n27934_;
  assign new_n27936_ = ~new_n27514_ & ~new_n27935_;
  assign new_n27937_ = \b[32]  & ~new_n27503_;
  assign new_n27938_ = ~new_n27501_ & new_n27937_;
  assign new_n27939_ = ~new_n27505_ & ~new_n27938_;
  assign new_n27940_ = ~new_n27936_ & new_n27939_;
  assign new_n27941_ = ~new_n27505_ & ~new_n27940_;
  assign new_n27942_ = \b[33]  & ~new_n27494_;
  assign new_n27943_ = ~new_n27492_ & new_n27942_;
  assign new_n27944_ = ~new_n27496_ & ~new_n27943_;
  assign new_n27945_ = ~new_n27941_ & new_n27944_;
  assign new_n27946_ = ~new_n27496_ & ~new_n27945_;
  assign new_n27947_ = \b[34]  & ~new_n27485_;
  assign new_n27948_ = ~new_n27483_ & new_n27947_;
  assign new_n27949_ = ~new_n27487_ & ~new_n27948_;
  assign new_n27950_ = ~new_n27946_ & new_n27949_;
  assign new_n27951_ = ~new_n27487_ & ~new_n27950_;
  assign new_n27952_ = \b[35]  & ~new_n27476_;
  assign new_n27953_ = ~new_n27474_ & new_n27952_;
  assign new_n27954_ = ~new_n27478_ & ~new_n27953_;
  assign new_n27955_ = ~new_n27951_ & new_n27954_;
  assign new_n27956_ = ~new_n27478_ & ~new_n27955_;
  assign new_n27957_ = \b[36]  & ~new_n27467_;
  assign new_n27958_ = ~new_n27465_ & new_n27957_;
  assign new_n27959_ = ~new_n27469_ & ~new_n27958_;
  assign new_n27960_ = ~new_n27956_ & new_n27959_;
  assign new_n27961_ = ~new_n27469_ & ~new_n27960_;
  assign new_n27962_ = \b[37]  & ~new_n27458_;
  assign new_n27963_ = ~new_n27456_ & new_n27962_;
  assign new_n27964_ = ~new_n27460_ & ~new_n27963_;
  assign new_n27965_ = ~new_n27961_ & new_n27964_;
  assign new_n27966_ = ~new_n27460_ & ~new_n27965_;
  assign new_n27967_ = \b[38]  & ~new_n27449_;
  assign new_n27968_ = ~new_n27447_ & new_n27967_;
  assign new_n27969_ = ~new_n27451_ & ~new_n27968_;
  assign new_n27970_ = ~new_n27966_ & new_n27969_;
  assign new_n27971_ = ~new_n27451_ & ~new_n27970_;
  assign new_n27972_ = \b[39]  & ~new_n27440_;
  assign new_n27973_ = ~new_n27438_ & new_n27972_;
  assign new_n27974_ = ~new_n27442_ & ~new_n27973_;
  assign new_n27975_ = ~new_n27971_ & new_n27974_;
  assign new_n27976_ = ~new_n27442_ & ~new_n27975_;
  assign new_n27977_ = \b[40]  & ~new_n27431_;
  assign new_n27978_ = ~new_n27429_ & new_n27977_;
  assign new_n27979_ = ~new_n27433_ & ~new_n27978_;
  assign new_n27980_ = ~new_n27976_ & new_n27979_;
  assign new_n27981_ = ~new_n27433_ & ~new_n27980_;
  assign new_n27982_ = \b[41]  & ~new_n27422_;
  assign new_n27983_ = ~new_n27420_ & new_n27982_;
  assign new_n27984_ = ~new_n27424_ & ~new_n27983_;
  assign new_n27985_ = ~new_n27981_ & new_n27984_;
  assign new_n27986_ = ~new_n27424_ & ~new_n27985_;
  assign new_n27987_ = \b[42]  & ~new_n27413_;
  assign new_n27988_ = ~new_n27411_ & new_n27987_;
  assign new_n27989_ = ~new_n27415_ & ~new_n27988_;
  assign new_n27990_ = ~new_n27986_ & new_n27989_;
  assign new_n27991_ = ~new_n27415_ & ~new_n27990_;
  assign new_n27992_ = \b[43]  & ~new_n27404_;
  assign new_n27993_ = ~new_n27402_ & new_n27992_;
  assign new_n27994_ = ~new_n27406_ & ~new_n27993_;
  assign new_n27995_ = ~new_n27991_ & new_n27994_;
  assign new_n27996_ = ~new_n27406_ & ~new_n27995_;
  assign new_n27997_ = \b[44]  & ~new_n27395_;
  assign new_n27998_ = ~new_n27393_ & new_n27997_;
  assign new_n27999_ = ~new_n27397_ & ~new_n27998_;
  assign new_n28000_ = ~new_n27996_ & new_n27999_;
  assign new_n28001_ = ~new_n27397_ & ~new_n28000_;
  assign new_n28002_ = \b[45]  & ~new_n27386_;
  assign new_n28003_ = ~new_n27384_ & new_n28002_;
  assign new_n28004_ = ~new_n27388_ & ~new_n28003_;
  assign new_n28005_ = ~new_n28001_ & new_n28004_;
  assign new_n28006_ = ~new_n27388_ & ~new_n28005_;
  assign new_n28007_ = \b[46]  & ~new_n27377_;
  assign new_n28008_ = ~new_n27375_ & new_n28007_;
  assign new_n28009_ = ~new_n27379_ & ~new_n28008_;
  assign new_n28010_ = ~new_n28006_ & new_n28009_;
  assign new_n28011_ = ~new_n27379_ & ~new_n28010_;
  assign new_n28012_ = \b[47]  & ~new_n27368_;
  assign new_n28013_ = ~new_n27366_ & new_n28012_;
  assign new_n28014_ = ~new_n27370_ & ~new_n28013_;
  assign new_n28015_ = ~new_n28011_ & new_n28014_;
  assign new_n28016_ = ~new_n27370_ & ~new_n28015_;
  assign new_n28017_ = \b[48]  & ~new_n27359_;
  assign new_n28018_ = ~new_n27357_ & new_n28017_;
  assign new_n28019_ = ~new_n27361_ & ~new_n28018_;
  assign new_n28020_ = ~new_n28016_ & new_n28019_;
  assign new_n28021_ = ~new_n27361_ & ~new_n28020_;
  assign new_n28022_ = \b[49]  & ~new_n27350_;
  assign new_n28023_ = ~new_n27348_ & new_n28022_;
  assign new_n28024_ = ~new_n27352_ & ~new_n28023_;
  assign new_n28025_ = ~new_n28021_ & new_n28024_;
  assign new_n28026_ = ~new_n27352_ & ~new_n28025_;
  assign new_n28027_ = \b[50]  & ~new_n27341_;
  assign new_n28028_ = ~new_n27339_ & new_n28027_;
  assign new_n28029_ = ~new_n27343_ & ~new_n28028_;
  assign new_n28030_ = ~new_n28026_ & new_n28029_;
  assign new_n28031_ = ~new_n27343_ & ~new_n28030_;
  assign new_n28032_ = \b[51]  & ~new_n27332_;
  assign new_n28033_ = ~new_n27330_ & new_n28032_;
  assign new_n28034_ = ~new_n27334_ & ~new_n28033_;
  assign new_n28035_ = ~new_n28031_ & new_n28034_;
  assign new_n28036_ = ~new_n27334_ & ~new_n28035_;
  assign new_n28037_ = \b[52]  & ~new_n27323_;
  assign new_n28038_ = ~new_n27321_ & new_n28037_;
  assign new_n28039_ = ~new_n27325_ & ~new_n28038_;
  assign new_n28040_ = ~new_n28036_ & new_n28039_;
  assign new_n28041_ = ~new_n27325_ & ~new_n28040_;
  assign new_n28042_ = \b[53]  & ~new_n27314_;
  assign new_n28043_ = ~new_n27312_ & new_n28042_;
  assign new_n28044_ = ~new_n27316_ & ~new_n28043_;
  assign new_n28045_ = ~new_n28041_ & new_n28044_;
  assign new_n28046_ = ~new_n27316_ & ~new_n28045_;
  assign new_n28047_ = \b[54]  & ~new_n27305_;
  assign new_n28048_ = ~new_n27303_ & new_n28047_;
  assign new_n28049_ = ~new_n27307_ & ~new_n28048_;
  assign new_n28050_ = ~new_n28046_ & new_n28049_;
  assign new_n28051_ = ~new_n27307_ & ~new_n28050_;
  assign new_n28052_ = \b[55]  & ~new_n27296_;
  assign new_n28053_ = ~new_n27294_ & new_n28052_;
  assign new_n28054_ = ~new_n27298_ & ~new_n28053_;
  assign new_n28055_ = ~new_n28051_ & new_n28054_;
  assign new_n28056_ = ~new_n27298_ & ~new_n28055_;
  assign new_n28057_ = \b[56]  & ~new_n27287_;
  assign new_n28058_ = ~new_n27285_ & new_n28057_;
  assign new_n28059_ = ~new_n27289_ & ~new_n28058_;
  assign new_n28060_ = ~new_n28056_ & new_n28059_;
  assign new_n28061_ = ~new_n27289_ & ~new_n28060_;
  assign new_n28062_ = \b[57]  & ~new_n27278_;
  assign new_n28063_ = ~new_n27276_ & new_n28062_;
  assign new_n28064_ = ~new_n27280_ & ~new_n28063_;
  assign new_n28065_ = ~new_n28061_ & new_n28064_;
  assign new_n28066_ = ~new_n27280_ & ~new_n28065_;
  assign new_n28067_ = \b[58]  & ~new_n27269_;
  assign new_n28068_ = ~new_n27267_ & new_n28067_;
  assign new_n28069_ = ~new_n27271_ & ~new_n28068_;
  assign new_n28070_ = ~new_n28066_ & new_n28069_;
  assign new_n28071_ = ~new_n27271_ & ~new_n28070_;
  assign new_n28072_ = \b[59]  & ~new_n27260_;
  assign new_n28073_ = ~new_n27258_ & new_n28072_;
  assign new_n28074_ = ~new_n27262_ & ~new_n28073_;
  assign new_n28075_ = ~new_n28071_ & new_n28074_;
  assign new_n28076_ = ~new_n27262_ & ~new_n28075_;
  assign new_n28077_ = \b[60]  & ~new_n27251_;
  assign new_n28078_ = ~new_n27249_ & new_n28077_;
  assign new_n28079_ = ~new_n27253_ & ~new_n28078_;
  assign new_n28080_ = ~new_n28076_ & new_n28079_;
  assign new_n28081_ = ~new_n27253_ & ~new_n28080_;
  assign new_n28082_ = \b[61]  & ~new_n27242_;
  assign new_n28083_ = ~new_n27240_ & new_n28082_;
  assign new_n28084_ = ~new_n27244_ & ~new_n28083_;
  assign new_n28085_ = ~new_n28081_ & new_n28084_;
  assign new_n28086_ = ~new_n27244_ & ~new_n28085_;
  assign new_n28087_ = ~new_n26389_ & ~new_n27230_;
  assign new_n28088_ = ~new_n27228_ & new_n28087_;
  assign new_n28089_ = ~new_n27216_ & new_n28088_;
  assign new_n28090_ = ~new_n27228_ & ~new_n27230_;
  assign new_n28091_ = ~new_n27217_ & ~new_n28090_;
  assign new_n28092_ = ~new_n28089_ & ~new_n28091_;
  assign new_n28093_ = \quotient[2]  & ~new_n28092_;
  assign new_n28094_ = ~new_n27227_ & ~new_n27234_;
  assign new_n28095_ = ~new_n27233_ & new_n28094_;
  assign new_n28096_ = ~new_n28093_ & ~new_n28095_;
  assign new_n28097_ = ~\b[62]  & ~new_n28096_;
  assign new_n28098_ = \b[62]  & ~new_n28095_;
  assign new_n28099_ = ~new_n28093_ & new_n28098_;
  assign new_n28100_ = ~\b[63]  & ~new_n28099_;
  assign new_n28101_ = ~new_n28097_ & new_n28100_;
  assign new_n28102_ = ~new_n28086_ & new_n28101_;
  assign new_n28103_ = new_n279_ & ~new_n28096_;
  assign \quotient[1]  = new_n28102_ | new_n28103_;
  assign new_n28105_ = ~new_n27262_ & new_n28079_;
  assign new_n28106_ = ~new_n28075_ & new_n28105_;
  assign new_n28107_ = ~new_n28076_ & ~new_n28079_;
  assign new_n28108_ = ~new_n28106_ & ~new_n28107_;
  assign new_n28109_ = \quotient[1]  & ~new_n28108_;
  assign new_n28110_ = ~new_n27252_ & ~new_n28103_;
  assign new_n28111_ = ~new_n28102_ & new_n28110_;
  assign new_n28112_ = ~new_n28109_ & ~new_n28111_;
  assign new_n28113_ = ~new_n27280_ & new_n28069_;
  assign new_n28114_ = ~new_n28065_ & new_n28113_;
  assign new_n28115_ = ~new_n28066_ & ~new_n28069_;
  assign new_n28116_ = ~new_n28114_ & ~new_n28115_;
  assign new_n28117_ = \quotient[1]  & ~new_n28116_;
  assign new_n28118_ = ~new_n27270_ & ~new_n28103_;
  assign new_n28119_ = ~new_n28102_ & new_n28118_;
  assign new_n28120_ = ~new_n28117_ & ~new_n28119_;
  assign new_n28121_ = ~new_n27298_ & new_n28059_;
  assign new_n28122_ = ~new_n28055_ & new_n28121_;
  assign new_n28123_ = ~new_n28056_ & ~new_n28059_;
  assign new_n28124_ = ~new_n28122_ & ~new_n28123_;
  assign new_n28125_ = \quotient[1]  & ~new_n28124_;
  assign new_n28126_ = ~new_n27288_ & ~new_n28103_;
  assign new_n28127_ = ~new_n28102_ & new_n28126_;
  assign new_n28128_ = ~new_n28125_ & ~new_n28127_;
  assign new_n28129_ = ~new_n27316_ & new_n28049_;
  assign new_n28130_ = ~new_n28045_ & new_n28129_;
  assign new_n28131_ = ~new_n28046_ & ~new_n28049_;
  assign new_n28132_ = ~new_n28130_ & ~new_n28131_;
  assign new_n28133_ = \quotient[1]  & ~new_n28132_;
  assign new_n28134_ = ~new_n27306_ & ~new_n28103_;
  assign new_n28135_ = ~new_n28102_ & new_n28134_;
  assign new_n28136_ = ~new_n28133_ & ~new_n28135_;
  assign new_n28137_ = ~new_n27334_ & new_n28039_;
  assign new_n28138_ = ~new_n28035_ & new_n28137_;
  assign new_n28139_ = ~new_n28036_ & ~new_n28039_;
  assign new_n28140_ = ~new_n28138_ & ~new_n28139_;
  assign new_n28141_ = \quotient[1]  & ~new_n28140_;
  assign new_n28142_ = ~new_n27324_ & ~new_n28103_;
  assign new_n28143_ = ~new_n28102_ & new_n28142_;
  assign new_n28144_ = ~new_n28141_ & ~new_n28143_;
  assign new_n28145_ = ~new_n27352_ & new_n28029_;
  assign new_n28146_ = ~new_n28025_ & new_n28145_;
  assign new_n28147_ = ~new_n28026_ & ~new_n28029_;
  assign new_n28148_ = ~new_n28146_ & ~new_n28147_;
  assign new_n28149_ = \quotient[1]  & ~new_n28148_;
  assign new_n28150_ = ~new_n27342_ & ~new_n28103_;
  assign new_n28151_ = ~new_n28102_ & new_n28150_;
  assign new_n28152_ = ~new_n28149_ & ~new_n28151_;
  assign new_n28153_ = ~new_n27370_ & new_n28019_;
  assign new_n28154_ = ~new_n28015_ & new_n28153_;
  assign new_n28155_ = ~new_n28016_ & ~new_n28019_;
  assign new_n28156_ = ~new_n28154_ & ~new_n28155_;
  assign new_n28157_ = \quotient[1]  & ~new_n28156_;
  assign new_n28158_ = ~new_n27360_ & ~new_n28103_;
  assign new_n28159_ = ~new_n28102_ & new_n28158_;
  assign new_n28160_ = ~new_n28157_ & ~new_n28159_;
  assign new_n28161_ = ~new_n27388_ & new_n28009_;
  assign new_n28162_ = ~new_n28005_ & new_n28161_;
  assign new_n28163_ = ~new_n28006_ & ~new_n28009_;
  assign new_n28164_ = ~new_n28162_ & ~new_n28163_;
  assign new_n28165_ = \quotient[1]  & ~new_n28164_;
  assign new_n28166_ = ~new_n27378_ & ~new_n28103_;
  assign new_n28167_ = ~new_n28102_ & new_n28166_;
  assign new_n28168_ = ~new_n28165_ & ~new_n28167_;
  assign new_n28169_ = ~new_n27406_ & new_n27999_;
  assign new_n28170_ = ~new_n27995_ & new_n28169_;
  assign new_n28171_ = ~new_n27996_ & ~new_n27999_;
  assign new_n28172_ = ~new_n28170_ & ~new_n28171_;
  assign new_n28173_ = \quotient[1]  & ~new_n28172_;
  assign new_n28174_ = ~new_n27396_ & ~new_n28103_;
  assign new_n28175_ = ~new_n28102_ & new_n28174_;
  assign new_n28176_ = ~new_n28173_ & ~new_n28175_;
  assign new_n28177_ = ~new_n27424_ & new_n27989_;
  assign new_n28178_ = ~new_n27985_ & new_n28177_;
  assign new_n28179_ = ~new_n27986_ & ~new_n27989_;
  assign new_n28180_ = ~new_n28178_ & ~new_n28179_;
  assign new_n28181_ = \quotient[1]  & ~new_n28180_;
  assign new_n28182_ = ~new_n27414_ & ~new_n28103_;
  assign new_n28183_ = ~new_n28102_ & new_n28182_;
  assign new_n28184_ = ~new_n28181_ & ~new_n28183_;
  assign new_n28185_ = ~new_n27442_ & new_n27979_;
  assign new_n28186_ = ~new_n27975_ & new_n28185_;
  assign new_n28187_ = ~new_n27976_ & ~new_n27979_;
  assign new_n28188_ = ~new_n28186_ & ~new_n28187_;
  assign new_n28189_ = \quotient[1]  & ~new_n28188_;
  assign new_n28190_ = ~new_n27432_ & ~new_n28103_;
  assign new_n28191_ = ~new_n28102_ & new_n28190_;
  assign new_n28192_ = ~new_n28189_ & ~new_n28191_;
  assign new_n28193_ = ~new_n27460_ & new_n27969_;
  assign new_n28194_ = ~new_n27965_ & new_n28193_;
  assign new_n28195_ = ~new_n27966_ & ~new_n27969_;
  assign new_n28196_ = ~new_n28194_ & ~new_n28195_;
  assign new_n28197_ = \quotient[1]  & ~new_n28196_;
  assign new_n28198_ = ~new_n27450_ & ~new_n28103_;
  assign new_n28199_ = ~new_n28102_ & new_n28198_;
  assign new_n28200_ = ~new_n28197_ & ~new_n28199_;
  assign new_n28201_ = ~new_n27478_ & new_n27959_;
  assign new_n28202_ = ~new_n27955_ & new_n28201_;
  assign new_n28203_ = ~new_n27956_ & ~new_n27959_;
  assign new_n28204_ = ~new_n28202_ & ~new_n28203_;
  assign new_n28205_ = \quotient[1]  & ~new_n28204_;
  assign new_n28206_ = ~new_n27468_ & ~new_n28103_;
  assign new_n28207_ = ~new_n28102_ & new_n28206_;
  assign new_n28208_ = ~new_n28205_ & ~new_n28207_;
  assign new_n28209_ = ~new_n27496_ & new_n27949_;
  assign new_n28210_ = ~new_n27945_ & new_n28209_;
  assign new_n28211_ = ~new_n27946_ & ~new_n27949_;
  assign new_n28212_ = ~new_n28210_ & ~new_n28211_;
  assign new_n28213_ = \quotient[1]  & ~new_n28212_;
  assign new_n28214_ = ~new_n27486_ & ~new_n28103_;
  assign new_n28215_ = ~new_n28102_ & new_n28214_;
  assign new_n28216_ = ~new_n28213_ & ~new_n28215_;
  assign new_n28217_ = ~new_n27514_ & new_n27939_;
  assign new_n28218_ = ~new_n27935_ & new_n28217_;
  assign new_n28219_ = ~new_n27936_ & ~new_n27939_;
  assign new_n28220_ = ~new_n28218_ & ~new_n28219_;
  assign new_n28221_ = \quotient[1]  & ~new_n28220_;
  assign new_n28222_ = ~new_n27504_ & ~new_n28103_;
  assign new_n28223_ = ~new_n28102_ & new_n28222_;
  assign new_n28224_ = ~new_n28221_ & ~new_n28223_;
  assign new_n28225_ = ~new_n27532_ & new_n27929_;
  assign new_n28226_ = ~new_n27925_ & new_n28225_;
  assign new_n28227_ = ~new_n27926_ & ~new_n27929_;
  assign new_n28228_ = ~new_n28226_ & ~new_n28227_;
  assign new_n28229_ = \quotient[1]  & ~new_n28228_;
  assign new_n28230_ = ~new_n27522_ & ~new_n28103_;
  assign new_n28231_ = ~new_n28102_ & new_n28230_;
  assign new_n28232_ = ~new_n28229_ & ~new_n28231_;
  assign new_n28233_ = ~new_n27550_ & new_n27919_;
  assign new_n28234_ = ~new_n27915_ & new_n28233_;
  assign new_n28235_ = ~new_n27916_ & ~new_n27919_;
  assign new_n28236_ = ~new_n28234_ & ~new_n28235_;
  assign new_n28237_ = \quotient[1]  & ~new_n28236_;
  assign new_n28238_ = ~new_n27540_ & ~new_n28103_;
  assign new_n28239_ = ~new_n28102_ & new_n28238_;
  assign new_n28240_ = ~new_n28237_ & ~new_n28239_;
  assign new_n28241_ = ~new_n27568_ & new_n27909_;
  assign new_n28242_ = ~new_n27905_ & new_n28241_;
  assign new_n28243_ = ~new_n27906_ & ~new_n27909_;
  assign new_n28244_ = ~new_n28242_ & ~new_n28243_;
  assign new_n28245_ = \quotient[1]  & ~new_n28244_;
  assign new_n28246_ = ~new_n27558_ & ~new_n28103_;
  assign new_n28247_ = ~new_n28102_ & new_n28246_;
  assign new_n28248_ = ~new_n28245_ & ~new_n28247_;
  assign new_n28249_ = ~new_n27586_ & new_n27899_;
  assign new_n28250_ = ~new_n27895_ & new_n28249_;
  assign new_n28251_ = ~new_n27896_ & ~new_n27899_;
  assign new_n28252_ = ~new_n28250_ & ~new_n28251_;
  assign new_n28253_ = \quotient[1]  & ~new_n28252_;
  assign new_n28254_ = ~new_n27576_ & ~new_n28103_;
  assign new_n28255_ = ~new_n28102_ & new_n28254_;
  assign new_n28256_ = ~new_n28253_ & ~new_n28255_;
  assign new_n28257_ = ~new_n27604_ & new_n27889_;
  assign new_n28258_ = ~new_n27885_ & new_n28257_;
  assign new_n28259_ = ~new_n27886_ & ~new_n27889_;
  assign new_n28260_ = ~new_n28258_ & ~new_n28259_;
  assign new_n28261_ = \quotient[1]  & ~new_n28260_;
  assign new_n28262_ = ~new_n27594_ & ~new_n28103_;
  assign new_n28263_ = ~new_n28102_ & new_n28262_;
  assign new_n28264_ = ~new_n28261_ & ~new_n28263_;
  assign new_n28265_ = ~new_n27622_ & new_n27879_;
  assign new_n28266_ = ~new_n27875_ & new_n28265_;
  assign new_n28267_ = ~new_n27876_ & ~new_n27879_;
  assign new_n28268_ = ~new_n28266_ & ~new_n28267_;
  assign new_n28269_ = \quotient[1]  & ~new_n28268_;
  assign new_n28270_ = ~new_n27612_ & ~new_n28103_;
  assign new_n28271_ = ~new_n28102_ & new_n28270_;
  assign new_n28272_ = ~new_n28269_ & ~new_n28271_;
  assign new_n28273_ = ~new_n27640_ & new_n27869_;
  assign new_n28274_ = ~new_n27865_ & new_n28273_;
  assign new_n28275_ = ~new_n27866_ & ~new_n27869_;
  assign new_n28276_ = ~new_n28274_ & ~new_n28275_;
  assign new_n28277_ = \quotient[1]  & ~new_n28276_;
  assign new_n28278_ = ~new_n27630_ & ~new_n28103_;
  assign new_n28279_ = ~new_n28102_ & new_n28278_;
  assign new_n28280_ = ~new_n28277_ & ~new_n28279_;
  assign new_n28281_ = ~new_n27658_ & new_n27859_;
  assign new_n28282_ = ~new_n27855_ & new_n28281_;
  assign new_n28283_ = ~new_n27856_ & ~new_n27859_;
  assign new_n28284_ = ~new_n28282_ & ~new_n28283_;
  assign new_n28285_ = \quotient[1]  & ~new_n28284_;
  assign new_n28286_ = ~new_n27648_ & ~new_n28103_;
  assign new_n28287_ = ~new_n28102_ & new_n28286_;
  assign new_n28288_ = ~new_n28285_ & ~new_n28287_;
  assign new_n28289_ = ~new_n27676_ & new_n27849_;
  assign new_n28290_ = ~new_n27845_ & new_n28289_;
  assign new_n28291_ = ~new_n27846_ & ~new_n27849_;
  assign new_n28292_ = ~new_n28290_ & ~new_n28291_;
  assign new_n28293_ = \quotient[1]  & ~new_n28292_;
  assign new_n28294_ = ~new_n27666_ & ~new_n28103_;
  assign new_n28295_ = ~new_n28102_ & new_n28294_;
  assign new_n28296_ = ~new_n28293_ & ~new_n28295_;
  assign new_n28297_ = ~new_n27694_ & new_n27839_;
  assign new_n28298_ = ~new_n27835_ & new_n28297_;
  assign new_n28299_ = ~new_n27836_ & ~new_n27839_;
  assign new_n28300_ = ~new_n28298_ & ~new_n28299_;
  assign new_n28301_ = \quotient[1]  & ~new_n28300_;
  assign new_n28302_ = ~new_n27684_ & ~new_n28103_;
  assign new_n28303_ = ~new_n28102_ & new_n28302_;
  assign new_n28304_ = ~new_n28301_ & ~new_n28303_;
  assign new_n28305_ = ~new_n27712_ & new_n27829_;
  assign new_n28306_ = ~new_n27825_ & new_n28305_;
  assign new_n28307_ = ~new_n27826_ & ~new_n27829_;
  assign new_n28308_ = ~new_n28306_ & ~new_n28307_;
  assign new_n28309_ = \quotient[1]  & ~new_n28308_;
  assign new_n28310_ = ~new_n27702_ & ~new_n28103_;
  assign new_n28311_ = ~new_n28102_ & new_n28310_;
  assign new_n28312_ = ~new_n28309_ & ~new_n28311_;
  assign new_n28313_ = ~new_n27730_ & new_n27819_;
  assign new_n28314_ = ~new_n27815_ & new_n28313_;
  assign new_n28315_ = ~new_n27816_ & ~new_n27819_;
  assign new_n28316_ = ~new_n28314_ & ~new_n28315_;
  assign new_n28317_ = \quotient[1]  & ~new_n28316_;
  assign new_n28318_ = ~new_n27720_ & ~new_n28103_;
  assign new_n28319_ = ~new_n28102_ & new_n28318_;
  assign new_n28320_ = ~new_n28317_ & ~new_n28319_;
  assign new_n28321_ = ~new_n27748_ & new_n27809_;
  assign new_n28322_ = ~new_n27805_ & new_n28321_;
  assign new_n28323_ = ~new_n27806_ & ~new_n27809_;
  assign new_n28324_ = ~new_n28322_ & ~new_n28323_;
  assign new_n28325_ = \quotient[1]  & ~new_n28324_;
  assign new_n28326_ = ~new_n27738_ & ~new_n28103_;
  assign new_n28327_ = ~new_n28102_ & new_n28326_;
  assign new_n28328_ = ~new_n28325_ & ~new_n28327_;
  assign new_n28329_ = ~new_n27766_ & new_n27799_;
  assign new_n28330_ = ~new_n27795_ & new_n28329_;
  assign new_n28331_ = ~new_n27796_ & ~new_n27799_;
  assign new_n28332_ = ~new_n28330_ & ~new_n28331_;
  assign new_n28333_ = \quotient[1]  & ~new_n28332_;
  assign new_n28334_ = ~new_n27756_ & ~new_n28103_;
  assign new_n28335_ = ~new_n28102_ & new_n28334_;
  assign new_n28336_ = ~new_n28333_ & ~new_n28335_;
  assign new_n28337_ = ~new_n27785_ & new_n27789_;
  assign new_n28338_ = ~new_n27784_ & new_n28337_;
  assign new_n28339_ = ~new_n27786_ & ~new_n27789_;
  assign new_n28340_ = ~new_n28338_ & ~new_n28339_;
  assign new_n28341_ = \quotient[1]  & ~new_n28340_;
  assign new_n28342_ = ~new_n27773_ & ~new_n28103_;
  assign new_n28343_ = ~new_n28102_ & new_n28342_;
  assign new_n28344_ = ~new_n28341_ & ~new_n28343_;
  assign new_n28345_ = ~\a[0]  & \b[0] ;
  assign new_n28346_ = \b[0]  & \quotient[1] ;
  assign new_n28347_ = \a[1]  & ~new_n28346_;
  assign new_n28348_ = new_n27783_ & \quotient[1] ;
  assign new_n28349_ = ~new_n28347_ & ~new_n28348_;
  assign new_n28350_ = ~new_n28345_ & ~new_n28349_;
  assign new_n28351_ = new_n28345_ & ~new_n28348_;
  assign new_n28352_ = ~new_n28347_ & new_n28351_;
  assign new_n28353_ = ~\b[1]  & ~new_n28352_;
  assign new_n28354_ = ~new_n27781_ & new_n27783_;
  assign new_n28355_ = ~new_n27779_ & new_n28354_;
  assign new_n28356_ = ~new_n27784_ & ~new_n28355_;
  assign new_n28357_ = \quotient[1]  & new_n28356_;
  assign new_n28358_ = ~new_n27778_ & ~new_n28103_;
  assign new_n28359_ = ~new_n28102_ & new_n28358_;
  assign new_n28360_ = ~new_n28357_ & ~new_n28359_;
  assign new_n28361_ = ~new_n28353_ & new_n28360_;
  assign new_n28362_ = ~new_n28350_ & new_n28361_;
  assign new_n28363_ = ~\b[2]  & ~new_n28362_;
  assign new_n28364_ = ~new_n28350_ & ~new_n28353_;
  assign new_n28365_ = ~new_n28360_ & ~new_n28364_;
  assign new_n28366_ = ~new_n28363_ & ~new_n28365_;
  assign new_n28367_ = ~new_n28344_ & ~new_n28366_;
  assign new_n28368_ = new_n28344_ & ~new_n28365_;
  assign new_n28369_ = ~new_n28363_ & new_n28368_;
  assign new_n28370_ = ~\b[3]  & ~new_n28369_;
  assign new_n28371_ = ~new_n27774_ & new_n27794_;
  assign new_n28372_ = ~new_n27790_ & new_n28371_;
  assign new_n28373_ = ~new_n27791_ & ~new_n27794_;
  assign new_n28374_ = ~new_n28372_ & ~new_n28373_;
  assign new_n28375_ = \quotient[1]  & ~new_n28374_;
  assign new_n28376_ = ~new_n27765_ & ~new_n28103_;
  assign new_n28377_ = ~new_n28102_ & new_n28376_;
  assign new_n28378_ = ~new_n28375_ & ~new_n28377_;
  assign new_n28379_ = ~new_n28370_ & new_n28378_;
  assign new_n28380_ = ~new_n28367_ & new_n28379_;
  assign new_n28381_ = ~\b[4]  & ~new_n28380_;
  assign new_n28382_ = ~new_n28367_ & ~new_n28370_;
  assign new_n28383_ = ~new_n28378_ & ~new_n28382_;
  assign new_n28384_ = ~new_n28381_ & ~new_n28383_;
  assign new_n28385_ = ~new_n28336_ & ~new_n28384_;
  assign new_n28386_ = new_n28336_ & ~new_n28383_;
  assign new_n28387_ = ~new_n28381_ & new_n28386_;
  assign new_n28388_ = ~\b[5]  & ~new_n28387_;
  assign new_n28389_ = ~new_n27757_ & new_n27804_;
  assign new_n28390_ = ~new_n27800_ & new_n28389_;
  assign new_n28391_ = ~new_n27801_ & ~new_n27804_;
  assign new_n28392_ = ~new_n28390_ & ~new_n28391_;
  assign new_n28393_ = \quotient[1]  & ~new_n28392_;
  assign new_n28394_ = ~new_n27747_ & ~new_n28103_;
  assign new_n28395_ = ~new_n28102_ & new_n28394_;
  assign new_n28396_ = ~new_n28393_ & ~new_n28395_;
  assign new_n28397_ = ~new_n28388_ & new_n28396_;
  assign new_n28398_ = ~new_n28385_ & new_n28397_;
  assign new_n28399_ = ~\b[6]  & ~new_n28398_;
  assign new_n28400_ = ~new_n28385_ & ~new_n28388_;
  assign new_n28401_ = ~new_n28396_ & ~new_n28400_;
  assign new_n28402_ = ~new_n28399_ & ~new_n28401_;
  assign new_n28403_ = ~new_n28328_ & ~new_n28402_;
  assign new_n28404_ = new_n28328_ & ~new_n28401_;
  assign new_n28405_ = ~new_n28399_ & new_n28404_;
  assign new_n28406_ = ~\b[7]  & ~new_n28405_;
  assign new_n28407_ = ~new_n27739_ & new_n27814_;
  assign new_n28408_ = ~new_n27810_ & new_n28407_;
  assign new_n28409_ = ~new_n27811_ & ~new_n27814_;
  assign new_n28410_ = ~new_n28408_ & ~new_n28409_;
  assign new_n28411_ = \quotient[1]  & ~new_n28410_;
  assign new_n28412_ = ~new_n27729_ & ~new_n28103_;
  assign new_n28413_ = ~new_n28102_ & new_n28412_;
  assign new_n28414_ = ~new_n28411_ & ~new_n28413_;
  assign new_n28415_ = ~new_n28406_ & new_n28414_;
  assign new_n28416_ = ~new_n28403_ & new_n28415_;
  assign new_n28417_ = ~\b[8]  & ~new_n28416_;
  assign new_n28418_ = ~new_n28403_ & ~new_n28406_;
  assign new_n28419_ = ~new_n28414_ & ~new_n28418_;
  assign new_n28420_ = ~new_n28417_ & ~new_n28419_;
  assign new_n28421_ = ~new_n28320_ & ~new_n28420_;
  assign new_n28422_ = new_n28320_ & ~new_n28419_;
  assign new_n28423_ = ~new_n28417_ & new_n28422_;
  assign new_n28424_ = ~\b[9]  & ~new_n28423_;
  assign new_n28425_ = ~new_n27721_ & new_n27824_;
  assign new_n28426_ = ~new_n27820_ & new_n28425_;
  assign new_n28427_ = ~new_n27821_ & ~new_n27824_;
  assign new_n28428_ = ~new_n28426_ & ~new_n28427_;
  assign new_n28429_ = \quotient[1]  & ~new_n28428_;
  assign new_n28430_ = ~new_n27711_ & ~new_n28103_;
  assign new_n28431_ = ~new_n28102_ & new_n28430_;
  assign new_n28432_ = ~new_n28429_ & ~new_n28431_;
  assign new_n28433_ = ~new_n28424_ & new_n28432_;
  assign new_n28434_ = ~new_n28421_ & new_n28433_;
  assign new_n28435_ = ~\b[10]  & ~new_n28434_;
  assign new_n28436_ = ~new_n28421_ & ~new_n28424_;
  assign new_n28437_ = ~new_n28432_ & ~new_n28436_;
  assign new_n28438_ = ~new_n28435_ & ~new_n28437_;
  assign new_n28439_ = ~new_n28312_ & ~new_n28438_;
  assign new_n28440_ = new_n28312_ & ~new_n28437_;
  assign new_n28441_ = ~new_n28435_ & new_n28440_;
  assign new_n28442_ = ~\b[11]  & ~new_n28441_;
  assign new_n28443_ = ~new_n27703_ & new_n27834_;
  assign new_n28444_ = ~new_n27830_ & new_n28443_;
  assign new_n28445_ = ~new_n27831_ & ~new_n27834_;
  assign new_n28446_ = ~new_n28444_ & ~new_n28445_;
  assign new_n28447_ = \quotient[1]  & ~new_n28446_;
  assign new_n28448_ = ~new_n27693_ & ~new_n28103_;
  assign new_n28449_ = ~new_n28102_ & new_n28448_;
  assign new_n28450_ = ~new_n28447_ & ~new_n28449_;
  assign new_n28451_ = ~new_n28442_ & new_n28450_;
  assign new_n28452_ = ~new_n28439_ & new_n28451_;
  assign new_n28453_ = ~\b[12]  & ~new_n28452_;
  assign new_n28454_ = ~new_n28439_ & ~new_n28442_;
  assign new_n28455_ = ~new_n28450_ & ~new_n28454_;
  assign new_n28456_ = ~new_n28453_ & ~new_n28455_;
  assign new_n28457_ = ~new_n28304_ & ~new_n28456_;
  assign new_n28458_ = new_n28304_ & ~new_n28455_;
  assign new_n28459_ = ~new_n28453_ & new_n28458_;
  assign new_n28460_ = ~\b[13]  & ~new_n28459_;
  assign new_n28461_ = ~new_n27685_ & new_n27844_;
  assign new_n28462_ = ~new_n27840_ & new_n28461_;
  assign new_n28463_ = ~new_n27841_ & ~new_n27844_;
  assign new_n28464_ = ~new_n28462_ & ~new_n28463_;
  assign new_n28465_ = \quotient[1]  & ~new_n28464_;
  assign new_n28466_ = ~new_n27675_ & ~new_n28103_;
  assign new_n28467_ = ~new_n28102_ & new_n28466_;
  assign new_n28468_ = ~new_n28465_ & ~new_n28467_;
  assign new_n28469_ = ~new_n28460_ & new_n28468_;
  assign new_n28470_ = ~new_n28457_ & new_n28469_;
  assign new_n28471_ = ~\b[14]  & ~new_n28470_;
  assign new_n28472_ = ~new_n28457_ & ~new_n28460_;
  assign new_n28473_ = ~new_n28468_ & ~new_n28472_;
  assign new_n28474_ = ~new_n28471_ & ~new_n28473_;
  assign new_n28475_ = ~new_n28296_ & ~new_n28474_;
  assign new_n28476_ = new_n28296_ & ~new_n28473_;
  assign new_n28477_ = ~new_n28471_ & new_n28476_;
  assign new_n28478_ = ~\b[15]  & ~new_n28477_;
  assign new_n28479_ = ~new_n27667_ & new_n27854_;
  assign new_n28480_ = ~new_n27850_ & new_n28479_;
  assign new_n28481_ = ~new_n27851_ & ~new_n27854_;
  assign new_n28482_ = ~new_n28480_ & ~new_n28481_;
  assign new_n28483_ = \quotient[1]  & ~new_n28482_;
  assign new_n28484_ = ~new_n27657_ & ~new_n28103_;
  assign new_n28485_ = ~new_n28102_ & new_n28484_;
  assign new_n28486_ = ~new_n28483_ & ~new_n28485_;
  assign new_n28487_ = ~new_n28478_ & new_n28486_;
  assign new_n28488_ = ~new_n28475_ & new_n28487_;
  assign new_n28489_ = ~\b[16]  & ~new_n28488_;
  assign new_n28490_ = ~new_n28475_ & ~new_n28478_;
  assign new_n28491_ = ~new_n28486_ & ~new_n28490_;
  assign new_n28492_ = ~new_n28489_ & ~new_n28491_;
  assign new_n28493_ = ~new_n28288_ & ~new_n28492_;
  assign new_n28494_ = new_n28288_ & ~new_n28491_;
  assign new_n28495_ = ~new_n28489_ & new_n28494_;
  assign new_n28496_ = ~\b[17]  & ~new_n28495_;
  assign new_n28497_ = ~new_n27649_ & new_n27864_;
  assign new_n28498_ = ~new_n27860_ & new_n28497_;
  assign new_n28499_ = ~new_n27861_ & ~new_n27864_;
  assign new_n28500_ = ~new_n28498_ & ~new_n28499_;
  assign new_n28501_ = \quotient[1]  & ~new_n28500_;
  assign new_n28502_ = ~new_n27639_ & ~new_n28103_;
  assign new_n28503_ = ~new_n28102_ & new_n28502_;
  assign new_n28504_ = ~new_n28501_ & ~new_n28503_;
  assign new_n28505_ = ~new_n28496_ & new_n28504_;
  assign new_n28506_ = ~new_n28493_ & new_n28505_;
  assign new_n28507_ = ~\b[18]  & ~new_n28506_;
  assign new_n28508_ = ~new_n28493_ & ~new_n28496_;
  assign new_n28509_ = ~new_n28504_ & ~new_n28508_;
  assign new_n28510_ = ~new_n28507_ & ~new_n28509_;
  assign new_n28511_ = ~new_n28280_ & ~new_n28510_;
  assign new_n28512_ = new_n28280_ & ~new_n28509_;
  assign new_n28513_ = ~new_n28507_ & new_n28512_;
  assign new_n28514_ = ~\b[19]  & ~new_n28513_;
  assign new_n28515_ = ~new_n27631_ & new_n27874_;
  assign new_n28516_ = ~new_n27870_ & new_n28515_;
  assign new_n28517_ = ~new_n27871_ & ~new_n27874_;
  assign new_n28518_ = ~new_n28516_ & ~new_n28517_;
  assign new_n28519_ = \quotient[1]  & ~new_n28518_;
  assign new_n28520_ = ~new_n27621_ & ~new_n28103_;
  assign new_n28521_ = ~new_n28102_ & new_n28520_;
  assign new_n28522_ = ~new_n28519_ & ~new_n28521_;
  assign new_n28523_ = ~new_n28514_ & new_n28522_;
  assign new_n28524_ = ~new_n28511_ & new_n28523_;
  assign new_n28525_ = ~\b[20]  & ~new_n28524_;
  assign new_n28526_ = ~new_n28511_ & ~new_n28514_;
  assign new_n28527_ = ~new_n28522_ & ~new_n28526_;
  assign new_n28528_ = ~new_n28525_ & ~new_n28527_;
  assign new_n28529_ = ~new_n28272_ & ~new_n28528_;
  assign new_n28530_ = new_n28272_ & ~new_n28527_;
  assign new_n28531_ = ~new_n28525_ & new_n28530_;
  assign new_n28532_ = ~\b[21]  & ~new_n28531_;
  assign new_n28533_ = ~new_n27613_ & new_n27884_;
  assign new_n28534_ = ~new_n27880_ & new_n28533_;
  assign new_n28535_ = ~new_n27881_ & ~new_n27884_;
  assign new_n28536_ = ~new_n28534_ & ~new_n28535_;
  assign new_n28537_ = \quotient[1]  & ~new_n28536_;
  assign new_n28538_ = ~new_n27603_ & ~new_n28103_;
  assign new_n28539_ = ~new_n28102_ & new_n28538_;
  assign new_n28540_ = ~new_n28537_ & ~new_n28539_;
  assign new_n28541_ = ~new_n28532_ & new_n28540_;
  assign new_n28542_ = ~new_n28529_ & new_n28541_;
  assign new_n28543_ = ~\b[22]  & ~new_n28542_;
  assign new_n28544_ = ~new_n28529_ & ~new_n28532_;
  assign new_n28545_ = ~new_n28540_ & ~new_n28544_;
  assign new_n28546_ = ~new_n28543_ & ~new_n28545_;
  assign new_n28547_ = ~new_n28264_ & ~new_n28546_;
  assign new_n28548_ = new_n28264_ & ~new_n28545_;
  assign new_n28549_ = ~new_n28543_ & new_n28548_;
  assign new_n28550_ = ~\b[23]  & ~new_n28549_;
  assign new_n28551_ = ~new_n27595_ & new_n27894_;
  assign new_n28552_ = ~new_n27890_ & new_n28551_;
  assign new_n28553_ = ~new_n27891_ & ~new_n27894_;
  assign new_n28554_ = ~new_n28552_ & ~new_n28553_;
  assign new_n28555_ = \quotient[1]  & ~new_n28554_;
  assign new_n28556_ = ~new_n27585_ & ~new_n28103_;
  assign new_n28557_ = ~new_n28102_ & new_n28556_;
  assign new_n28558_ = ~new_n28555_ & ~new_n28557_;
  assign new_n28559_ = ~new_n28550_ & new_n28558_;
  assign new_n28560_ = ~new_n28547_ & new_n28559_;
  assign new_n28561_ = ~\b[24]  & ~new_n28560_;
  assign new_n28562_ = ~new_n28547_ & ~new_n28550_;
  assign new_n28563_ = ~new_n28558_ & ~new_n28562_;
  assign new_n28564_ = ~new_n28561_ & ~new_n28563_;
  assign new_n28565_ = ~new_n28256_ & ~new_n28564_;
  assign new_n28566_ = new_n28256_ & ~new_n28563_;
  assign new_n28567_ = ~new_n28561_ & new_n28566_;
  assign new_n28568_ = ~\b[25]  & ~new_n28567_;
  assign new_n28569_ = ~new_n27577_ & new_n27904_;
  assign new_n28570_ = ~new_n27900_ & new_n28569_;
  assign new_n28571_ = ~new_n27901_ & ~new_n27904_;
  assign new_n28572_ = ~new_n28570_ & ~new_n28571_;
  assign new_n28573_ = \quotient[1]  & ~new_n28572_;
  assign new_n28574_ = ~new_n27567_ & ~new_n28103_;
  assign new_n28575_ = ~new_n28102_ & new_n28574_;
  assign new_n28576_ = ~new_n28573_ & ~new_n28575_;
  assign new_n28577_ = ~new_n28568_ & new_n28576_;
  assign new_n28578_ = ~new_n28565_ & new_n28577_;
  assign new_n28579_ = ~\b[26]  & ~new_n28578_;
  assign new_n28580_ = ~new_n28565_ & ~new_n28568_;
  assign new_n28581_ = ~new_n28576_ & ~new_n28580_;
  assign new_n28582_ = ~new_n28579_ & ~new_n28581_;
  assign new_n28583_ = ~new_n28248_ & ~new_n28582_;
  assign new_n28584_ = new_n28248_ & ~new_n28581_;
  assign new_n28585_ = ~new_n28579_ & new_n28584_;
  assign new_n28586_ = ~\b[27]  & ~new_n28585_;
  assign new_n28587_ = ~new_n27559_ & new_n27914_;
  assign new_n28588_ = ~new_n27910_ & new_n28587_;
  assign new_n28589_ = ~new_n27911_ & ~new_n27914_;
  assign new_n28590_ = ~new_n28588_ & ~new_n28589_;
  assign new_n28591_ = \quotient[1]  & ~new_n28590_;
  assign new_n28592_ = ~new_n27549_ & ~new_n28103_;
  assign new_n28593_ = ~new_n28102_ & new_n28592_;
  assign new_n28594_ = ~new_n28591_ & ~new_n28593_;
  assign new_n28595_ = ~new_n28586_ & new_n28594_;
  assign new_n28596_ = ~new_n28583_ & new_n28595_;
  assign new_n28597_ = ~\b[28]  & ~new_n28596_;
  assign new_n28598_ = ~new_n28583_ & ~new_n28586_;
  assign new_n28599_ = ~new_n28594_ & ~new_n28598_;
  assign new_n28600_ = ~new_n28597_ & ~new_n28599_;
  assign new_n28601_ = ~new_n28240_ & ~new_n28600_;
  assign new_n28602_ = new_n28240_ & ~new_n28599_;
  assign new_n28603_ = ~new_n28597_ & new_n28602_;
  assign new_n28604_ = ~\b[29]  & ~new_n28603_;
  assign new_n28605_ = ~new_n27541_ & new_n27924_;
  assign new_n28606_ = ~new_n27920_ & new_n28605_;
  assign new_n28607_ = ~new_n27921_ & ~new_n27924_;
  assign new_n28608_ = ~new_n28606_ & ~new_n28607_;
  assign new_n28609_ = \quotient[1]  & ~new_n28608_;
  assign new_n28610_ = ~new_n27531_ & ~new_n28103_;
  assign new_n28611_ = ~new_n28102_ & new_n28610_;
  assign new_n28612_ = ~new_n28609_ & ~new_n28611_;
  assign new_n28613_ = ~new_n28604_ & new_n28612_;
  assign new_n28614_ = ~new_n28601_ & new_n28613_;
  assign new_n28615_ = ~\b[30]  & ~new_n28614_;
  assign new_n28616_ = ~new_n28601_ & ~new_n28604_;
  assign new_n28617_ = ~new_n28612_ & ~new_n28616_;
  assign new_n28618_ = ~new_n28615_ & ~new_n28617_;
  assign new_n28619_ = ~new_n28232_ & ~new_n28618_;
  assign new_n28620_ = new_n28232_ & ~new_n28617_;
  assign new_n28621_ = ~new_n28615_ & new_n28620_;
  assign new_n28622_ = ~\b[31]  & ~new_n28621_;
  assign new_n28623_ = ~new_n27523_ & new_n27934_;
  assign new_n28624_ = ~new_n27930_ & new_n28623_;
  assign new_n28625_ = ~new_n27931_ & ~new_n27934_;
  assign new_n28626_ = ~new_n28624_ & ~new_n28625_;
  assign new_n28627_ = \quotient[1]  & ~new_n28626_;
  assign new_n28628_ = ~new_n27513_ & ~new_n28103_;
  assign new_n28629_ = ~new_n28102_ & new_n28628_;
  assign new_n28630_ = ~new_n28627_ & ~new_n28629_;
  assign new_n28631_ = ~new_n28622_ & new_n28630_;
  assign new_n28632_ = ~new_n28619_ & new_n28631_;
  assign new_n28633_ = ~\b[32]  & ~new_n28632_;
  assign new_n28634_ = ~new_n28619_ & ~new_n28622_;
  assign new_n28635_ = ~new_n28630_ & ~new_n28634_;
  assign new_n28636_ = ~new_n28633_ & ~new_n28635_;
  assign new_n28637_ = ~new_n28224_ & ~new_n28636_;
  assign new_n28638_ = new_n28224_ & ~new_n28635_;
  assign new_n28639_ = ~new_n28633_ & new_n28638_;
  assign new_n28640_ = ~\b[33]  & ~new_n28639_;
  assign new_n28641_ = ~new_n27505_ & new_n27944_;
  assign new_n28642_ = ~new_n27940_ & new_n28641_;
  assign new_n28643_ = ~new_n27941_ & ~new_n27944_;
  assign new_n28644_ = ~new_n28642_ & ~new_n28643_;
  assign new_n28645_ = \quotient[1]  & ~new_n28644_;
  assign new_n28646_ = ~new_n27495_ & ~new_n28103_;
  assign new_n28647_ = ~new_n28102_ & new_n28646_;
  assign new_n28648_ = ~new_n28645_ & ~new_n28647_;
  assign new_n28649_ = ~new_n28640_ & new_n28648_;
  assign new_n28650_ = ~new_n28637_ & new_n28649_;
  assign new_n28651_ = ~\b[34]  & ~new_n28650_;
  assign new_n28652_ = ~new_n28637_ & ~new_n28640_;
  assign new_n28653_ = ~new_n28648_ & ~new_n28652_;
  assign new_n28654_ = ~new_n28651_ & ~new_n28653_;
  assign new_n28655_ = ~new_n28216_ & ~new_n28654_;
  assign new_n28656_ = new_n28216_ & ~new_n28653_;
  assign new_n28657_ = ~new_n28651_ & new_n28656_;
  assign new_n28658_ = ~\b[35]  & ~new_n28657_;
  assign new_n28659_ = ~new_n27487_ & new_n27954_;
  assign new_n28660_ = ~new_n27950_ & new_n28659_;
  assign new_n28661_ = ~new_n27951_ & ~new_n27954_;
  assign new_n28662_ = ~new_n28660_ & ~new_n28661_;
  assign new_n28663_ = \quotient[1]  & ~new_n28662_;
  assign new_n28664_ = ~new_n27477_ & ~new_n28103_;
  assign new_n28665_ = ~new_n28102_ & new_n28664_;
  assign new_n28666_ = ~new_n28663_ & ~new_n28665_;
  assign new_n28667_ = ~new_n28658_ & new_n28666_;
  assign new_n28668_ = ~new_n28655_ & new_n28667_;
  assign new_n28669_ = ~\b[36]  & ~new_n28668_;
  assign new_n28670_ = ~new_n28655_ & ~new_n28658_;
  assign new_n28671_ = ~new_n28666_ & ~new_n28670_;
  assign new_n28672_ = ~new_n28669_ & ~new_n28671_;
  assign new_n28673_ = ~new_n28208_ & ~new_n28672_;
  assign new_n28674_ = new_n28208_ & ~new_n28671_;
  assign new_n28675_ = ~new_n28669_ & new_n28674_;
  assign new_n28676_ = ~\b[37]  & ~new_n28675_;
  assign new_n28677_ = ~new_n27469_ & new_n27964_;
  assign new_n28678_ = ~new_n27960_ & new_n28677_;
  assign new_n28679_ = ~new_n27961_ & ~new_n27964_;
  assign new_n28680_ = ~new_n28678_ & ~new_n28679_;
  assign new_n28681_ = \quotient[1]  & ~new_n28680_;
  assign new_n28682_ = ~new_n27459_ & ~new_n28103_;
  assign new_n28683_ = ~new_n28102_ & new_n28682_;
  assign new_n28684_ = ~new_n28681_ & ~new_n28683_;
  assign new_n28685_ = ~new_n28676_ & new_n28684_;
  assign new_n28686_ = ~new_n28673_ & new_n28685_;
  assign new_n28687_ = ~\b[38]  & ~new_n28686_;
  assign new_n28688_ = ~new_n28673_ & ~new_n28676_;
  assign new_n28689_ = ~new_n28684_ & ~new_n28688_;
  assign new_n28690_ = ~new_n28687_ & ~new_n28689_;
  assign new_n28691_ = ~new_n28200_ & ~new_n28690_;
  assign new_n28692_ = new_n28200_ & ~new_n28689_;
  assign new_n28693_ = ~new_n28687_ & new_n28692_;
  assign new_n28694_ = ~\b[39]  & ~new_n28693_;
  assign new_n28695_ = ~new_n27451_ & new_n27974_;
  assign new_n28696_ = ~new_n27970_ & new_n28695_;
  assign new_n28697_ = ~new_n27971_ & ~new_n27974_;
  assign new_n28698_ = ~new_n28696_ & ~new_n28697_;
  assign new_n28699_ = \quotient[1]  & ~new_n28698_;
  assign new_n28700_ = ~new_n27441_ & ~new_n28103_;
  assign new_n28701_ = ~new_n28102_ & new_n28700_;
  assign new_n28702_ = ~new_n28699_ & ~new_n28701_;
  assign new_n28703_ = ~new_n28694_ & new_n28702_;
  assign new_n28704_ = ~new_n28691_ & new_n28703_;
  assign new_n28705_ = ~\b[40]  & ~new_n28704_;
  assign new_n28706_ = ~new_n28691_ & ~new_n28694_;
  assign new_n28707_ = ~new_n28702_ & ~new_n28706_;
  assign new_n28708_ = ~new_n28705_ & ~new_n28707_;
  assign new_n28709_ = ~new_n28192_ & ~new_n28708_;
  assign new_n28710_ = new_n28192_ & ~new_n28707_;
  assign new_n28711_ = ~new_n28705_ & new_n28710_;
  assign new_n28712_ = ~\b[41]  & ~new_n28711_;
  assign new_n28713_ = ~new_n27433_ & new_n27984_;
  assign new_n28714_ = ~new_n27980_ & new_n28713_;
  assign new_n28715_ = ~new_n27981_ & ~new_n27984_;
  assign new_n28716_ = ~new_n28714_ & ~new_n28715_;
  assign new_n28717_ = \quotient[1]  & ~new_n28716_;
  assign new_n28718_ = ~new_n27423_ & ~new_n28103_;
  assign new_n28719_ = ~new_n28102_ & new_n28718_;
  assign new_n28720_ = ~new_n28717_ & ~new_n28719_;
  assign new_n28721_ = ~new_n28712_ & new_n28720_;
  assign new_n28722_ = ~new_n28709_ & new_n28721_;
  assign new_n28723_ = ~\b[42]  & ~new_n28722_;
  assign new_n28724_ = ~new_n28709_ & ~new_n28712_;
  assign new_n28725_ = ~new_n28720_ & ~new_n28724_;
  assign new_n28726_ = ~new_n28723_ & ~new_n28725_;
  assign new_n28727_ = ~new_n28184_ & ~new_n28726_;
  assign new_n28728_ = new_n28184_ & ~new_n28725_;
  assign new_n28729_ = ~new_n28723_ & new_n28728_;
  assign new_n28730_ = ~\b[43]  & ~new_n28729_;
  assign new_n28731_ = ~new_n27415_ & new_n27994_;
  assign new_n28732_ = ~new_n27990_ & new_n28731_;
  assign new_n28733_ = ~new_n27991_ & ~new_n27994_;
  assign new_n28734_ = ~new_n28732_ & ~new_n28733_;
  assign new_n28735_ = \quotient[1]  & ~new_n28734_;
  assign new_n28736_ = ~new_n27405_ & ~new_n28103_;
  assign new_n28737_ = ~new_n28102_ & new_n28736_;
  assign new_n28738_ = ~new_n28735_ & ~new_n28737_;
  assign new_n28739_ = ~new_n28730_ & new_n28738_;
  assign new_n28740_ = ~new_n28727_ & new_n28739_;
  assign new_n28741_ = ~\b[44]  & ~new_n28740_;
  assign new_n28742_ = ~new_n28727_ & ~new_n28730_;
  assign new_n28743_ = ~new_n28738_ & ~new_n28742_;
  assign new_n28744_ = ~new_n28741_ & ~new_n28743_;
  assign new_n28745_ = ~new_n28176_ & ~new_n28744_;
  assign new_n28746_ = new_n28176_ & ~new_n28743_;
  assign new_n28747_ = ~new_n28741_ & new_n28746_;
  assign new_n28748_ = ~\b[45]  & ~new_n28747_;
  assign new_n28749_ = ~new_n27397_ & new_n28004_;
  assign new_n28750_ = ~new_n28000_ & new_n28749_;
  assign new_n28751_ = ~new_n28001_ & ~new_n28004_;
  assign new_n28752_ = ~new_n28750_ & ~new_n28751_;
  assign new_n28753_ = \quotient[1]  & ~new_n28752_;
  assign new_n28754_ = ~new_n27387_ & ~new_n28103_;
  assign new_n28755_ = ~new_n28102_ & new_n28754_;
  assign new_n28756_ = ~new_n28753_ & ~new_n28755_;
  assign new_n28757_ = ~new_n28748_ & new_n28756_;
  assign new_n28758_ = ~new_n28745_ & new_n28757_;
  assign new_n28759_ = ~\b[46]  & ~new_n28758_;
  assign new_n28760_ = ~new_n28745_ & ~new_n28748_;
  assign new_n28761_ = ~new_n28756_ & ~new_n28760_;
  assign new_n28762_ = ~new_n28759_ & ~new_n28761_;
  assign new_n28763_ = ~new_n28168_ & ~new_n28762_;
  assign new_n28764_ = new_n28168_ & ~new_n28761_;
  assign new_n28765_ = ~new_n28759_ & new_n28764_;
  assign new_n28766_ = ~\b[47]  & ~new_n28765_;
  assign new_n28767_ = ~new_n27379_ & new_n28014_;
  assign new_n28768_ = ~new_n28010_ & new_n28767_;
  assign new_n28769_ = ~new_n28011_ & ~new_n28014_;
  assign new_n28770_ = ~new_n28768_ & ~new_n28769_;
  assign new_n28771_ = \quotient[1]  & ~new_n28770_;
  assign new_n28772_ = ~new_n27369_ & ~new_n28103_;
  assign new_n28773_ = ~new_n28102_ & new_n28772_;
  assign new_n28774_ = ~new_n28771_ & ~new_n28773_;
  assign new_n28775_ = ~new_n28766_ & new_n28774_;
  assign new_n28776_ = ~new_n28763_ & new_n28775_;
  assign new_n28777_ = ~\b[48]  & ~new_n28776_;
  assign new_n28778_ = ~new_n28763_ & ~new_n28766_;
  assign new_n28779_ = ~new_n28774_ & ~new_n28778_;
  assign new_n28780_ = ~new_n28777_ & ~new_n28779_;
  assign new_n28781_ = ~new_n28160_ & ~new_n28780_;
  assign new_n28782_ = new_n28160_ & ~new_n28779_;
  assign new_n28783_ = ~new_n28777_ & new_n28782_;
  assign new_n28784_ = ~\b[49]  & ~new_n28783_;
  assign new_n28785_ = ~new_n27361_ & new_n28024_;
  assign new_n28786_ = ~new_n28020_ & new_n28785_;
  assign new_n28787_ = ~new_n28021_ & ~new_n28024_;
  assign new_n28788_ = ~new_n28786_ & ~new_n28787_;
  assign new_n28789_ = \quotient[1]  & ~new_n28788_;
  assign new_n28790_ = ~new_n27351_ & ~new_n28103_;
  assign new_n28791_ = ~new_n28102_ & new_n28790_;
  assign new_n28792_ = ~new_n28789_ & ~new_n28791_;
  assign new_n28793_ = ~new_n28784_ & new_n28792_;
  assign new_n28794_ = ~new_n28781_ & new_n28793_;
  assign new_n28795_ = ~\b[50]  & ~new_n28794_;
  assign new_n28796_ = ~new_n28781_ & ~new_n28784_;
  assign new_n28797_ = ~new_n28792_ & ~new_n28796_;
  assign new_n28798_ = ~new_n28795_ & ~new_n28797_;
  assign new_n28799_ = ~new_n28152_ & ~new_n28798_;
  assign new_n28800_ = new_n28152_ & ~new_n28797_;
  assign new_n28801_ = ~new_n28795_ & new_n28800_;
  assign new_n28802_ = ~\b[51]  & ~new_n28801_;
  assign new_n28803_ = ~new_n27343_ & new_n28034_;
  assign new_n28804_ = ~new_n28030_ & new_n28803_;
  assign new_n28805_ = ~new_n28031_ & ~new_n28034_;
  assign new_n28806_ = ~new_n28804_ & ~new_n28805_;
  assign new_n28807_ = \quotient[1]  & ~new_n28806_;
  assign new_n28808_ = ~new_n27333_ & ~new_n28103_;
  assign new_n28809_ = ~new_n28102_ & new_n28808_;
  assign new_n28810_ = ~new_n28807_ & ~new_n28809_;
  assign new_n28811_ = ~new_n28802_ & new_n28810_;
  assign new_n28812_ = ~new_n28799_ & new_n28811_;
  assign new_n28813_ = ~\b[52]  & ~new_n28812_;
  assign new_n28814_ = ~new_n28799_ & ~new_n28802_;
  assign new_n28815_ = ~new_n28810_ & ~new_n28814_;
  assign new_n28816_ = ~new_n28813_ & ~new_n28815_;
  assign new_n28817_ = ~new_n28144_ & ~new_n28816_;
  assign new_n28818_ = new_n28144_ & ~new_n28815_;
  assign new_n28819_ = ~new_n28813_ & new_n28818_;
  assign new_n28820_ = ~\b[53]  & ~new_n28819_;
  assign new_n28821_ = ~new_n27325_ & new_n28044_;
  assign new_n28822_ = ~new_n28040_ & new_n28821_;
  assign new_n28823_ = ~new_n28041_ & ~new_n28044_;
  assign new_n28824_ = ~new_n28822_ & ~new_n28823_;
  assign new_n28825_ = \quotient[1]  & ~new_n28824_;
  assign new_n28826_ = ~new_n27315_ & ~new_n28103_;
  assign new_n28827_ = ~new_n28102_ & new_n28826_;
  assign new_n28828_ = ~new_n28825_ & ~new_n28827_;
  assign new_n28829_ = ~new_n28820_ & new_n28828_;
  assign new_n28830_ = ~new_n28817_ & new_n28829_;
  assign new_n28831_ = ~\b[54]  & ~new_n28830_;
  assign new_n28832_ = ~new_n28817_ & ~new_n28820_;
  assign new_n28833_ = ~new_n28828_ & ~new_n28832_;
  assign new_n28834_ = ~new_n28831_ & ~new_n28833_;
  assign new_n28835_ = ~new_n28136_ & ~new_n28834_;
  assign new_n28836_ = new_n28136_ & ~new_n28833_;
  assign new_n28837_ = ~new_n28831_ & new_n28836_;
  assign new_n28838_ = ~\b[55]  & ~new_n28837_;
  assign new_n28839_ = ~new_n27307_ & new_n28054_;
  assign new_n28840_ = ~new_n28050_ & new_n28839_;
  assign new_n28841_ = ~new_n28051_ & ~new_n28054_;
  assign new_n28842_ = ~new_n28840_ & ~new_n28841_;
  assign new_n28843_ = \quotient[1]  & ~new_n28842_;
  assign new_n28844_ = ~new_n27297_ & ~new_n28103_;
  assign new_n28845_ = ~new_n28102_ & new_n28844_;
  assign new_n28846_ = ~new_n28843_ & ~new_n28845_;
  assign new_n28847_ = ~new_n28838_ & new_n28846_;
  assign new_n28848_ = ~new_n28835_ & new_n28847_;
  assign new_n28849_ = ~\b[56]  & ~new_n28848_;
  assign new_n28850_ = ~new_n28835_ & ~new_n28838_;
  assign new_n28851_ = ~new_n28846_ & ~new_n28850_;
  assign new_n28852_ = ~new_n28849_ & ~new_n28851_;
  assign new_n28853_ = ~new_n28128_ & ~new_n28852_;
  assign new_n28854_ = new_n28128_ & ~new_n28851_;
  assign new_n28855_ = ~new_n28849_ & new_n28854_;
  assign new_n28856_ = ~\b[57]  & ~new_n28855_;
  assign new_n28857_ = ~new_n27289_ & new_n28064_;
  assign new_n28858_ = ~new_n28060_ & new_n28857_;
  assign new_n28859_ = ~new_n28061_ & ~new_n28064_;
  assign new_n28860_ = ~new_n28858_ & ~new_n28859_;
  assign new_n28861_ = \quotient[1]  & ~new_n28860_;
  assign new_n28862_ = ~new_n27279_ & ~new_n28103_;
  assign new_n28863_ = ~new_n28102_ & new_n28862_;
  assign new_n28864_ = ~new_n28861_ & ~new_n28863_;
  assign new_n28865_ = ~new_n28856_ & new_n28864_;
  assign new_n28866_ = ~new_n28853_ & new_n28865_;
  assign new_n28867_ = ~\b[58]  & ~new_n28866_;
  assign new_n28868_ = ~new_n28853_ & ~new_n28856_;
  assign new_n28869_ = ~new_n28864_ & ~new_n28868_;
  assign new_n28870_ = ~new_n28867_ & ~new_n28869_;
  assign new_n28871_ = ~new_n28120_ & ~new_n28870_;
  assign new_n28872_ = new_n28120_ & ~new_n28869_;
  assign new_n28873_ = ~new_n28867_ & new_n28872_;
  assign new_n28874_ = ~\b[59]  & ~new_n28873_;
  assign new_n28875_ = ~new_n27271_ & new_n28074_;
  assign new_n28876_ = ~new_n28070_ & new_n28875_;
  assign new_n28877_ = ~new_n28071_ & ~new_n28074_;
  assign new_n28878_ = ~new_n28876_ & ~new_n28877_;
  assign new_n28879_ = \quotient[1]  & ~new_n28878_;
  assign new_n28880_ = ~new_n27261_ & ~new_n28103_;
  assign new_n28881_ = ~new_n28102_ & new_n28880_;
  assign new_n28882_ = ~new_n28879_ & ~new_n28881_;
  assign new_n28883_ = ~new_n28874_ & new_n28882_;
  assign new_n28884_ = ~new_n28871_ & new_n28883_;
  assign new_n28885_ = ~\b[60]  & ~new_n28884_;
  assign new_n28886_ = ~new_n28871_ & ~new_n28874_;
  assign new_n28887_ = ~new_n28882_ & ~new_n28886_;
  assign new_n28888_ = ~new_n28885_ & ~new_n28887_;
  assign new_n28889_ = ~new_n28112_ & ~new_n28888_;
  assign new_n28890_ = new_n28112_ & ~new_n28887_;
  assign new_n28891_ = ~new_n28885_ & new_n28890_;
  assign new_n28892_ = ~\b[61]  & ~new_n28891_;
  assign new_n28893_ = ~new_n27253_ & new_n28084_;
  assign new_n28894_ = ~new_n28080_ & new_n28893_;
  assign new_n28895_ = ~new_n28081_ & ~new_n28084_;
  assign new_n28896_ = ~new_n28894_ & ~new_n28895_;
  assign new_n28897_ = \quotient[1]  & ~new_n28896_;
  assign new_n28898_ = ~new_n27243_ & ~new_n28103_;
  assign new_n28899_ = ~new_n28102_ & new_n28898_;
  assign new_n28900_ = ~new_n28897_ & ~new_n28899_;
  assign new_n28901_ = ~new_n28892_ & new_n28900_;
  assign new_n28902_ = ~new_n28889_ & new_n28901_;
  assign new_n28903_ = ~\b[62]  & ~new_n28902_;
  assign new_n28904_ = ~new_n28889_ & ~new_n28892_;
  assign new_n28905_ = ~new_n28900_ & ~new_n28904_;
  assign new_n28906_ = ~new_n27244_ & ~new_n28099_;
  assign new_n28907_ = ~new_n28097_ & new_n28906_;
  assign new_n28908_ = ~new_n28085_ & new_n28907_;
  assign new_n28909_ = ~new_n28097_ & ~new_n28099_;
  assign new_n28910_ = ~new_n28086_ & ~new_n28909_;
  assign new_n28911_ = ~new_n28908_ & ~new_n28910_;
  assign new_n28912_ = \quotient[1]  & ~new_n28911_;
  assign new_n28913_ = ~new_n28096_ & ~new_n28103_;
  assign new_n28914_ = ~new_n28102_ & new_n28913_;
  assign new_n28915_ = ~new_n28912_ & ~new_n28914_;
  assign new_n28916_ = ~new_n28905_ & new_n28915_;
  assign new_n28917_ = ~new_n28903_ & new_n28916_;
  assign new_n28918_ = ~\b[63]  & ~new_n28917_;
  assign new_n28919_ = ~new_n28903_ & ~new_n28905_;
  assign new_n28920_ = ~new_n28915_ & ~new_n28919_;
  assign \quotient[0]  = new_n28918_ | new_n28920_;
  assign \quotient[59]  = ~new_n583_ & new_n600_;
  assign new_n28923_ = new_n334_ & new_n344_;
  assign new_n28924_ = new_n432_ & new_n28923_;
  assign \quotient[62]  = ~new_n327_ & new_n28924_;
  assign new_n28926_ = ~\b[1]  & ~\b[2] ;
  assign new_n28927_ = new_n383_ & new_n28926_;
  assign new_n28928_ = ~new_n257_ & new_n28927_;
  assign new_n28929_ = new_n592_ & new_n28928_;
  assign \quotient[63]  = new_n643_ & new_n28929_;
  assign new_n28931_ = new_n260_ & new_n267_;
  assign new_n28932_ = new_n333_ & new_n28931_;
  assign new_n28933_ = new_n344_ & new_n28932_;
  assign new_n28934_ = new_n432_ & new_n28933_;
  assign new_n28935_ = new_n324_ & ~new_n28934_;
  assign new_n28936_ = ~new_n326_ & ~new_n28935_;
  assign new_n28937_ = \a[63]  & ~new_n28934_;
  assign new_n28938_ = new_n347_ & ~new_n28937_;
  assign new_n28939_ = ~new_n28936_ & new_n28938_;
  assign new_n28940_ = new_n358_ & ~new_n28936_;
  assign new_n28941_ = new_n28937_ & ~new_n28940_;
  assign new_n28942_ = ~new_n28939_ & ~new_n28941_;
  assign new_n28943_ = new_n425_ & ~new_n28936_;
  assign new_n28944_ = \a[62]  & ~new_n28943_;
  assign new_n28945_ = new_n433_ & ~new_n28936_;
  assign new_n28946_ = ~new_n28944_ & ~new_n28945_;
  assign new_n28947_ = ~new_n363_ & ~new_n28946_;
  assign new_n28948_ = ~new_n437_ & ~new_n28947_;
  assign new_n28949_ = \b[2]  & ~new_n28939_;
  assign new_n28950_ = ~new_n28941_ & new_n28949_;
  assign new_n28951_ = ~\b[2]  & ~new_n28942_;
  assign new_n28952_ = ~new_n28950_ & ~new_n28951_;
  assign new_n28953_ = new_n28948_ & ~new_n28952_;
  assign new_n28954_ = ~\b[2]  & ~new_n28953_;
  assign new_n28955_ = ~new_n28948_ & ~new_n28950_;
  assign new_n28956_ = ~new_n28951_ & ~new_n28955_;
  assign new_n28957_ = new_n450_ & ~new_n28956_;
  assign new_n28958_ = ~new_n28954_ & new_n28957_;
  assign new_n28959_ = ~new_n28942_ & ~new_n28958_;
  assign new_n28960_ = new_n450_ & ~new_n28955_;
  assign new_n28961_ = ~new_n28953_ & new_n28960_;
  assign new_n28962_ = ~new_n28956_ & new_n28961_;
  assign new_n28963_ = \b[3]  & ~new_n28962_;
  assign new_n28964_ = ~new_n28959_ & new_n28963_;
  assign new_n28965_ = new_n467_ & ~new_n28956_;
  assign new_n28966_ = ~new_n28946_ & ~new_n28965_;
  assign new_n28967_ = new_n476_ & ~new_n28945_;
  assign new_n28968_ = ~new_n28944_ & new_n28967_;
  assign new_n28969_ = ~new_n28956_ & new_n28968_;
  assign new_n28970_ = ~new_n28966_ & ~new_n28969_;
  assign new_n28971_ = ~\b[2]  & ~new_n28970_;
  assign new_n28972_ = \b[2]  & ~new_n28969_;
  assign new_n28973_ = ~new_n28966_ & new_n28972_;
  assign new_n28974_ = new_n488_ & ~new_n28956_;
  assign new_n28975_ = \a[61]  & ~new_n28974_;
  assign new_n28976_ = new_n495_ & ~new_n28956_;
  assign new_n28977_ = ~new_n28975_ & ~new_n28976_;
  assign new_n28978_ = ~new_n499_ & ~new_n28977_;
  assign new_n28979_ = ~new_n501_ & ~new_n28978_;
  assign new_n28980_ = ~new_n28973_ & ~new_n28979_;
  assign new_n28981_ = ~new_n28971_ & ~new_n28980_;
  assign new_n28982_ = ~new_n28964_ & ~new_n28981_;
  assign new_n28983_ = ~new_n28959_ & ~new_n28962_;
  assign new_n28984_ = ~\b[3]  & ~new_n28983_;
  assign new_n28985_ = ~new_n28982_ & ~new_n28984_;
  assign new_n28986_ = ~new_n28964_ & ~new_n28984_;
  assign new_n28987_ = ~new_n28981_ & new_n28986_;
  assign new_n28988_ = new_n28981_ & ~new_n28986_;
  assign new_n28989_ = new_n513_ & ~new_n28988_;
  assign new_n28990_ = ~new_n28987_ & new_n28989_;
  assign new_n28991_ = ~new_n28985_ & new_n28990_;
  assign new_n28992_ = new_n513_ & ~new_n28985_;
  assign new_n28993_ = ~new_n28983_ & ~new_n28992_;
  assign new_n28994_ = \b[4]  & ~new_n28993_;
  assign new_n28995_ = ~new_n28991_ & new_n28994_;
  assign new_n28996_ = ~new_n28971_ & ~new_n28973_;
  assign new_n28997_ = new_n28979_ & ~new_n28996_;
  assign new_n28998_ = new_n513_ & ~new_n28980_;
  assign new_n28999_ = ~new_n28997_ & new_n28998_;
  assign new_n29000_ = ~new_n28985_ & new_n28999_;
  assign new_n29001_ = ~\b[2]  & ~new_n28997_;
  assign new_n29002_ = new_n513_ & ~new_n29001_;
  assign new_n29003_ = ~new_n28985_ & new_n29002_;
  assign new_n29004_ = ~new_n28970_ & ~new_n29003_;
  assign new_n29005_ = ~new_n29000_ & ~new_n29004_;
  assign new_n29006_ = ~\b[3]  & ~new_n29005_;
  assign new_n29007_ = \b[3]  & ~new_n29000_;
  assign new_n29008_ = ~new_n29004_ & new_n29007_;
  assign new_n29009_ = new_n543_ & ~new_n28985_;
  assign new_n29010_ = ~new_n28977_ & ~new_n29009_;
  assign new_n29011_ = new_n550_ & ~new_n28976_;
  assign new_n29012_ = ~new_n28975_ & new_n29011_;
  assign new_n29013_ = ~new_n28985_ & new_n29012_;
  assign new_n29014_ = ~new_n29010_ & ~new_n29013_;
  assign new_n29015_ = ~\b[2]  & ~new_n29014_;
  assign new_n29016_ = \b[2]  & ~new_n29013_;
  assign new_n29017_ = ~new_n29010_ & new_n29016_;
  assign new_n29018_ = new_n564_ & ~new_n28985_;
  assign new_n29019_ = \a[60]  & ~new_n29018_;
  assign new_n29020_ = new_n570_ & ~new_n28985_;
  assign new_n29021_ = ~new_n29019_ & ~new_n29020_;
  assign new_n29022_ = ~new_n559_ & ~new_n29021_;
  assign new_n29023_ = ~new_n574_ & ~new_n29022_;
  assign new_n29024_ = ~new_n29017_ & ~new_n29023_;
  assign new_n29025_ = ~new_n29015_ & ~new_n29024_;
  assign new_n29026_ = ~new_n29008_ & ~new_n29025_;
  assign new_n29027_ = ~new_n29006_ & ~new_n29026_;
  assign new_n29028_ = ~new_n28995_ & ~new_n29027_;
  assign new_n29029_ = ~new_n28991_ & ~new_n28993_;
  assign new_n29030_ = ~\b[4]  & ~new_n29029_;
  assign new_n29031_ = ~new_n29028_ & ~new_n29030_;
  assign new_n29032_ = ~new_n29006_ & ~new_n29008_;
  assign new_n29033_ = ~new_n29015_ & ~new_n29032_;
  assign new_n29034_ = ~new_n29024_ & new_n29033_;
  assign new_n29035_ = new_n600_ & ~new_n29034_;
  assign new_n29036_ = ~new_n29026_ & new_n29035_;
  assign new_n29037_ = ~new_n29031_ & new_n29036_;
  assign new_n29038_ = ~\b[3]  & ~new_n29034_;
  assign new_n29039_ = new_n600_ & ~new_n29038_;
  assign new_n29040_ = ~new_n29031_ & new_n29039_;
  assign new_n29041_ = ~new_n29005_ & ~new_n29040_;
  assign new_n29042_ = ~new_n29037_ & ~new_n29041_;
  assign new_n29043_ = \b[4]  & ~new_n29042_;
  assign new_n29044_ = ~\b[4]  & ~new_n29037_;
  assign new_n29045_ = ~new_n29041_ & new_n29044_;
  assign new_n29046_ = ~new_n29043_ & ~new_n29045_;
  assign new_n29047_ = ~new_n29015_ & ~new_n29017_;
  assign new_n29048_ = new_n29023_ & ~new_n29047_;
  assign new_n29049_ = new_n600_ & ~new_n29024_;
  assign new_n29050_ = ~new_n29048_ & new_n29049_;
  assign new_n29051_ = ~new_n29031_ & new_n29050_;
  assign new_n29052_ = ~\b[2]  & ~new_n29048_;
  assign new_n29053_ = new_n600_ & ~new_n29052_;
  assign new_n29054_ = ~new_n29031_ & new_n29053_;
  assign new_n29055_ = ~new_n29014_ & ~new_n29054_;
  assign new_n29056_ = ~new_n29051_ & ~new_n29055_;
  assign new_n29057_ = \b[3]  & ~new_n29056_;
  assign new_n29058_ = ~\b[3]  & ~new_n29051_;
  assign new_n29059_ = ~new_n29055_ & new_n29058_;
  assign new_n29060_ = ~new_n29057_ & ~new_n29059_;
  assign new_n29061_ = new_n635_ & ~new_n29031_;
  assign new_n29062_ = ~new_n29021_ & ~new_n29061_;
  assign new_n29063_ = new_n644_ & ~new_n29020_;
  assign new_n29064_ = ~new_n29019_ & new_n29063_;
  assign new_n29065_ = ~new_n29031_ & new_n29064_;
  assign new_n29066_ = ~new_n29062_ & ~new_n29065_;
  assign new_n29067_ = ~\b[2]  & ~new_n29066_;
  assign new_n29068_ = new_n655_ & ~new_n29031_;
  assign new_n29069_ = \a[59]  & ~new_n29068_;
  assign new_n29070_ = new_n661_ & ~new_n29031_;
  assign new_n29071_ = ~new_n29069_ & ~new_n29070_;
  assign new_n29072_ = \b[1]  & ~new_n29071_;
  assign new_n29073_ = ~\b[1]  & ~new_n29070_;
  assign new_n29074_ = ~new_n29069_ & new_n29073_;
  assign new_n29075_ = ~new_n29072_ & ~new_n29074_;
  assign new_n29076_ = ~new_n668_ & ~new_n29075_;
  assign new_n29077_ = ~\b[1]  & ~new_n29071_;
  assign new_n29078_ = ~new_n29076_ & ~new_n29077_;
  assign new_n29079_ = \b[2]  & ~new_n29065_;
  assign new_n29080_ = ~new_n29062_ & new_n29079_;
  assign new_n29081_ = ~new_n29067_ & ~new_n29080_;
  assign new_n29082_ = ~new_n29078_ & new_n29081_;
  assign new_n29083_ = ~new_n29067_ & ~new_n29082_;
  assign new_n29084_ = ~new_n29060_ & ~new_n29083_;
  assign new_n29085_ = ~\b[3]  & ~new_n29056_;
  assign new_n29086_ = ~new_n29084_ & ~new_n29085_;
  assign new_n29087_ = ~new_n29046_ & ~new_n29086_;
  assign new_n29088_ = ~\b[4]  & ~new_n29042_;
  assign new_n29089_ = ~new_n29087_ & ~new_n29088_;
  assign new_n29090_ = ~new_n28995_ & ~new_n29030_;
  assign new_n29091_ = ~new_n29006_ & ~new_n29090_;
  assign new_n29092_ = ~new_n29026_ & new_n29091_;
  assign new_n29093_ = new_n600_ & ~new_n29092_;
  assign new_n29094_ = ~new_n29028_ & new_n29093_;
  assign new_n29095_ = ~new_n29031_ & new_n29094_;
  assign new_n29096_ = ~\b[4]  & ~new_n29092_;
  assign new_n29097_ = new_n600_ & ~new_n29096_;
  assign new_n29098_ = ~new_n29031_ & new_n29097_;
  assign new_n29099_ = ~new_n29029_ & ~new_n29098_;
  assign new_n29100_ = ~new_n29095_ & ~new_n29099_;
  assign new_n29101_ = \b[5]  & ~new_n29100_;
  assign new_n29102_ = ~\b[5]  & ~new_n29095_;
  assign new_n29103_ = ~new_n29099_ & new_n29102_;
  assign new_n29104_ = ~new_n29101_ & ~new_n29103_;
  assign new_n29105_ = new_n701_ & ~new_n29104_;
  assign new_n29106_ = ~new_n29089_ & new_n29105_;
  assign new_n29107_ = new_n600_ & ~new_n29100_;
  assign new_n29108_ = ~new_n29106_ & ~new_n29107_;
  assign new_n29109_ = new_n29046_ & ~new_n29085_;
  assign new_n29110_ = ~new_n29084_ & new_n29109_;
  assign new_n29111_ = ~new_n29087_ & ~new_n29110_;
  assign new_n29112_ = ~new_n29108_ & new_n29111_;
  assign new_n29113_ = ~new_n29042_ & ~new_n29107_;
  assign new_n29114_ = ~new_n29106_ & new_n29113_;
  assign new_n29115_ = ~new_n29112_ & ~new_n29114_;
  assign new_n29116_ = ~new_n29089_ & ~new_n29104_;
  assign new_n29117_ = ~new_n29088_ & new_n29104_;
  assign new_n29118_ = ~new_n29087_ & new_n29117_;
  assign new_n29119_ = ~new_n29116_ & ~new_n29118_;
  assign new_n29120_ = ~new_n29108_ & new_n29119_;
  assign new_n29121_ = ~new_n29100_ & ~new_n29107_;
  assign new_n29122_ = ~new_n29106_ & new_n29121_;
  assign new_n29123_ = ~new_n29120_ & ~new_n29122_;
  assign new_n29124_ = ~\b[6]  & ~new_n29123_;
  assign new_n29125_ = ~\b[5]  & ~new_n29115_;
  assign new_n29126_ = new_n29060_ & ~new_n29067_;
  assign new_n29127_ = ~new_n29082_ & new_n29126_;
  assign new_n29128_ = ~new_n29084_ & ~new_n29127_;
  assign new_n29129_ = ~new_n29108_ & new_n29128_;
  assign new_n29130_ = ~new_n29056_ & ~new_n29107_;
  assign new_n29131_ = ~new_n29106_ & new_n29130_;
  assign new_n29132_ = ~new_n29129_ & ~new_n29131_;
  assign new_n29133_ = ~\b[4]  & ~new_n29132_;
  assign new_n29134_ = ~new_n29077_ & new_n29081_;
  assign new_n29135_ = ~new_n29076_ & new_n29134_;
  assign new_n29136_ = ~new_n29078_ & ~new_n29081_;
  assign new_n29137_ = ~new_n29135_ & ~new_n29136_;
  assign new_n29138_ = ~new_n29108_ & ~new_n29137_;
  assign new_n29139_ = ~new_n29066_ & ~new_n29107_;
  assign new_n29140_ = ~new_n29106_ & new_n29139_;
  assign new_n29141_ = ~new_n29138_ & ~new_n29140_;
  assign new_n29142_ = ~\b[3]  & ~new_n29141_;
  assign new_n29143_ = new_n668_ & ~new_n29074_;
  assign new_n29144_ = ~new_n29072_ & new_n29143_;
  assign new_n29145_ = ~new_n29076_ & ~new_n29144_;
  assign new_n29146_ = ~new_n29108_ & new_n29145_;
  assign new_n29147_ = ~new_n29071_ & ~new_n29107_;
  assign new_n29148_ = ~new_n29106_ & new_n29147_;
  assign new_n29149_ = ~new_n29146_ & ~new_n29148_;
  assign new_n29150_ = ~\b[2]  & ~new_n29149_;
  assign new_n29151_ = \b[0]  & ~new_n29108_;
  assign new_n29152_ = \a[58]  & ~new_n29151_;
  assign new_n29153_ = new_n668_ & ~new_n29108_;
  assign new_n29154_ = ~new_n29152_ & ~new_n29153_;
  assign new_n29155_ = \b[1]  & ~new_n29154_;
  assign new_n29156_ = ~\b[1]  & ~new_n29153_;
  assign new_n29157_ = ~new_n29152_ & new_n29156_;
  assign new_n29158_ = ~new_n29155_ & ~new_n29157_;
  assign new_n29159_ = ~new_n756_ & ~new_n29158_;
  assign new_n29160_ = ~\b[1]  & ~new_n29154_;
  assign new_n29161_ = ~new_n29159_ & ~new_n29160_;
  assign new_n29162_ = \b[2]  & ~new_n29148_;
  assign new_n29163_ = ~new_n29146_ & new_n29162_;
  assign new_n29164_ = ~new_n29150_ & ~new_n29163_;
  assign new_n29165_ = ~new_n29161_ & new_n29164_;
  assign new_n29166_ = ~new_n29150_ & ~new_n29165_;
  assign new_n29167_ = \b[3]  & ~new_n29140_;
  assign new_n29168_ = ~new_n29138_ & new_n29167_;
  assign new_n29169_ = ~new_n29142_ & ~new_n29168_;
  assign new_n29170_ = ~new_n29166_ & new_n29169_;
  assign new_n29171_ = ~new_n29142_ & ~new_n29170_;
  assign new_n29172_ = \b[4]  & ~new_n29131_;
  assign new_n29173_ = ~new_n29129_ & new_n29172_;
  assign new_n29174_ = ~new_n29133_ & ~new_n29173_;
  assign new_n29175_ = ~new_n29171_ & new_n29174_;
  assign new_n29176_ = ~new_n29133_ & ~new_n29175_;
  assign new_n29177_ = \b[5]  & ~new_n29114_;
  assign new_n29178_ = ~new_n29112_ & new_n29177_;
  assign new_n29179_ = ~new_n29125_ & ~new_n29178_;
  assign new_n29180_ = ~new_n29176_ & new_n29179_;
  assign new_n29181_ = ~new_n29125_ & ~new_n29180_;
  assign new_n29182_ = \b[6]  & ~new_n29122_;
  assign new_n29183_ = ~new_n29120_ & new_n29182_;
  assign new_n29184_ = ~new_n29124_ & ~new_n29183_;
  assign new_n29185_ = ~new_n29181_ & new_n29184_;
  assign new_n29186_ = ~new_n29124_ & ~new_n29185_;
  assign new_n29187_ = new_n788_ & ~new_n29186_;
  assign new_n29188_ = ~new_n29115_ & ~new_n29187_;
  assign new_n29189_ = ~new_n29133_ & new_n29179_;
  assign new_n29190_ = ~new_n29175_ & new_n29189_;
  assign new_n29191_ = ~new_n29176_ & ~new_n29179_;
  assign new_n29192_ = ~new_n29190_ & ~new_n29191_;
  assign new_n29193_ = new_n788_ & ~new_n29192_;
  assign new_n29194_ = ~new_n29186_ & new_n29193_;
  assign new_n29195_ = ~new_n29188_ & ~new_n29194_;
  assign new_n29196_ = ~new_n29123_ & ~new_n29187_;
  assign new_n29197_ = ~new_n29125_ & new_n29184_;
  assign new_n29198_ = ~new_n29180_ & new_n29197_;
  assign new_n29199_ = ~new_n29181_ & ~new_n29184_;
  assign new_n29200_ = ~new_n29198_ & ~new_n29199_;
  assign new_n29201_ = new_n29187_ & ~new_n29200_;
  assign new_n29202_ = ~new_n29196_ & ~new_n29201_;
  assign new_n29203_ = ~\b[7]  & ~new_n29202_;
  assign new_n29204_ = ~\b[6]  & ~new_n29195_;
  assign new_n29205_ = ~new_n29132_ & ~new_n29187_;
  assign new_n29206_ = ~new_n29142_ & new_n29174_;
  assign new_n29207_ = ~new_n29170_ & new_n29206_;
  assign new_n29208_ = ~new_n29171_ & ~new_n29174_;
  assign new_n29209_ = ~new_n29207_ & ~new_n29208_;
  assign new_n29210_ = new_n788_ & ~new_n29209_;
  assign new_n29211_ = ~new_n29186_ & new_n29210_;
  assign new_n29212_ = ~new_n29205_ & ~new_n29211_;
  assign new_n29213_ = ~\b[5]  & ~new_n29212_;
  assign new_n29214_ = ~new_n29141_ & ~new_n29187_;
  assign new_n29215_ = ~new_n29150_ & new_n29169_;
  assign new_n29216_ = ~new_n29165_ & new_n29215_;
  assign new_n29217_ = ~new_n29166_ & ~new_n29169_;
  assign new_n29218_ = ~new_n29216_ & ~new_n29217_;
  assign new_n29219_ = new_n788_ & ~new_n29218_;
  assign new_n29220_ = ~new_n29186_ & new_n29219_;
  assign new_n29221_ = ~new_n29214_ & ~new_n29220_;
  assign new_n29222_ = ~\b[4]  & ~new_n29221_;
  assign new_n29223_ = ~new_n29149_ & ~new_n29187_;
  assign new_n29224_ = ~new_n29160_ & new_n29164_;
  assign new_n29225_ = ~new_n29159_ & new_n29224_;
  assign new_n29226_ = ~new_n29161_ & ~new_n29164_;
  assign new_n29227_ = ~new_n29225_ & ~new_n29226_;
  assign new_n29228_ = new_n788_ & ~new_n29227_;
  assign new_n29229_ = ~new_n29186_ & new_n29228_;
  assign new_n29230_ = ~new_n29223_ & ~new_n29229_;
  assign new_n29231_ = ~\b[3]  & ~new_n29230_;
  assign new_n29232_ = ~new_n29154_ & ~new_n29187_;
  assign new_n29233_ = new_n756_ & ~new_n29157_;
  assign new_n29234_ = ~new_n29155_ & new_n29233_;
  assign new_n29235_ = new_n788_ & ~new_n29234_;
  assign new_n29236_ = ~new_n29159_ & new_n29235_;
  assign new_n29237_ = ~new_n29186_ & new_n29236_;
  assign new_n29238_ = ~new_n29232_ & ~new_n29237_;
  assign new_n29239_ = ~\b[2]  & ~new_n29238_;
  assign new_n29240_ = new_n846_ & ~new_n29186_;
  assign new_n29241_ = \a[57]  & ~new_n29240_;
  assign new_n29242_ = new_n853_ & ~new_n29186_;
  assign new_n29243_ = ~new_n29241_ & ~new_n29242_;
  assign new_n29244_ = \b[1]  & ~new_n29243_;
  assign new_n29245_ = ~\b[1]  & ~new_n29242_;
  assign new_n29246_ = ~new_n29241_ & new_n29245_;
  assign new_n29247_ = ~new_n29244_ & ~new_n29246_;
  assign new_n29248_ = ~new_n860_ & ~new_n29247_;
  assign new_n29249_ = ~\b[1]  & ~new_n29243_;
  assign new_n29250_ = ~new_n29248_ & ~new_n29249_;
  assign new_n29251_ = \b[2]  & ~new_n29237_;
  assign new_n29252_ = ~new_n29232_ & new_n29251_;
  assign new_n29253_ = ~new_n29239_ & ~new_n29252_;
  assign new_n29254_ = ~new_n29250_ & new_n29253_;
  assign new_n29255_ = ~new_n29239_ & ~new_n29254_;
  assign new_n29256_ = \b[3]  & ~new_n29229_;
  assign new_n29257_ = ~new_n29223_ & new_n29256_;
  assign new_n29258_ = ~new_n29231_ & ~new_n29257_;
  assign new_n29259_ = ~new_n29255_ & new_n29258_;
  assign new_n29260_ = ~new_n29231_ & ~new_n29259_;
  assign new_n29261_ = \b[4]  & ~new_n29220_;
  assign new_n29262_ = ~new_n29214_ & new_n29261_;
  assign new_n29263_ = ~new_n29222_ & ~new_n29262_;
  assign new_n29264_ = ~new_n29260_ & new_n29263_;
  assign new_n29265_ = ~new_n29222_ & ~new_n29264_;
  assign new_n29266_ = \b[5]  & ~new_n29211_;
  assign new_n29267_ = ~new_n29205_ & new_n29266_;
  assign new_n29268_ = ~new_n29213_ & ~new_n29267_;
  assign new_n29269_ = ~new_n29265_ & new_n29268_;
  assign new_n29270_ = ~new_n29213_ & ~new_n29269_;
  assign new_n29271_ = \b[6]  & ~new_n29194_;
  assign new_n29272_ = ~new_n29188_ & new_n29271_;
  assign new_n29273_ = ~new_n29204_ & ~new_n29272_;
  assign new_n29274_ = ~new_n29270_ & new_n29273_;
  assign new_n29275_ = ~new_n29204_ & ~new_n29274_;
  assign new_n29276_ = \b[7]  & ~new_n29196_;
  assign new_n29277_ = ~new_n29201_ & new_n29276_;
  assign new_n29278_ = ~new_n29203_ & ~new_n29277_;
  assign new_n29279_ = ~new_n29275_ & new_n29278_;
  assign new_n29280_ = ~new_n29203_ & ~new_n29279_;
  assign new_n29281_ = new_n895_ & ~new_n29280_;
  assign new_n29282_ = ~new_n29195_ & ~new_n29281_;
  assign new_n29283_ = ~new_n29213_ & new_n29273_;
  assign new_n29284_ = ~new_n29269_ & new_n29283_;
  assign new_n29285_ = ~new_n29270_ & ~new_n29273_;
  assign new_n29286_ = ~new_n29284_ & ~new_n29285_;
  assign new_n29287_ = new_n895_ & ~new_n29286_;
  assign new_n29288_ = ~new_n29280_ & new_n29287_;
  assign new_n29289_ = ~new_n29282_ & ~new_n29288_;
  assign new_n29290_ = ~\b[7]  & ~new_n29289_;
  assign new_n29291_ = ~new_n29212_ & ~new_n29281_;
  assign new_n29292_ = ~new_n29222_ & new_n29268_;
  assign new_n29293_ = ~new_n29264_ & new_n29292_;
  assign new_n29294_ = ~new_n29265_ & ~new_n29268_;
  assign new_n29295_ = ~new_n29293_ & ~new_n29294_;
  assign new_n29296_ = new_n895_ & ~new_n29295_;
  assign new_n29297_ = ~new_n29280_ & new_n29296_;
  assign new_n29298_ = ~new_n29291_ & ~new_n29297_;
  assign new_n29299_ = ~\b[6]  & ~new_n29298_;
  assign new_n29300_ = ~new_n29221_ & ~new_n29281_;
  assign new_n29301_ = ~new_n29231_ & new_n29263_;
  assign new_n29302_ = ~new_n29259_ & new_n29301_;
  assign new_n29303_ = ~new_n29260_ & ~new_n29263_;
  assign new_n29304_ = ~new_n29302_ & ~new_n29303_;
  assign new_n29305_ = new_n895_ & ~new_n29304_;
  assign new_n29306_ = ~new_n29280_ & new_n29305_;
  assign new_n29307_ = ~new_n29300_ & ~new_n29306_;
  assign new_n29308_ = ~\b[5]  & ~new_n29307_;
  assign new_n29309_ = ~new_n29230_ & ~new_n29281_;
  assign new_n29310_ = ~new_n29239_ & new_n29258_;
  assign new_n29311_ = ~new_n29254_ & new_n29310_;
  assign new_n29312_ = ~new_n29255_ & ~new_n29258_;
  assign new_n29313_ = ~new_n29311_ & ~new_n29312_;
  assign new_n29314_ = new_n895_ & ~new_n29313_;
  assign new_n29315_ = ~new_n29280_ & new_n29314_;
  assign new_n29316_ = ~new_n29309_ & ~new_n29315_;
  assign new_n29317_ = ~\b[4]  & ~new_n29316_;
  assign new_n29318_ = ~new_n29238_ & ~new_n29281_;
  assign new_n29319_ = ~new_n29249_ & new_n29253_;
  assign new_n29320_ = ~new_n29248_ & new_n29319_;
  assign new_n29321_ = ~new_n29250_ & ~new_n29253_;
  assign new_n29322_ = ~new_n29320_ & ~new_n29321_;
  assign new_n29323_ = new_n895_ & ~new_n29322_;
  assign new_n29324_ = ~new_n29280_ & new_n29323_;
  assign new_n29325_ = ~new_n29318_ & ~new_n29324_;
  assign new_n29326_ = ~\b[3]  & ~new_n29325_;
  assign new_n29327_ = ~new_n29243_ & ~new_n29281_;
  assign new_n29328_ = new_n860_ & ~new_n29246_;
  assign new_n29329_ = ~new_n29244_ & new_n29328_;
  assign new_n29330_ = new_n895_ & ~new_n29329_;
  assign new_n29331_ = ~new_n29248_ & new_n29330_;
  assign new_n29332_ = ~new_n29280_ & new_n29331_;
  assign new_n29333_ = ~new_n29327_ & ~new_n29332_;
  assign new_n29334_ = ~\b[2]  & ~new_n29333_;
  assign new_n29335_ = new_n954_ & ~new_n29280_;
  assign new_n29336_ = \a[56]  & ~new_n29335_;
  assign new_n29337_ = new_n960_ & ~new_n29280_;
  assign new_n29338_ = ~new_n29336_ & ~new_n29337_;
  assign new_n29339_ = \b[1]  & ~new_n29338_;
  assign new_n29340_ = ~\b[1]  & ~new_n29337_;
  assign new_n29341_ = ~new_n29336_ & new_n29340_;
  assign new_n29342_ = ~new_n29339_ & ~new_n29341_;
  assign new_n29343_ = ~new_n967_ & ~new_n29342_;
  assign new_n29344_ = ~\b[1]  & ~new_n29338_;
  assign new_n29345_ = ~new_n29343_ & ~new_n29344_;
  assign new_n29346_ = \b[2]  & ~new_n29332_;
  assign new_n29347_ = ~new_n29327_ & new_n29346_;
  assign new_n29348_ = ~new_n29334_ & ~new_n29347_;
  assign new_n29349_ = ~new_n29345_ & new_n29348_;
  assign new_n29350_ = ~new_n29334_ & ~new_n29349_;
  assign new_n29351_ = \b[3]  & ~new_n29324_;
  assign new_n29352_ = ~new_n29318_ & new_n29351_;
  assign new_n29353_ = ~new_n29326_ & ~new_n29352_;
  assign new_n29354_ = ~new_n29350_ & new_n29353_;
  assign new_n29355_ = ~new_n29326_ & ~new_n29354_;
  assign new_n29356_ = \b[4]  & ~new_n29315_;
  assign new_n29357_ = ~new_n29309_ & new_n29356_;
  assign new_n29358_ = ~new_n29317_ & ~new_n29357_;
  assign new_n29359_ = ~new_n29355_ & new_n29358_;
  assign new_n29360_ = ~new_n29317_ & ~new_n29359_;
  assign new_n29361_ = \b[5]  & ~new_n29306_;
  assign new_n29362_ = ~new_n29300_ & new_n29361_;
  assign new_n29363_ = ~new_n29308_ & ~new_n29362_;
  assign new_n29364_ = ~new_n29360_ & new_n29363_;
  assign new_n29365_ = ~new_n29308_ & ~new_n29364_;
  assign new_n29366_ = \b[6]  & ~new_n29297_;
  assign new_n29367_ = ~new_n29291_ & new_n29366_;
  assign new_n29368_ = ~new_n29299_ & ~new_n29367_;
  assign new_n29369_ = ~new_n29365_ & new_n29368_;
  assign new_n29370_ = ~new_n29299_ & ~new_n29369_;
  assign new_n29371_ = \b[7]  & ~new_n29288_;
  assign new_n29372_ = ~new_n29282_ & new_n29371_;
  assign new_n29373_ = ~new_n29290_ & ~new_n29372_;
  assign new_n29374_ = ~new_n29370_ & new_n29373_;
  assign new_n29375_ = ~new_n29290_ & ~new_n29374_;
  assign new_n29376_ = ~new_n29202_ & ~new_n29281_;
  assign new_n29377_ = ~new_n29204_ & new_n29278_;
  assign new_n29378_ = ~new_n29274_ & new_n29377_;
  assign new_n29379_ = ~new_n29275_ & ~new_n29278_;
  assign new_n29380_ = ~new_n29378_ & ~new_n29379_;
  assign new_n29381_ = new_n29281_ & ~new_n29380_;
  assign new_n29382_ = ~new_n29376_ & ~new_n29381_;
  assign new_n29383_ = ~\b[8]  & ~new_n29382_;
  assign new_n29384_ = \b[8]  & ~new_n29376_;
  assign new_n29385_ = ~new_n29381_ & new_n29384_;
  assign new_n29386_ = new_n1012_ & ~new_n29385_;
  assign new_n29387_ = ~new_n29383_ & new_n29386_;
  assign new_n29388_ = ~new_n29375_ & new_n29387_;
  assign new_n29389_ = new_n895_ & ~new_n29382_;
  assign new_n29390_ = ~new_n29388_ & ~new_n29389_;
  assign new_n29391_ = ~new_n29299_ & new_n29373_;
  assign new_n29392_ = ~new_n29369_ & new_n29391_;
  assign new_n29393_ = ~new_n29370_ & ~new_n29373_;
  assign new_n29394_ = ~new_n29392_ & ~new_n29393_;
  assign new_n29395_ = ~new_n29390_ & ~new_n29394_;
  assign new_n29396_ = ~new_n29289_ & ~new_n29389_;
  assign new_n29397_ = ~new_n29388_ & new_n29396_;
  assign new_n29398_ = ~new_n29395_ & ~new_n29397_;
  assign new_n29399_ = ~new_n29290_ & ~new_n29385_;
  assign new_n29400_ = ~new_n29383_ & new_n29399_;
  assign new_n29401_ = ~new_n29374_ & new_n29400_;
  assign new_n29402_ = ~new_n29383_ & ~new_n29385_;
  assign new_n29403_ = ~new_n29375_ & ~new_n29402_;
  assign new_n29404_ = ~new_n29401_ & ~new_n29403_;
  assign new_n29405_ = ~new_n29390_ & ~new_n29404_;
  assign new_n29406_ = ~new_n29382_ & ~new_n29389_;
  assign new_n29407_ = ~new_n29388_ & new_n29406_;
  assign new_n29408_ = ~new_n29405_ & ~new_n29407_;
  assign new_n29409_ = ~\b[9]  & ~new_n29408_;
  assign new_n29410_ = ~\b[8]  & ~new_n29398_;
  assign new_n29411_ = ~new_n29308_ & new_n29368_;
  assign new_n29412_ = ~new_n29364_ & new_n29411_;
  assign new_n29413_ = ~new_n29365_ & ~new_n29368_;
  assign new_n29414_ = ~new_n29412_ & ~new_n29413_;
  assign new_n29415_ = ~new_n29390_ & ~new_n29414_;
  assign new_n29416_ = ~new_n29298_ & ~new_n29389_;
  assign new_n29417_ = ~new_n29388_ & new_n29416_;
  assign new_n29418_ = ~new_n29415_ & ~new_n29417_;
  assign new_n29419_ = ~\b[7]  & ~new_n29418_;
  assign new_n29420_ = ~new_n29317_ & new_n29363_;
  assign new_n29421_ = ~new_n29359_ & new_n29420_;
  assign new_n29422_ = ~new_n29360_ & ~new_n29363_;
  assign new_n29423_ = ~new_n29421_ & ~new_n29422_;
  assign new_n29424_ = ~new_n29390_ & ~new_n29423_;
  assign new_n29425_ = ~new_n29307_ & ~new_n29389_;
  assign new_n29426_ = ~new_n29388_ & new_n29425_;
  assign new_n29427_ = ~new_n29424_ & ~new_n29426_;
  assign new_n29428_ = ~\b[6]  & ~new_n29427_;
  assign new_n29429_ = ~new_n29326_ & new_n29358_;
  assign new_n29430_ = ~new_n29354_ & new_n29429_;
  assign new_n29431_ = ~new_n29355_ & ~new_n29358_;
  assign new_n29432_ = ~new_n29430_ & ~new_n29431_;
  assign new_n29433_ = ~new_n29390_ & ~new_n29432_;
  assign new_n29434_ = ~new_n29316_ & ~new_n29389_;
  assign new_n29435_ = ~new_n29388_ & new_n29434_;
  assign new_n29436_ = ~new_n29433_ & ~new_n29435_;
  assign new_n29437_ = ~\b[5]  & ~new_n29436_;
  assign new_n29438_ = ~new_n29334_ & new_n29353_;
  assign new_n29439_ = ~new_n29349_ & new_n29438_;
  assign new_n29440_ = ~new_n29350_ & ~new_n29353_;
  assign new_n29441_ = ~new_n29439_ & ~new_n29440_;
  assign new_n29442_ = ~new_n29390_ & ~new_n29441_;
  assign new_n29443_ = ~new_n29325_ & ~new_n29389_;
  assign new_n29444_ = ~new_n29388_ & new_n29443_;
  assign new_n29445_ = ~new_n29442_ & ~new_n29444_;
  assign new_n29446_ = ~\b[4]  & ~new_n29445_;
  assign new_n29447_ = ~new_n29344_ & new_n29348_;
  assign new_n29448_ = ~new_n29343_ & new_n29447_;
  assign new_n29449_ = ~new_n29345_ & ~new_n29348_;
  assign new_n29450_ = ~new_n29448_ & ~new_n29449_;
  assign new_n29451_ = ~new_n29390_ & ~new_n29450_;
  assign new_n29452_ = ~new_n29333_ & ~new_n29389_;
  assign new_n29453_ = ~new_n29388_ & new_n29452_;
  assign new_n29454_ = ~new_n29451_ & ~new_n29453_;
  assign new_n29455_ = ~\b[3]  & ~new_n29454_;
  assign new_n29456_ = new_n967_ & ~new_n29341_;
  assign new_n29457_ = ~new_n29339_ & new_n29456_;
  assign new_n29458_ = ~new_n29343_ & ~new_n29457_;
  assign new_n29459_ = ~new_n29390_ & new_n29458_;
  assign new_n29460_ = ~new_n29338_ & ~new_n29389_;
  assign new_n29461_ = ~new_n29388_ & new_n29460_;
  assign new_n29462_ = ~new_n29459_ & ~new_n29461_;
  assign new_n29463_ = ~\b[2]  & ~new_n29462_;
  assign new_n29464_ = \b[0]  & ~new_n29390_;
  assign new_n29465_ = \a[55]  & ~new_n29464_;
  assign new_n29466_ = new_n967_ & ~new_n29390_;
  assign new_n29467_ = ~new_n29465_ & ~new_n29466_;
  assign new_n29468_ = \b[1]  & ~new_n29467_;
  assign new_n29469_ = ~\b[1]  & ~new_n29466_;
  assign new_n29470_ = ~new_n29465_ & new_n29469_;
  assign new_n29471_ = ~new_n29468_ & ~new_n29470_;
  assign new_n29472_ = ~new_n1099_ & ~new_n29471_;
  assign new_n29473_ = ~\b[1]  & ~new_n29467_;
  assign new_n29474_ = ~new_n29472_ & ~new_n29473_;
  assign new_n29475_ = \b[2]  & ~new_n29461_;
  assign new_n29476_ = ~new_n29459_ & new_n29475_;
  assign new_n29477_ = ~new_n29463_ & ~new_n29476_;
  assign new_n29478_ = ~new_n29474_ & new_n29477_;
  assign new_n29479_ = ~new_n29463_ & ~new_n29478_;
  assign new_n29480_ = \b[3]  & ~new_n29453_;
  assign new_n29481_ = ~new_n29451_ & new_n29480_;
  assign new_n29482_ = ~new_n29455_ & ~new_n29481_;
  assign new_n29483_ = ~new_n29479_ & new_n29482_;
  assign new_n29484_ = ~new_n29455_ & ~new_n29483_;
  assign new_n29485_ = \b[4]  & ~new_n29444_;
  assign new_n29486_ = ~new_n29442_ & new_n29485_;
  assign new_n29487_ = ~new_n29446_ & ~new_n29486_;
  assign new_n29488_ = ~new_n29484_ & new_n29487_;
  assign new_n29489_ = ~new_n29446_ & ~new_n29488_;
  assign new_n29490_ = \b[5]  & ~new_n29435_;
  assign new_n29491_ = ~new_n29433_ & new_n29490_;
  assign new_n29492_ = ~new_n29437_ & ~new_n29491_;
  assign new_n29493_ = ~new_n29489_ & new_n29492_;
  assign new_n29494_ = ~new_n29437_ & ~new_n29493_;
  assign new_n29495_ = \b[6]  & ~new_n29426_;
  assign new_n29496_ = ~new_n29424_ & new_n29495_;
  assign new_n29497_ = ~new_n29428_ & ~new_n29496_;
  assign new_n29498_ = ~new_n29494_ & new_n29497_;
  assign new_n29499_ = ~new_n29428_ & ~new_n29498_;
  assign new_n29500_ = \b[7]  & ~new_n29417_;
  assign new_n29501_ = ~new_n29415_ & new_n29500_;
  assign new_n29502_ = ~new_n29419_ & ~new_n29501_;
  assign new_n29503_ = ~new_n29499_ & new_n29502_;
  assign new_n29504_ = ~new_n29419_ & ~new_n29503_;
  assign new_n29505_ = \b[8]  & ~new_n29397_;
  assign new_n29506_ = ~new_n29395_ & new_n29505_;
  assign new_n29507_ = ~new_n29410_ & ~new_n29506_;
  assign new_n29508_ = ~new_n29504_ & new_n29507_;
  assign new_n29509_ = ~new_n29410_ & ~new_n29508_;
  assign new_n29510_ = \b[9]  & ~new_n29407_;
  assign new_n29511_ = ~new_n29405_ & new_n29510_;
  assign new_n29512_ = ~new_n29409_ & ~new_n29511_;
  assign new_n29513_ = ~new_n29509_ & new_n29512_;
  assign new_n29514_ = ~new_n29409_ & ~new_n29513_;
  assign new_n29515_ = new_n1145_ & ~new_n29514_;
  assign new_n29516_ = ~new_n29398_ & ~new_n29515_;
  assign new_n29517_ = ~new_n29419_ & new_n29507_;
  assign new_n29518_ = ~new_n29503_ & new_n29517_;
  assign new_n29519_ = ~new_n29504_ & ~new_n29507_;
  assign new_n29520_ = ~new_n29518_ & ~new_n29519_;
  assign new_n29521_ = new_n1145_ & ~new_n29520_;
  assign new_n29522_ = ~new_n29514_ & new_n29521_;
  assign new_n29523_ = ~new_n29516_ & ~new_n29522_;
  assign new_n29524_ = ~new_n29408_ & ~new_n29515_;
  assign new_n29525_ = ~new_n29410_ & new_n29512_;
  assign new_n29526_ = ~new_n29508_ & new_n29525_;
  assign new_n29527_ = ~new_n29509_ & ~new_n29512_;
  assign new_n29528_ = ~new_n29526_ & ~new_n29527_;
  assign new_n29529_ = new_n29515_ & ~new_n29528_;
  assign new_n29530_ = ~new_n29524_ & ~new_n29529_;
  assign new_n29531_ = ~\b[10]  & ~new_n29530_;
  assign new_n29532_ = ~\b[9]  & ~new_n29523_;
  assign new_n29533_ = ~new_n29418_ & ~new_n29515_;
  assign new_n29534_ = ~new_n29428_ & new_n29502_;
  assign new_n29535_ = ~new_n29498_ & new_n29534_;
  assign new_n29536_ = ~new_n29499_ & ~new_n29502_;
  assign new_n29537_ = ~new_n29535_ & ~new_n29536_;
  assign new_n29538_ = new_n1145_ & ~new_n29537_;
  assign new_n29539_ = ~new_n29514_ & new_n29538_;
  assign new_n29540_ = ~new_n29533_ & ~new_n29539_;
  assign new_n29541_ = ~\b[8]  & ~new_n29540_;
  assign new_n29542_ = ~new_n29427_ & ~new_n29515_;
  assign new_n29543_ = ~new_n29437_ & new_n29497_;
  assign new_n29544_ = ~new_n29493_ & new_n29543_;
  assign new_n29545_ = ~new_n29494_ & ~new_n29497_;
  assign new_n29546_ = ~new_n29544_ & ~new_n29545_;
  assign new_n29547_ = new_n1145_ & ~new_n29546_;
  assign new_n29548_ = ~new_n29514_ & new_n29547_;
  assign new_n29549_ = ~new_n29542_ & ~new_n29548_;
  assign new_n29550_ = ~\b[7]  & ~new_n29549_;
  assign new_n29551_ = ~new_n29436_ & ~new_n29515_;
  assign new_n29552_ = ~new_n29446_ & new_n29492_;
  assign new_n29553_ = ~new_n29488_ & new_n29552_;
  assign new_n29554_ = ~new_n29489_ & ~new_n29492_;
  assign new_n29555_ = ~new_n29553_ & ~new_n29554_;
  assign new_n29556_ = new_n1145_ & ~new_n29555_;
  assign new_n29557_ = ~new_n29514_ & new_n29556_;
  assign new_n29558_ = ~new_n29551_ & ~new_n29557_;
  assign new_n29559_ = ~\b[6]  & ~new_n29558_;
  assign new_n29560_ = ~new_n29445_ & ~new_n29515_;
  assign new_n29561_ = ~new_n29455_ & new_n29487_;
  assign new_n29562_ = ~new_n29483_ & new_n29561_;
  assign new_n29563_ = ~new_n29484_ & ~new_n29487_;
  assign new_n29564_ = ~new_n29562_ & ~new_n29563_;
  assign new_n29565_ = new_n1145_ & ~new_n29564_;
  assign new_n29566_ = ~new_n29514_ & new_n29565_;
  assign new_n29567_ = ~new_n29560_ & ~new_n29566_;
  assign new_n29568_ = ~\b[5]  & ~new_n29567_;
  assign new_n29569_ = ~new_n29454_ & ~new_n29515_;
  assign new_n29570_ = ~new_n29463_ & new_n29482_;
  assign new_n29571_ = ~new_n29478_ & new_n29570_;
  assign new_n29572_ = ~new_n29479_ & ~new_n29482_;
  assign new_n29573_ = ~new_n29571_ & ~new_n29572_;
  assign new_n29574_ = new_n1145_ & ~new_n29573_;
  assign new_n29575_ = ~new_n29514_ & new_n29574_;
  assign new_n29576_ = ~new_n29569_ & ~new_n29575_;
  assign new_n29577_ = ~\b[4]  & ~new_n29576_;
  assign new_n29578_ = ~new_n29462_ & ~new_n29515_;
  assign new_n29579_ = ~new_n29473_ & new_n29477_;
  assign new_n29580_ = ~new_n29472_ & new_n29579_;
  assign new_n29581_ = ~new_n29474_ & ~new_n29477_;
  assign new_n29582_ = ~new_n29580_ & ~new_n29581_;
  assign new_n29583_ = new_n1145_ & ~new_n29582_;
  assign new_n29584_ = ~new_n29514_ & new_n29583_;
  assign new_n29585_ = ~new_n29578_ & ~new_n29584_;
  assign new_n29586_ = ~\b[3]  & ~new_n29585_;
  assign new_n29587_ = ~new_n29467_ & ~new_n29515_;
  assign new_n29588_ = new_n1099_ & ~new_n29470_;
  assign new_n29589_ = ~new_n29468_ & new_n29588_;
  assign new_n29590_ = new_n1145_ & ~new_n29589_;
  assign new_n29591_ = ~new_n29472_ & new_n29590_;
  assign new_n29592_ = ~new_n29514_ & new_n29591_;
  assign new_n29593_ = ~new_n29587_ & ~new_n29592_;
  assign new_n29594_ = ~\b[2]  & ~new_n29593_;
  assign new_n29595_ = new_n1230_ & ~new_n29514_;
  assign new_n29596_ = \a[54]  & ~new_n29595_;
  assign new_n29597_ = new_n1236_ & ~new_n29514_;
  assign new_n29598_ = ~new_n29596_ & ~new_n29597_;
  assign new_n29599_ = \b[1]  & ~new_n29598_;
  assign new_n29600_ = ~\b[1]  & ~new_n29597_;
  assign new_n29601_ = ~new_n29596_ & new_n29600_;
  assign new_n29602_ = ~new_n29599_ & ~new_n29601_;
  assign new_n29603_ = ~new_n1243_ & ~new_n29602_;
  assign new_n29604_ = ~\b[1]  & ~new_n29598_;
  assign new_n29605_ = ~new_n29603_ & ~new_n29604_;
  assign new_n29606_ = \b[2]  & ~new_n29592_;
  assign new_n29607_ = ~new_n29587_ & new_n29606_;
  assign new_n29608_ = ~new_n29594_ & ~new_n29607_;
  assign new_n29609_ = ~new_n29605_ & new_n29608_;
  assign new_n29610_ = ~new_n29594_ & ~new_n29609_;
  assign new_n29611_ = \b[3]  & ~new_n29584_;
  assign new_n29612_ = ~new_n29578_ & new_n29611_;
  assign new_n29613_ = ~new_n29586_ & ~new_n29612_;
  assign new_n29614_ = ~new_n29610_ & new_n29613_;
  assign new_n29615_ = ~new_n29586_ & ~new_n29614_;
  assign new_n29616_ = \b[4]  & ~new_n29575_;
  assign new_n29617_ = ~new_n29569_ & new_n29616_;
  assign new_n29618_ = ~new_n29577_ & ~new_n29617_;
  assign new_n29619_ = ~new_n29615_ & new_n29618_;
  assign new_n29620_ = ~new_n29577_ & ~new_n29619_;
  assign new_n29621_ = \b[5]  & ~new_n29566_;
  assign new_n29622_ = ~new_n29560_ & new_n29621_;
  assign new_n29623_ = ~new_n29568_ & ~new_n29622_;
  assign new_n29624_ = ~new_n29620_ & new_n29623_;
  assign new_n29625_ = ~new_n29568_ & ~new_n29624_;
  assign new_n29626_ = \b[6]  & ~new_n29557_;
  assign new_n29627_ = ~new_n29551_ & new_n29626_;
  assign new_n29628_ = ~new_n29559_ & ~new_n29627_;
  assign new_n29629_ = ~new_n29625_ & new_n29628_;
  assign new_n29630_ = ~new_n29559_ & ~new_n29629_;
  assign new_n29631_ = \b[7]  & ~new_n29548_;
  assign new_n29632_ = ~new_n29542_ & new_n29631_;
  assign new_n29633_ = ~new_n29550_ & ~new_n29632_;
  assign new_n29634_ = ~new_n29630_ & new_n29633_;
  assign new_n29635_ = ~new_n29550_ & ~new_n29634_;
  assign new_n29636_ = \b[8]  & ~new_n29539_;
  assign new_n29637_ = ~new_n29533_ & new_n29636_;
  assign new_n29638_ = ~new_n29541_ & ~new_n29637_;
  assign new_n29639_ = ~new_n29635_ & new_n29638_;
  assign new_n29640_ = ~new_n29541_ & ~new_n29639_;
  assign new_n29641_ = \b[9]  & ~new_n29522_;
  assign new_n29642_ = ~new_n29516_ & new_n29641_;
  assign new_n29643_ = ~new_n29532_ & ~new_n29642_;
  assign new_n29644_ = ~new_n29640_ & new_n29643_;
  assign new_n29645_ = ~new_n29532_ & ~new_n29644_;
  assign new_n29646_ = \b[10]  & ~new_n29524_;
  assign new_n29647_ = ~new_n29529_ & new_n29646_;
  assign new_n29648_ = ~new_n29531_ & ~new_n29647_;
  assign new_n29649_ = ~new_n29645_ & new_n29648_;
  assign new_n29650_ = ~new_n29531_ & ~new_n29649_;
  assign new_n29651_ = new_n1294_ & ~new_n29650_;
  assign new_n29652_ = ~new_n29523_ & ~new_n29651_;
  assign new_n29653_ = ~new_n29541_ & new_n29643_;
  assign new_n29654_ = ~new_n29639_ & new_n29653_;
  assign new_n29655_ = ~new_n29640_ & ~new_n29643_;
  assign new_n29656_ = ~new_n29654_ & ~new_n29655_;
  assign new_n29657_ = new_n1294_ & ~new_n29656_;
  assign new_n29658_ = ~new_n29650_ & new_n29657_;
  assign new_n29659_ = ~new_n29652_ & ~new_n29658_;
  assign new_n29660_ = ~\b[10]  & ~new_n29659_;
  assign new_n29661_ = ~new_n29540_ & ~new_n29651_;
  assign new_n29662_ = ~new_n29550_ & new_n29638_;
  assign new_n29663_ = ~new_n29634_ & new_n29662_;
  assign new_n29664_ = ~new_n29635_ & ~new_n29638_;
  assign new_n29665_ = ~new_n29663_ & ~new_n29664_;
  assign new_n29666_ = new_n1294_ & ~new_n29665_;
  assign new_n29667_ = ~new_n29650_ & new_n29666_;
  assign new_n29668_ = ~new_n29661_ & ~new_n29667_;
  assign new_n29669_ = ~\b[9]  & ~new_n29668_;
  assign new_n29670_ = ~new_n29549_ & ~new_n29651_;
  assign new_n29671_ = ~new_n29559_ & new_n29633_;
  assign new_n29672_ = ~new_n29629_ & new_n29671_;
  assign new_n29673_ = ~new_n29630_ & ~new_n29633_;
  assign new_n29674_ = ~new_n29672_ & ~new_n29673_;
  assign new_n29675_ = new_n1294_ & ~new_n29674_;
  assign new_n29676_ = ~new_n29650_ & new_n29675_;
  assign new_n29677_ = ~new_n29670_ & ~new_n29676_;
  assign new_n29678_ = ~\b[8]  & ~new_n29677_;
  assign new_n29679_ = ~new_n29558_ & ~new_n29651_;
  assign new_n29680_ = ~new_n29568_ & new_n29628_;
  assign new_n29681_ = ~new_n29624_ & new_n29680_;
  assign new_n29682_ = ~new_n29625_ & ~new_n29628_;
  assign new_n29683_ = ~new_n29681_ & ~new_n29682_;
  assign new_n29684_ = new_n1294_ & ~new_n29683_;
  assign new_n29685_ = ~new_n29650_ & new_n29684_;
  assign new_n29686_ = ~new_n29679_ & ~new_n29685_;
  assign new_n29687_ = ~\b[7]  & ~new_n29686_;
  assign new_n29688_ = ~new_n29567_ & ~new_n29651_;
  assign new_n29689_ = ~new_n29577_ & new_n29623_;
  assign new_n29690_ = ~new_n29619_ & new_n29689_;
  assign new_n29691_ = ~new_n29620_ & ~new_n29623_;
  assign new_n29692_ = ~new_n29690_ & ~new_n29691_;
  assign new_n29693_ = new_n1294_ & ~new_n29692_;
  assign new_n29694_ = ~new_n29650_ & new_n29693_;
  assign new_n29695_ = ~new_n29688_ & ~new_n29694_;
  assign new_n29696_ = ~\b[6]  & ~new_n29695_;
  assign new_n29697_ = ~new_n29576_ & ~new_n29651_;
  assign new_n29698_ = ~new_n29586_ & new_n29618_;
  assign new_n29699_ = ~new_n29614_ & new_n29698_;
  assign new_n29700_ = ~new_n29615_ & ~new_n29618_;
  assign new_n29701_ = ~new_n29699_ & ~new_n29700_;
  assign new_n29702_ = new_n1294_ & ~new_n29701_;
  assign new_n29703_ = ~new_n29650_ & new_n29702_;
  assign new_n29704_ = ~new_n29697_ & ~new_n29703_;
  assign new_n29705_ = ~\b[5]  & ~new_n29704_;
  assign new_n29706_ = ~new_n29585_ & ~new_n29651_;
  assign new_n29707_ = ~new_n29594_ & new_n29613_;
  assign new_n29708_ = ~new_n29609_ & new_n29707_;
  assign new_n29709_ = ~new_n29610_ & ~new_n29613_;
  assign new_n29710_ = ~new_n29708_ & ~new_n29709_;
  assign new_n29711_ = new_n1294_ & ~new_n29710_;
  assign new_n29712_ = ~new_n29650_ & new_n29711_;
  assign new_n29713_ = ~new_n29706_ & ~new_n29712_;
  assign new_n29714_ = ~\b[4]  & ~new_n29713_;
  assign new_n29715_ = ~new_n29593_ & ~new_n29651_;
  assign new_n29716_ = ~new_n29604_ & new_n29608_;
  assign new_n29717_ = ~new_n29603_ & new_n29716_;
  assign new_n29718_ = ~new_n29605_ & ~new_n29608_;
  assign new_n29719_ = ~new_n29717_ & ~new_n29718_;
  assign new_n29720_ = new_n1294_ & ~new_n29719_;
  assign new_n29721_ = ~new_n29650_ & new_n29720_;
  assign new_n29722_ = ~new_n29715_ & ~new_n29721_;
  assign new_n29723_ = ~\b[3]  & ~new_n29722_;
  assign new_n29724_ = ~new_n29598_ & ~new_n29651_;
  assign new_n29725_ = new_n1243_ & ~new_n29601_;
  assign new_n29726_ = ~new_n29599_ & new_n29725_;
  assign new_n29727_ = new_n1294_ & ~new_n29726_;
  assign new_n29728_ = ~new_n29603_ & new_n29727_;
  assign new_n29729_ = ~new_n29650_ & new_n29728_;
  assign new_n29730_ = ~new_n29724_ & ~new_n29729_;
  assign new_n29731_ = ~\b[2]  & ~new_n29730_;
  assign new_n29732_ = new_n1379_ & ~new_n29650_;
  assign new_n29733_ = \a[53]  & ~new_n29732_;
  assign new_n29734_ = new_n1385_ & ~new_n29650_;
  assign new_n29735_ = ~new_n29733_ & ~new_n29734_;
  assign new_n29736_ = \b[1]  & ~new_n29735_;
  assign new_n29737_ = ~\b[1]  & ~new_n29734_;
  assign new_n29738_ = ~new_n29733_ & new_n29737_;
  assign new_n29739_ = ~new_n29736_ & ~new_n29738_;
  assign new_n29740_ = ~new_n1392_ & ~new_n29739_;
  assign new_n29741_ = ~\b[1]  & ~new_n29735_;
  assign new_n29742_ = ~new_n29740_ & ~new_n29741_;
  assign new_n29743_ = \b[2]  & ~new_n29729_;
  assign new_n29744_ = ~new_n29724_ & new_n29743_;
  assign new_n29745_ = ~new_n29731_ & ~new_n29744_;
  assign new_n29746_ = ~new_n29742_ & new_n29745_;
  assign new_n29747_ = ~new_n29731_ & ~new_n29746_;
  assign new_n29748_ = \b[3]  & ~new_n29721_;
  assign new_n29749_ = ~new_n29715_ & new_n29748_;
  assign new_n29750_ = ~new_n29723_ & ~new_n29749_;
  assign new_n29751_ = ~new_n29747_ & new_n29750_;
  assign new_n29752_ = ~new_n29723_ & ~new_n29751_;
  assign new_n29753_ = \b[4]  & ~new_n29712_;
  assign new_n29754_ = ~new_n29706_ & new_n29753_;
  assign new_n29755_ = ~new_n29714_ & ~new_n29754_;
  assign new_n29756_ = ~new_n29752_ & new_n29755_;
  assign new_n29757_ = ~new_n29714_ & ~new_n29756_;
  assign new_n29758_ = \b[5]  & ~new_n29703_;
  assign new_n29759_ = ~new_n29697_ & new_n29758_;
  assign new_n29760_ = ~new_n29705_ & ~new_n29759_;
  assign new_n29761_ = ~new_n29757_ & new_n29760_;
  assign new_n29762_ = ~new_n29705_ & ~new_n29761_;
  assign new_n29763_ = \b[6]  & ~new_n29694_;
  assign new_n29764_ = ~new_n29688_ & new_n29763_;
  assign new_n29765_ = ~new_n29696_ & ~new_n29764_;
  assign new_n29766_ = ~new_n29762_ & new_n29765_;
  assign new_n29767_ = ~new_n29696_ & ~new_n29766_;
  assign new_n29768_ = \b[7]  & ~new_n29685_;
  assign new_n29769_ = ~new_n29679_ & new_n29768_;
  assign new_n29770_ = ~new_n29687_ & ~new_n29769_;
  assign new_n29771_ = ~new_n29767_ & new_n29770_;
  assign new_n29772_ = ~new_n29687_ & ~new_n29771_;
  assign new_n29773_ = \b[8]  & ~new_n29676_;
  assign new_n29774_ = ~new_n29670_ & new_n29773_;
  assign new_n29775_ = ~new_n29678_ & ~new_n29774_;
  assign new_n29776_ = ~new_n29772_ & new_n29775_;
  assign new_n29777_ = ~new_n29678_ & ~new_n29776_;
  assign new_n29778_ = \b[9]  & ~new_n29667_;
  assign new_n29779_ = ~new_n29661_ & new_n29778_;
  assign new_n29780_ = ~new_n29669_ & ~new_n29779_;
  assign new_n29781_ = ~new_n29777_ & new_n29780_;
  assign new_n29782_ = ~new_n29669_ & ~new_n29781_;
  assign new_n29783_ = \b[10]  & ~new_n29658_;
  assign new_n29784_ = ~new_n29652_ & new_n29783_;
  assign new_n29785_ = ~new_n29660_ & ~new_n29784_;
  assign new_n29786_ = ~new_n29782_ & new_n29785_;
  assign new_n29787_ = ~new_n29660_ & ~new_n29786_;
  assign new_n29788_ = ~new_n29530_ & ~new_n29651_;
  assign new_n29789_ = ~new_n29532_ & new_n29648_;
  assign new_n29790_ = ~new_n29644_ & new_n29789_;
  assign new_n29791_ = ~new_n29645_ & ~new_n29648_;
  assign new_n29792_ = ~new_n29790_ & ~new_n29791_;
  assign new_n29793_ = new_n29651_ & ~new_n29792_;
  assign new_n29794_ = ~new_n29788_ & ~new_n29793_;
  assign new_n29795_ = ~\b[11]  & ~new_n29794_;
  assign new_n29796_ = \b[11]  & ~new_n29788_;
  assign new_n29797_ = ~new_n29793_ & new_n29796_;
  assign new_n29798_ = new_n1452_ & ~new_n29797_;
  assign new_n29799_ = ~new_n29795_ & new_n29798_;
  assign new_n29800_ = ~new_n29787_ & new_n29799_;
  assign new_n29801_ = new_n1294_ & ~new_n29794_;
  assign new_n29802_ = ~new_n29800_ & ~new_n29801_;
  assign new_n29803_ = ~new_n29669_ & new_n29785_;
  assign new_n29804_ = ~new_n29781_ & new_n29803_;
  assign new_n29805_ = ~new_n29782_ & ~new_n29785_;
  assign new_n29806_ = ~new_n29804_ & ~new_n29805_;
  assign new_n29807_ = ~new_n29802_ & ~new_n29806_;
  assign new_n29808_ = ~new_n29659_ & ~new_n29801_;
  assign new_n29809_ = ~new_n29800_ & new_n29808_;
  assign new_n29810_ = ~new_n29807_ & ~new_n29809_;
  assign new_n29811_ = ~new_n29660_ & ~new_n29797_;
  assign new_n29812_ = ~new_n29795_ & new_n29811_;
  assign new_n29813_ = ~new_n29786_ & new_n29812_;
  assign new_n29814_ = ~new_n29795_ & ~new_n29797_;
  assign new_n29815_ = ~new_n29787_ & ~new_n29814_;
  assign new_n29816_ = ~new_n29813_ & ~new_n29815_;
  assign new_n29817_ = ~new_n29802_ & ~new_n29816_;
  assign new_n29818_ = ~new_n29794_ & ~new_n29801_;
  assign new_n29819_ = ~new_n29800_ & new_n29818_;
  assign new_n29820_ = ~new_n29817_ & ~new_n29819_;
  assign new_n29821_ = ~\b[12]  & ~new_n29820_;
  assign new_n29822_ = ~\b[11]  & ~new_n29810_;
  assign new_n29823_ = ~new_n29678_ & new_n29780_;
  assign new_n29824_ = ~new_n29776_ & new_n29823_;
  assign new_n29825_ = ~new_n29777_ & ~new_n29780_;
  assign new_n29826_ = ~new_n29824_ & ~new_n29825_;
  assign new_n29827_ = ~new_n29802_ & ~new_n29826_;
  assign new_n29828_ = ~new_n29668_ & ~new_n29801_;
  assign new_n29829_ = ~new_n29800_ & new_n29828_;
  assign new_n29830_ = ~new_n29827_ & ~new_n29829_;
  assign new_n29831_ = ~\b[10]  & ~new_n29830_;
  assign new_n29832_ = ~new_n29687_ & new_n29775_;
  assign new_n29833_ = ~new_n29771_ & new_n29832_;
  assign new_n29834_ = ~new_n29772_ & ~new_n29775_;
  assign new_n29835_ = ~new_n29833_ & ~new_n29834_;
  assign new_n29836_ = ~new_n29802_ & ~new_n29835_;
  assign new_n29837_ = ~new_n29677_ & ~new_n29801_;
  assign new_n29838_ = ~new_n29800_ & new_n29837_;
  assign new_n29839_ = ~new_n29836_ & ~new_n29838_;
  assign new_n29840_ = ~\b[9]  & ~new_n29839_;
  assign new_n29841_ = ~new_n29696_ & new_n29770_;
  assign new_n29842_ = ~new_n29766_ & new_n29841_;
  assign new_n29843_ = ~new_n29767_ & ~new_n29770_;
  assign new_n29844_ = ~new_n29842_ & ~new_n29843_;
  assign new_n29845_ = ~new_n29802_ & ~new_n29844_;
  assign new_n29846_ = ~new_n29686_ & ~new_n29801_;
  assign new_n29847_ = ~new_n29800_ & new_n29846_;
  assign new_n29848_ = ~new_n29845_ & ~new_n29847_;
  assign new_n29849_ = ~\b[8]  & ~new_n29848_;
  assign new_n29850_ = ~new_n29705_ & new_n29765_;
  assign new_n29851_ = ~new_n29761_ & new_n29850_;
  assign new_n29852_ = ~new_n29762_ & ~new_n29765_;
  assign new_n29853_ = ~new_n29851_ & ~new_n29852_;
  assign new_n29854_ = ~new_n29802_ & ~new_n29853_;
  assign new_n29855_ = ~new_n29695_ & ~new_n29801_;
  assign new_n29856_ = ~new_n29800_ & new_n29855_;
  assign new_n29857_ = ~new_n29854_ & ~new_n29856_;
  assign new_n29858_ = ~\b[7]  & ~new_n29857_;
  assign new_n29859_ = ~new_n29714_ & new_n29760_;
  assign new_n29860_ = ~new_n29756_ & new_n29859_;
  assign new_n29861_ = ~new_n29757_ & ~new_n29760_;
  assign new_n29862_ = ~new_n29860_ & ~new_n29861_;
  assign new_n29863_ = ~new_n29802_ & ~new_n29862_;
  assign new_n29864_ = ~new_n29704_ & ~new_n29801_;
  assign new_n29865_ = ~new_n29800_ & new_n29864_;
  assign new_n29866_ = ~new_n29863_ & ~new_n29865_;
  assign new_n29867_ = ~\b[6]  & ~new_n29866_;
  assign new_n29868_ = ~new_n29723_ & new_n29755_;
  assign new_n29869_ = ~new_n29751_ & new_n29868_;
  assign new_n29870_ = ~new_n29752_ & ~new_n29755_;
  assign new_n29871_ = ~new_n29869_ & ~new_n29870_;
  assign new_n29872_ = ~new_n29802_ & ~new_n29871_;
  assign new_n29873_ = ~new_n29713_ & ~new_n29801_;
  assign new_n29874_ = ~new_n29800_ & new_n29873_;
  assign new_n29875_ = ~new_n29872_ & ~new_n29874_;
  assign new_n29876_ = ~\b[5]  & ~new_n29875_;
  assign new_n29877_ = ~new_n29731_ & new_n29750_;
  assign new_n29878_ = ~new_n29746_ & new_n29877_;
  assign new_n29879_ = ~new_n29747_ & ~new_n29750_;
  assign new_n29880_ = ~new_n29878_ & ~new_n29879_;
  assign new_n29881_ = ~new_n29802_ & ~new_n29880_;
  assign new_n29882_ = ~new_n29722_ & ~new_n29801_;
  assign new_n29883_ = ~new_n29800_ & new_n29882_;
  assign new_n29884_ = ~new_n29881_ & ~new_n29883_;
  assign new_n29885_ = ~\b[4]  & ~new_n29884_;
  assign new_n29886_ = ~new_n29741_ & new_n29745_;
  assign new_n29887_ = ~new_n29740_ & new_n29886_;
  assign new_n29888_ = ~new_n29742_ & ~new_n29745_;
  assign new_n29889_ = ~new_n29887_ & ~new_n29888_;
  assign new_n29890_ = ~new_n29802_ & ~new_n29889_;
  assign new_n29891_ = ~new_n29730_ & ~new_n29801_;
  assign new_n29892_ = ~new_n29800_ & new_n29891_;
  assign new_n29893_ = ~new_n29890_ & ~new_n29892_;
  assign new_n29894_ = ~\b[3]  & ~new_n29893_;
  assign new_n29895_ = new_n1392_ & ~new_n29738_;
  assign new_n29896_ = ~new_n29736_ & new_n29895_;
  assign new_n29897_ = ~new_n29740_ & ~new_n29896_;
  assign new_n29898_ = ~new_n29802_ & new_n29897_;
  assign new_n29899_ = ~new_n29735_ & ~new_n29801_;
  assign new_n29900_ = ~new_n29800_ & new_n29899_;
  assign new_n29901_ = ~new_n29898_ & ~new_n29900_;
  assign new_n29902_ = ~\b[2]  & ~new_n29901_;
  assign new_n29903_ = \b[0]  & ~new_n29802_;
  assign new_n29904_ = \a[52]  & ~new_n29903_;
  assign new_n29905_ = new_n1392_ & ~new_n29802_;
  assign new_n29906_ = ~new_n29904_ & ~new_n29905_;
  assign new_n29907_ = \b[1]  & ~new_n29906_;
  assign new_n29908_ = ~\b[1]  & ~new_n29905_;
  assign new_n29909_ = ~new_n29904_ & new_n29908_;
  assign new_n29910_ = ~new_n29907_ & ~new_n29909_;
  assign new_n29911_ = ~new_n1566_ & ~new_n29910_;
  assign new_n29912_ = ~\b[1]  & ~new_n29906_;
  assign new_n29913_ = ~new_n29911_ & ~new_n29912_;
  assign new_n29914_ = \b[2]  & ~new_n29900_;
  assign new_n29915_ = ~new_n29898_ & new_n29914_;
  assign new_n29916_ = ~new_n29902_ & ~new_n29915_;
  assign new_n29917_ = ~new_n29913_ & new_n29916_;
  assign new_n29918_ = ~new_n29902_ & ~new_n29917_;
  assign new_n29919_ = \b[3]  & ~new_n29892_;
  assign new_n29920_ = ~new_n29890_ & new_n29919_;
  assign new_n29921_ = ~new_n29894_ & ~new_n29920_;
  assign new_n29922_ = ~new_n29918_ & new_n29921_;
  assign new_n29923_ = ~new_n29894_ & ~new_n29922_;
  assign new_n29924_ = \b[4]  & ~new_n29883_;
  assign new_n29925_ = ~new_n29881_ & new_n29924_;
  assign new_n29926_ = ~new_n29885_ & ~new_n29925_;
  assign new_n29927_ = ~new_n29923_ & new_n29926_;
  assign new_n29928_ = ~new_n29885_ & ~new_n29927_;
  assign new_n29929_ = \b[5]  & ~new_n29874_;
  assign new_n29930_ = ~new_n29872_ & new_n29929_;
  assign new_n29931_ = ~new_n29876_ & ~new_n29930_;
  assign new_n29932_ = ~new_n29928_ & new_n29931_;
  assign new_n29933_ = ~new_n29876_ & ~new_n29932_;
  assign new_n29934_ = \b[6]  & ~new_n29865_;
  assign new_n29935_ = ~new_n29863_ & new_n29934_;
  assign new_n29936_ = ~new_n29867_ & ~new_n29935_;
  assign new_n29937_ = ~new_n29933_ & new_n29936_;
  assign new_n29938_ = ~new_n29867_ & ~new_n29937_;
  assign new_n29939_ = \b[7]  & ~new_n29856_;
  assign new_n29940_ = ~new_n29854_ & new_n29939_;
  assign new_n29941_ = ~new_n29858_ & ~new_n29940_;
  assign new_n29942_ = ~new_n29938_ & new_n29941_;
  assign new_n29943_ = ~new_n29858_ & ~new_n29942_;
  assign new_n29944_ = \b[8]  & ~new_n29847_;
  assign new_n29945_ = ~new_n29845_ & new_n29944_;
  assign new_n29946_ = ~new_n29849_ & ~new_n29945_;
  assign new_n29947_ = ~new_n29943_ & new_n29946_;
  assign new_n29948_ = ~new_n29849_ & ~new_n29947_;
  assign new_n29949_ = \b[9]  & ~new_n29838_;
  assign new_n29950_ = ~new_n29836_ & new_n29949_;
  assign new_n29951_ = ~new_n29840_ & ~new_n29950_;
  assign new_n29952_ = ~new_n29948_ & new_n29951_;
  assign new_n29953_ = ~new_n29840_ & ~new_n29952_;
  assign new_n29954_ = \b[10]  & ~new_n29829_;
  assign new_n29955_ = ~new_n29827_ & new_n29954_;
  assign new_n29956_ = ~new_n29831_ & ~new_n29955_;
  assign new_n29957_ = ~new_n29953_ & new_n29956_;
  assign new_n29958_ = ~new_n29831_ & ~new_n29957_;
  assign new_n29959_ = \b[11]  & ~new_n29809_;
  assign new_n29960_ = ~new_n29807_ & new_n29959_;
  assign new_n29961_ = ~new_n29822_ & ~new_n29960_;
  assign new_n29962_ = ~new_n29958_ & new_n29961_;
  assign new_n29963_ = ~new_n29822_ & ~new_n29962_;
  assign new_n29964_ = \b[12]  & ~new_n29819_;
  assign new_n29965_ = ~new_n29817_ & new_n29964_;
  assign new_n29966_ = ~new_n29821_ & ~new_n29965_;
  assign new_n29967_ = ~new_n29963_ & new_n29966_;
  assign new_n29968_ = ~new_n29821_ & ~new_n29967_;
  assign new_n29969_ = new_n1626_ & ~new_n29968_;
  assign new_n29970_ = ~new_n29810_ & ~new_n29969_;
  assign new_n29971_ = ~new_n29831_ & new_n29961_;
  assign new_n29972_ = ~new_n29957_ & new_n29971_;
  assign new_n29973_ = ~new_n29958_ & ~new_n29961_;
  assign new_n29974_ = ~new_n29972_ & ~new_n29973_;
  assign new_n29975_ = new_n1626_ & ~new_n29974_;
  assign new_n29976_ = ~new_n29968_ & new_n29975_;
  assign new_n29977_ = ~new_n29970_ & ~new_n29976_;
  assign new_n29978_ = ~new_n29820_ & ~new_n29969_;
  assign new_n29979_ = ~new_n29822_ & new_n29966_;
  assign new_n29980_ = ~new_n29962_ & new_n29979_;
  assign new_n29981_ = ~new_n29963_ & ~new_n29966_;
  assign new_n29982_ = ~new_n29980_ & ~new_n29981_;
  assign new_n29983_ = new_n29969_ & ~new_n29982_;
  assign new_n29984_ = ~new_n29978_ & ~new_n29983_;
  assign new_n29985_ = ~\b[13]  & ~new_n29984_;
  assign new_n29986_ = ~\b[12]  & ~new_n29977_;
  assign new_n29987_ = ~new_n29830_ & ~new_n29969_;
  assign new_n29988_ = ~new_n29840_ & new_n29956_;
  assign new_n29989_ = ~new_n29952_ & new_n29988_;
  assign new_n29990_ = ~new_n29953_ & ~new_n29956_;
  assign new_n29991_ = ~new_n29989_ & ~new_n29990_;
  assign new_n29992_ = new_n1626_ & ~new_n29991_;
  assign new_n29993_ = ~new_n29968_ & new_n29992_;
  assign new_n29994_ = ~new_n29987_ & ~new_n29993_;
  assign new_n29995_ = ~\b[11]  & ~new_n29994_;
  assign new_n29996_ = ~new_n29839_ & ~new_n29969_;
  assign new_n29997_ = ~new_n29849_ & new_n29951_;
  assign new_n29998_ = ~new_n29947_ & new_n29997_;
  assign new_n29999_ = ~new_n29948_ & ~new_n29951_;
  assign new_n30000_ = ~new_n29998_ & ~new_n29999_;
  assign new_n30001_ = new_n1626_ & ~new_n30000_;
  assign new_n30002_ = ~new_n29968_ & new_n30001_;
  assign new_n30003_ = ~new_n29996_ & ~new_n30002_;
  assign new_n30004_ = ~\b[10]  & ~new_n30003_;
  assign new_n30005_ = ~new_n29848_ & ~new_n29969_;
  assign new_n30006_ = ~new_n29858_ & new_n29946_;
  assign new_n30007_ = ~new_n29942_ & new_n30006_;
  assign new_n30008_ = ~new_n29943_ & ~new_n29946_;
  assign new_n30009_ = ~new_n30007_ & ~new_n30008_;
  assign new_n30010_ = new_n1626_ & ~new_n30009_;
  assign new_n30011_ = ~new_n29968_ & new_n30010_;
  assign new_n30012_ = ~new_n30005_ & ~new_n30011_;
  assign new_n30013_ = ~\b[9]  & ~new_n30012_;
  assign new_n30014_ = ~new_n29857_ & ~new_n29969_;
  assign new_n30015_ = ~new_n29867_ & new_n29941_;
  assign new_n30016_ = ~new_n29937_ & new_n30015_;
  assign new_n30017_ = ~new_n29938_ & ~new_n29941_;
  assign new_n30018_ = ~new_n30016_ & ~new_n30017_;
  assign new_n30019_ = new_n1626_ & ~new_n30018_;
  assign new_n30020_ = ~new_n29968_ & new_n30019_;
  assign new_n30021_ = ~new_n30014_ & ~new_n30020_;
  assign new_n30022_ = ~\b[8]  & ~new_n30021_;
  assign new_n30023_ = ~new_n29866_ & ~new_n29969_;
  assign new_n30024_ = ~new_n29876_ & new_n29936_;
  assign new_n30025_ = ~new_n29932_ & new_n30024_;
  assign new_n30026_ = ~new_n29933_ & ~new_n29936_;
  assign new_n30027_ = ~new_n30025_ & ~new_n30026_;
  assign new_n30028_ = new_n1626_ & ~new_n30027_;
  assign new_n30029_ = ~new_n29968_ & new_n30028_;
  assign new_n30030_ = ~new_n30023_ & ~new_n30029_;
  assign new_n30031_ = ~\b[7]  & ~new_n30030_;
  assign new_n30032_ = ~new_n29875_ & ~new_n29969_;
  assign new_n30033_ = ~new_n29885_ & new_n29931_;
  assign new_n30034_ = ~new_n29927_ & new_n30033_;
  assign new_n30035_ = ~new_n29928_ & ~new_n29931_;
  assign new_n30036_ = ~new_n30034_ & ~new_n30035_;
  assign new_n30037_ = new_n1626_ & ~new_n30036_;
  assign new_n30038_ = ~new_n29968_ & new_n30037_;
  assign new_n30039_ = ~new_n30032_ & ~new_n30038_;
  assign new_n30040_ = ~\b[6]  & ~new_n30039_;
  assign new_n30041_ = ~new_n29884_ & ~new_n29969_;
  assign new_n30042_ = ~new_n29894_ & new_n29926_;
  assign new_n30043_ = ~new_n29922_ & new_n30042_;
  assign new_n30044_ = ~new_n29923_ & ~new_n29926_;
  assign new_n30045_ = ~new_n30043_ & ~new_n30044_;
  assign new_n30046_ = new_n1626_ & ~new_n30045_;
  assign new_n30047_ = ~new_n29968_ & new_n30046_;
  assign new_n30048_ = ~new_n30041_ & ~new_n30047_;
  assign new_n30049_ = ~\b[5]  & ~new_n30048_;
  assign new_n30050_ = ~new_n29893_ & ~new_n29969_;
  assign new_n30051_ = ~new_n29902_ & new_n29921_;
  assign new_n30052_ = ~new_n29917_ & new_n30051_;
  assign new_n30053_ = ~new_n29918_ & ~new_n29921_;
  assign new_n30054_ = ~new_n30052_ & ~new_n30053_;
  assign new_n30055_ = new_n1626_ & ~new_n30054_;
  assign new_n30056_ = ~new_n29968_ & new_n30055_;
  assign new_n30057_ = ~new_n30050_ & ~new_n30056_;
  assign new_n30058_ = ~\b[4]  & ~new_n30057_;
  assign new_n30059_ = ~new_n29901_ & ~new_n29969_;
  assign new_n30060_ = ~new_n29912_ & new_n29916_;
  assign new_n30061_ = ~new_n29911_ & new_n30060_;
  assign new_n30062_ = ~new_n29913_ & ~new_n29916_;
  assign new_n30063_ = ~new_n30061_ & ~new_n30062_;
  assign new_n30064_ = new_n1626_ & ~new_n30063_;
  assign new_n30065_ = ~new_n29968_ & new_n30064_;
  assign new_n30066_ = ~new_n30059_ & ~new_n30065_;
  assign new_n30067_ = ~\b[3]  & ~new_n30066_;
  assign new_n30068_ = ~new_n29906_ & ~new_n29969_;
  assign new_n30069_ = new_n1566_ & ~new_n29909_;
  assign new_n30070_ = ~new_n29907_ & new_n30069_;
  assign new_n30071_ = new_n1626_ & ~new_n30070_;
  assign new_n30072_ = ~new_n29911_ & new_n30071_;
  assign new_n30073_ = ~new_n29968_ & new_n30072_;
  assign new_n30074_ = ~new_n30068_ & ~new_n30073_;
  assign new_n30075_ = ~\b[2]  & ~new_n30074_;
  assign new_n30076_ = new_n1738_ & ~new_n29968_;
  assign new_n30077_ = \a[51]  & ~new_n30076_;
  assign new_n30078_ = new_n1743_ & ~new_n29968_;
  assign new_n30079_ = ~new_n30077_ & ~new_n30078_;
  assign new_n30080_ = \b[1]  & ~new_n30079_;
  assign new_n30081_ = ~\b[1]  & ~new_n30078_;
  assign new_n30082_ = ~new_n30077_ & new_n30081_;
  assign new_n30083_ = ~new_n30080_ & ~new_n30082_;
  assign new_n30084_ = ~new_n1750_ & ~new_n30083_;
  assign new_n30085_ = ~\b[1]  & ~new_n30079_;
  assign new_n30086_ = ~new_n30084_ & ~new_n30085_;
  assign new_n30087_ = \b[2]  & ~new_n30073_;
  assign new_n30088_ = ~new_n30068_ & new_n30087_;
  assign new_n30089_ = ~new_n30075_ & ~new_n30088_;
  assign new_n30090_ = ~new_n30086_ & new_n30089_;
  assign new_n30091_ = ~new_n30075_ & ~new_n30090_;
  assign new_n30092_ = \b[3]  & ~new_n30065_;
  assign new_n30093_ = ~new_n30059_ & new_n30092_;
  assign new_n30094_ = ~new_n30067_ & ~new_n30093_;
  assign new_n30095_ = ~new_n30091_ & new_n30094_;
  assign new_n30096_ = ~new_n30067_ & ~new_n30095_;
  assign new_n30097_ = \b[4]  & ~new_n30056_;
  assign new_n30098_ = ~new_n30050_ & new_n30097_;
  assign new_n30099_ = ~new_n30058_ & ~new_n30098_;
  assign new_n30100_ = ~new_n30096_ & new_n30099_;
  assign new_n30101_ = ~new_n30058_ & ~new_n30100_;
  assign new_n30102_ = \b[5]  & ~new_n30047_;
  assign new_n30103_ = ~new_n30041_ & new_n30102_;
  assign new_n30104_ = ~new_n30049_ & ~new_n30103_;
  assign new_n30105_ = ~new_n30101_ & new_n30104_;
  assign new_n30106_ = ~new_n30049_ & ~new_n30105_;
  assign new_n30107_ = \b[6]  & ~new_n30038_;
  assign new_n30108_ = ~new_n30032_ & new_n30107_;
  assign new_n30109_ = ~new_n30040_ & ~new_n30108_;
  assign new_n30110_ = ~new_n30106_ & new_n30109_;
  assign new_n30111_ = ~new_n30040_ & ~new_n30110_;
  assign new_n30112_ = \b[7]  & ~new_n30029_;
  assign new_n30113_ = ~new_n30023_ & new_n30112_;
  assign new_n30114_ = ~new_n30031_ & ~new_n30113_;
  assign new_n30115_ = ~new_n30111_ & new_n30114_;
  assign new_n30116_ = ~new_n30031_ & ~new_n30115_;
  assign new_n30117_ = \b[8]  & ~new_n30020_;
  assign new_n30118_ = ~new_n30014_ & new_n30117_;
  assign new_n30119_ = ~new_n30022_ & ~new_n30118_;
  assign new_n30120_ = ~new_n30116_ & new_n30119_;
  assign new_n30121_ = ~new_n30022_ & ~new_n30120_;
  assign new_n30122_ = \b[9]  & ~new_n30011_;
  assign new_n30123_ = ~new_n30005_ & new_n30122_;
  assign new_n30124_ = ~new_n30013_ & ~new_n30123_;
  assign new_n30125_ = ~new_n30121_ & new_n30124_;
  assign new_n30126_ = ~new_n30013_ & ~new_n30125_;
  assign new_n30127_ = \b[10]  & ~new_n30002_;
  assign new_n30128_ = ~new_n29996_ & new_n30127_;
  assign new_n30129_ = ~new_n30004_ & ~new_n30128_;
  assign new_n30130_ = ~new_n30126_ & new_n30129_;
  assign new_n30131_ = ~new_n30004_ & ~new_n30130_;
  assign new_n30132_ = \b[11]  & ~new_n29993_;
  assign new_n30133_ = ~new_n29987_ & new_n30132_;
  assign new_n30134_ = ~new_n29995_ & ~new_n30133_;
  assign new_n30135_ = ~new_n30131_ & new_n30134_;
  assign new_n30136_ = ~new_n29995_ & ~new_n30135_;
  assign new_n30137_ = \b[12]  & ~new_n29976_;
  assign new_n30138_ = ~new_n29970_ & new_n30137_;
  assign new_n30139_ = ~new_n29986_ & ~new_n30138_;
  assign new_n30140_ = ~new_n30136_ & new_n30139_;
  assign new_n30141_ = ~new_n29986_ & ~new_n30140_;
  assign new_n30142_ = \b[13]  & ~new_n29978_;
  assign new_n30143_ = ~new_n29983_ & new_n30142_;
  assign new_n30144_ = ~new_n29985_ & ~new_n30143_;
  assign new_n30145_ = ~new_n30141_ & new_n30144_;
  assign new_n30146_ = ~new_n29985_ & ~new_n30145_;
  assign new_n30147_ = new_n1816_ & ~new_n30146_;
  assign new_n30148_ = ~new_n29977_ & ~new_n30147_;
  assign new_n30149_ = ~new_n29995_ & new_n30139_;
  assign new_n30150_ = ~new_n30135_ & new_n30149_;
  assign new_n30151_ = ~new_n30136_ & ~new_n30139_;
  assign new_n30152_ = ~new_n30150_ & ~new_n30151_;
  assign new_n30153_ = new_n1816_ & ~new_n30152_;
  assign new_n30154_ = ~new_n30146_ & new_n30153_;
  assign new_n30155_ = ~new_n30148_ & ~new_n30154_;
  assign new_n30156_ = ~\b[13]  & ~new_n30155_;
  assign new_n30157_ = ~new_n29994_ & ~new_n30147_;
  assign new_n30158_ = ~new_n30004_ & new_n30134_;
  assign new_n30159_ = ~new_n30130_ & new_n30158_;
  assign new_n30160_ = ~new_n30131_ & ~new_n30134_;
  assign new_n30161_ = ~new_n30159_ & ~new_n30160_;
  assign new_n30162_ = new_n1816_ & ~new_n30161_;
  assign new_n30163_ = ~new_n30146_ & new_n30162_;
  assign new_n30164_ = ~new_n30157_ & ~new_n30163_;
  assign new_n30165_ = ~\b[12]  & ~new_n30164_;
  assign new_n30166_ = ~new_n30003_ & ~new_n30147_;
  assign new_n30167_ = ~new_n30013_ & new_n30129_;
  assign new_n30168_ = ~new_n30125_ & new_n30167_;
  assign new_n30169_ = ~new_n30126_ & ~new_n30129_;
  assign new_n30170_ = ~new_n30168_ & ~new_n30169_;
  assign new_n30171_ = new_n1816_ & ~new_n30170_;
  assign new_n30172_ = ~new_n30146_ & new_n30171_;
  assign new_n30173_ = ~new_n30166_ & ~new_n30172_;
  assign new_n30174_ = ~\b[11]  & ~new_n30173_;
  assign new_n30175_ = ~new_n30012_ & ~new_n30147_;
  assign new_n30176_ = ~new_n30022_ & new_n30124_;
  assign new_n30177_ = ~new_n30120_ & new_n30176_;
  assign new_n30178_ = ~new_n30121_ & ~new_n30124_;
  assign new_n30179_ = ~new_n30177_ & ~new_n30178_;
  assign new_n30180_ = new_n1816_ & ~new_n30179_;
  assign new_n30181_ = ~new_n30146_ & new_n30180_;
  assign new_n30182_ = ~new_n30175_ & ~new_n30181_;
  assign new_n30183_ = ~\b[10]  & ~new_n30182_;
  assign new_n30184_ = ~new_n30021_ & ~new_n30147_;
  assign new_n30185_ = ~new_n30031_ & new_n30119_;
  assign new_n30186_ = ~new_n30115_ & new_n30185_;
  assign new_n30187_ = ~new_n30116_ & ~new_n30119_;
  assign new_n30188_ = ~new_n30186_ & ~new_n30187_;
  assign new_n30189_ = new_n1816_ & ~new_n30188_;
  assign new_n30190_ = ~new_n30146_ & new_n30189_;
  assign new_n30191_ = ~new_n30184_ & ~new_n30190_;
  assign new_n30192_ = ~\b[9]  & ~new_n30191_;
  assign new_n30193_ = ~new_n30030_ & ~new_n30147_;
  assign new_n30194_ = ~new_n30040_ & new_n30114_;
  assign new_n30195_ = ~new_n30110_ & new_n30194_;
  assign new_n30196_ = ~new_n30111_ & ~new_n30114_;
  assign new_n30197_ = ~new_n30195_ & ~new_n30196_;
  assign new_n30198_ = new_n1816_ & ~new_n30197_;
  assign new_n30199_ = ~new_n30146_ & new_n30198_;
  assign new_n30200_ = ~new_n30193_ & ~new_n30199_;
  assign new_n30201_ = ~\b[8]  & ~new_n30200_;
  assign new_n30202_ = ~new_n30039_ & ~new_n30147_;
  assign new_n30203_ = ~new_n30049_ & new_n30109_;
  assign new_n30204_ = ~new_n30105_ & new_n30203_;
  assign new_n30205_ = ~new_n30106_ & ~new_n30109_;
  assign new_n30206_ = ~new_n30204_ & ~new_n30205_;
  assign new_n30207_ = new_n1816_ & ~new_n30206_;
  assign new_n30208_ = ~new_n30146_ & new_n30207_;
  assign new_n30209_ = ~new_n30202_ & ~new_n30208_;
  assign new_n30210_ = ~\b[7]  & ~new_n30209_;
  assign new_n30211_ = ~new_n30048_ & ~new_n30147_;
  assign new_n30212_ = ~new_n30058_ & new_n30104_;
  assign new_n30213_ = ~new_n30100_ & new_n30212_;
  assign new_n30214_ = ~new_n30101_ & ~new_n30104_;
  assign new_n30215_ = ~new_n30213_ & ~new_n30214_;
  assign new_n30216_ = new_n1816_ & ~new_n30215_;
  assign new_n30217_ = ~new_n30146_ & new_n30216_;
  assign new_n30218_ = ~new_n30211_ & ~new_n30217_;
  assign new_n30219_ = ~\b[6]  & ~new_n30218_;
  assign new_n30220_ = ~new_n30057_ & ~new_n30147_;
  assign new_n30221_ = ~new_n30067_ & new_n30099_;
  assign new_n30222_ = ~new_n30095_ & new_n30221_;
  assign new_n30223_ = ~new_n30096_ & ~new_n30099_;
  assign new_n30224_ = ~new_n30222_ & ~new_n30223_;
  assign new_n30225_ = new_n1816_ & ~new_n30224_;
  assign new_n30226_ = ~new_n30146_ & new_n30225_;
  assign new_n30227_ = ~new_n30220_ & ~new_n30226_;
  assign new_n30228_ = ~\b[5]  & ~new_n30227_;
  assign new_n30229_ = ~new_n30066_ & ~new_n30147_;
  assign new_n30230_ = ~new_n30075_ & new_n30094_;
  assign new_n30231_ = ~new_n30090_ & new_n30230_;
  assign new_n30232_ = ~new_n30091_ & ~new_n30094_;
  assign new_n30233_ = ~new_n30231_ & ~new_n30232_;
  assign new_n30234_ = new_n1816_ & ~new_n30233_;
  assign new_n30235_ = ~new_n30146_ & new_n30234_;
  assign new_n30236_ = ~new_n30229_ & ~new_n30235_;
  assign new_n30237_ = ~\b[4]  & ~new_n30236_;
  assign new_n30238_ = ~new_n30074_ & ~new_n30147_;
  assign new_n30239_ = ~new_n30085_ & new_n30089_;
  assign new_n30240_ = ~new_n30084_ & new_n30239_;
  assign new_n30241_ = ~new_n30086_ & ~new_n30089_;
  assign new_n30242_ = ~new_n30240_ & ~new_n30241_;
  assign new_n30243_ = new_n1816_ & ~new_n30242_;
  assign new_n30244_ = ~new_n30146_ & new_n30243_;
  assign new_n30245_ = ~new_n30238_ & ~new_n30244_;
  assign new_n30246_ = ~\b[3]  & ~new_n30245_;
  assign new_n30247_ = ~new_n30079_ & ~new_n30147_;
  assign new_n30248_ = new_n1750_ & ~new_n30082_;
  assign new_n30249_ = ~new_n30080_ & new_n30248_;
  assign new_n30250_ = new_n1816_ & ~new_n30249_;
  assign new_n30251_ = ~new_n30084_ & new_n30250_;
  assign new_n30252_ = ~new_n30146_ & new_n30251_;
  assign new_n30253_ = ~new_n30247_ & ~new_n30252_;
  assign new_n30254_ = ~\b[2]  & ~new_n30253_;
  assign new_n30255_ = new_n1929_ & ~new_n30146_;
  assign new_n30256_ = \a[50]  & ~new_n30255_;
  assign new_n30257_ = new_n1935_ & ~new_n30146_;
  assign new_n30258_ = ~new_n30256_ & ~new_n30257_;
  assign new_n30259_ = \b[1]  & ~new_n30258_;
  assign new_n30260_ = ~\b[1]  & ~new_n30257_;
  assign new_n30261_ = ~new_n30256_ & new_n30260_;
  assign new_n30262_ = ~new_n30259_ & ~new_n30261_;
  assign new_n30263_ = ~new_n1942_ & ~new_n30262_;
  assign new_n30264_ = ~\b[1]  & ~new_n30258_;
  assign new_n30265_ = ~new_n30263_ & ~new_n30264_;
  assign new_n30266_ = \b[2]  & ~new_n30252_;
  assign new_n30267_ = ~new_n30247_ & new_n30266_;
  assign new_n30268_ = ~new_n30254_ & ~new_n30267_;
  assign new_n30269_ = ~new_n30265_ & new_n30268_;
  assign new_n30270_ = ~new_n30254_ & ~new_n30269_;
  assign new_n30271_ = \b[3]  & ~new_n30244_;
  assign new_n30272_ = ~new_n30238_ & new_n30271_;
  assign new_n30273_ = ~new_n30246_ & ~new_n30272_;
  assign new_n30274_ = ~new_n30270_ & new_n30273_;
  assign new_n30275_ = ~new_n30246_ & ~new_n30274_;
  assign new_n30276_ = \b[4]  & ~new_n30235_;
  assign new_n30277_ = ~new_n30229_ & new_n30276_;
  assign new_n30278_ = ~new_n30237_ & ~new_n30277_;
  assign new_n30279_ = ~new_n30275_ & new_n30278_;
  assign new_n30280_ = ~new_n30237_ & ~new_n30279_;
  assign new_n30281_ = \b[5]  & ~new_n30226_;
  assign new_n30282_ = ~new_n30220_ & new_n30281_;
  assign new_n30283_ = ~new_n30228_ & ~new_n30282_;
  assign new_n30284_ = ~new_n30280_ & new_n30283_;
  assign new_n30285_ = ~new_n30228_ & ~new_n30284_;
  assign new_n30286_ = \b[6]  & ~new_n30217_;
  assign new_n30287_ = ~new_n30211_ & new_n30286_;
  assign new_n30288_ = ~new_n30219_ & ~new_n30287_;
  assign new_n30289_ = ~new_n30285_ & new_n30288_;
  assign new_n30290_ = ~new_n30219_ & ~new_n30289_;
  assign new_n30291_ = \b[7]  & ~new_n30208_;
  assign new_n30292_ = ~new_n30202_ & new_n30291_;
  assign new_n30293_ = ~new_n30210_ & ~new_n30292_;
  assign new_n30294_ = ~new_n30290_ & new_n30293_;
  assign new_n30295_ = ~new_n30210_ & ~new_n30294_;
  assign new_n30296_ = \b[8]  & ~new_n30199_;
  assign new_n30297_ = ~new_n30193_ & new_n30296_;
  assign new_n30298_ = ~new_n30201_ & ~new_n30297_;
  assign new_n30299_ = ~new_n30295_ & new_n30298_;
  assign new_n30300_ = ~new_n30201_ & ~new_n30299_;
  assign new_n30301_ = \b[9]  & ~new_n30190_;
  assign new_n30302_ = ~new_n30184_ & new_n30301_;
  assign new_n30303_ = ~new_n30192_ & ~new_n30302_;
  assign new_n30304_ = ~new_n30300_ & new_n30303_;
  assign new_n30305_ = ~new_n30192_ & ~new_n30304_;
  assign new_n30306_ = \b[10]  & ~new_n30181_;
  assign new_n30307_ = ~new_n30175_ & new_n30306_;
  assign new_n30308_ = ~new_n30183_ & ~new_n30307_;
  assign new_n30309_ = ~new_n30305_ & new_n30308_;
  assign new_n30310_ = ~new_n30183_ & ~new_n30309_;
  assign new_n30311_ = \b[11]  & ~new_n30172_;
  assign new_n30312_ = ~new_n30166_ & new_n30311_;
  assign new_n30313_ = ~new_n30174_ & ~new_n30312_;
  assign new_n30314_ = ~new_n30310_ & new_n30313_;
  assign new_n30315_ = ~new_n30174_ & ~new_n30314_;
  assign new_n30316_ = \b[12]  & ~new_n30163_;
  assign new_n30317_ = ~new_n30157_ & new_n30316_;
  assign new_n30318_ = ~new_n30165_ & ~new_n30317_;
  assign new_n30319_ = ~new_n30315_ & new_n30318_;
  assign new_n30320_ = ~new_n30165_ & ~new_n30319_;
  assign new_n30321_ = \b[13]  & ~new_n30154_;
  assign new_n30322_ = ~new_n30148_ & new_n30321_;
  assign new_n30323_ = ~new_n30156_ & ~new_n30322_;
  assign new_n30324_ = ~new_n30320_ & new_n30323_;
  assign new_n30325_ = ~new_n30156_ & ~new_n30324_;
  assign new_n30326_ = ~new_n29984_ & ~new_n30147_;
  assign new_n30327_ = ~new_n29986_ & new_n30144_;
  assign new_n30328_ = ~new_n30140_ & new_n30327_;
  assign new_n30329_ = ~new_n30141_ & ~new_n30144_;
  assign new_n30330_ = ~new_n30328_ & ~new_n30329_;
  assign new_n30331_ = new_n30147_ & ~new_n30330_;
  assign new_n30332_ = ~new_n30326_ & ~new_n30331_;
  assign new_n30333_ = ~\b[14]  & ~new_n30332_;
  assign new_n30334_ = \b[14]  & ~new_n30326_;
  assign new_n30335_ = ~new_n30331_ & new_n30334_;
  assign new_n30336_ = new_n2018_ & ~new_n30335_;
  assign new_n30337_ = ~new_n30333_ & new_n30336_;
  assign new_n30338_ = ~new_n30325_ & new_n30337_;
  assign new_n30339_ = new_n1816_ & ~new_n30332_;
  assign new_n30340_ = ~new_n30338_ & ~new_n30339_;
  assign new_n30341_ = ~new_n30165_ & new_n30323_;
  assign new_n30342_ = ~new_n30319_ & new_n30341_;
  assign new_n30343_ = ~new_n30320_ & ~new_n30323_;
  assign new_n30344_ = ~new_n30342_ & ~new_n30343_;
  assign new_n30345_ = ~new_n30340_ & ~new_n30344_;
  assign new_n30346_ = ~new_n30155_ & ~new_n30339_;
  assign new_n30347_ = ~new_n30338_ & new_n30346_;
  assign new_n30348_ = ~new_n30345_ & ~new_n30347_;
  assign new_n30349_ = ~new_n30156_ & ~new_n30335_;
  assign new_n30350_ = ~new_n30333_ & new_n30349_;
  assign new_n30351_ = ~new_n30324_ & new_n30350_;
  assign new_n30352_ = ~new_n30333_ & ~new_n30335_;
  assign new_n30353_ = ~new_n30325_ & ~new_n30352_;
  assign new_n30354_ = ~new_n30351_ & ~new_n30353_;
  assign new_n30355_ = ~new_n30340_ & ~new_n30354_;
  assign new_n30356_ = ~new_n30332_ & ~new_n30339_;
  assign new_n30357_ = ~new_n30338_ & new_n30356_;
  assign new_n30358_ = ~new_n30355_ & ~new_n30357_;
  assign new_n30359_ = ~\b[15]  & ~new_n30358_;
  assign new_n30360_ = ~\b[14]  & ~new_n30348_;
  assign new_n30361_ = ~new_n30174_ & new_n30318_;
  assign new_n30362_ = ~new_n30314_ & new_n30361_;
  assign new_n30363_ = ~new_n30315_ & ~new_n30318_;
  assign new_n30364_ = ~new_n30362_ & ~new_n30363_;
  assign new_n30365_ = ~new_n30340_ & ~new_n30364_;
  assign new_n30366_ = ~new_n30164_ & ~new_n30339_;
  assign new_n30367_ = ~new_n30338_ & new_n30366_;
  assign new_n30368_ = ~new_n30365_ & ~new_n30367_;
  assign new_n30369_ = ~\b[13]  & ~new_n30368_;
  assign new_n30370_ = ~new_n30183_ & new_n30313_;
  assign new_n30371_ = ~new_n30309_ & new_n30370_;
  assign new_n30372_ = ~new_n30310_ & ~new_n30313_;
  assign new_n30373_ = ~new_n30371_ & ~new_n30372_;
  assign new_n30374_ = ~new_n30340_ & ~new_n30373_;
  assign new_n30375_ = ~new_n30173_ & ~new_n30339_;
  assign new_n30376_ = ~new_n30338_ & new_n30375_;
  assign new_n30377_ = ~new_n30374_ & ~new_n30376_;
  assign new_n30378_ = ~\b[12]  & ~new_n30377_;
  assign new_n30379_ = ~new_n30192_ & new_n30308_;
  assign new_n30380_ = ~new_n30304_ & new_n30379_;
  assign new_n30381_ = ~new_n30305_ & ~new_n30308_;
  assign new_n30382_ = ~new_n30380_ & ~new_n30381_;
  assign new_n30383_ = ~new_n30340_ & ~new_n30382_;
  assign new_n30384_ = ~new_n30182_ & ~new_n30339_;
  assign new_n30385_ = ~new_n30338_ & new_n30384_;
  assign new_n30386_ = ~new_n30383_ & ~new_n30385_;
  assign new_n30387_ = ~\b[11]  & ~new_n30386_;
  assign new_n30388_ = ~new_n30201_ & new_n30303_;
  assign new_n30389_ = ~new_n30299_ & new_n30388_;
  assign new_n30390_ = ~new_n30300_ & ~new_n30303_;
  assign new_n30391_ = ~new_n30389_ & ~new_n30390_;
  assign new_n30392_ = ~new_n30340_ & ~new_n30391_;
  assign new_n30393_ = ~new_n30191_ & ~new_n30339_;
  assign new_n30394_ = ~new_n30338_ & new_n30393_;
  assign new_n30395_ = ~new_n30392_ & ~new_n30394_;
  assign new_n30396_ = ~\b[10]  & ~new_n30395_;
  assign new_n30397_ = ~new_n30210_ & new_n30298_;
  assign new_n30398_ = ~new_n30294_ & new_n30397_;
  assign new_n30399_ = ~new_n30295_ & ~new_n30298_;
  assign new_n30400_ = ~new_n30398_ & ~new_n30399_;
  assign new_n30401_ = ~new_n30340_ & ~new_n30400_;
  assign new_n30402_ = ~new_n30200_ & ~new_n30339_;
  assign new_n30403_ = ~new_n30338_ & new_n30402_;
  assign new_n30404_ = ~new_n30401_ & ~new_n30403_;
  assign new_n30405_ = ~\b[9]  & ~new_n30404_;
  assign new_n30406_ = ~new_n30219_ & new_n30293_;
  assign new_n30407_ = ~new_n30289_ & new_n30406_;
  assign new_n30408_ = ~new_n30290_ & ~new_n30293_;
  assign new_n30409_ = ~new_n30407_ & ~new_n30408_;
  assign new_n30410_ = ~new_n30340_ & ~new_n30409_;
  assign new_n30411_ = ~new_n30209_ & ~new_n30339_;
  assign new_n30412_ = ~new_n30338_ & new_n30411_;
  assign new_n30413_ = ~new_n30410_ & ~new_n30412_;
  assign new_n30414_ = ~\b[8]  & ~new_n30413_;
  assign new_n30415_ = ~new_n30228_ & new_n30288_;
  assign new_n30416_ = ~new_n30284_ & new_n30415_;
  assign new_n30417_ = ~new_n30285_ & ~new_n30288_;
  assign new_n30418_ = ~new_n30416_ & ~new_n30417_;
  assign new_n30419_ = ~new_n30340_ & ~new_n30418_;
  assign new_n30420_ = ~new_n30218_ & ~new_n30339_;
  assign new_n30421_ = ~new_n30338_ & new_n30420_;
  assign new_n30422_ = ~new_n30419_ & ~new_n30421_;
  assign new_n30423_ = ~\b[7]  & ~new_n30422_;
  assign new_n30424_ = ~new_n30237_ & new_n30283_;
  assign new_n30425_ = ~new_n30279_ & new_n30424_;
  assign new_n30426_ = ~new_n30280_ & ~new_n30283_;
  assign new_n30427_ = ~new_n30425_ & ~new_n30426_;
  assign new_n30428_ = ~new_n30340_ & ~new_n30427_;
  assign new_n30429_ = ~new_n30227_ & ~new_n30339_;
  assign new_n30430_ = ~new_n30338_ & new_n30429_;
  assign new_n30431_ = ~new_n30428_ & ~new_n30430_;
  assign new_n30432_ = ~\b[6]  & ~new_n30431_;
  assign new_n30433_ = ~new_n30246_ & new_n30278_;
  assign new_n30434_ = ~new_n30274_ & new_n30433_;
  assign new_n30435_ = ~new_n30275_ & ~new_n30278_;
  assign new_n30436_ = ~new_n30434_ & ~new_n30435_;
  assign new_n30437_ = ~new_n30340_ & ~new_n30436_;
  assign new_n30438_ = ~new_n30236_ & ~new_n30339_;
  assign new_n30439_ = ~new_n30338_ & new_n30438_;
  assign new_n30440_ = ~new_n30437_ & ~new_n30439_;
  assign new_n30441_ = ~\b[5]  & ~new_n30440_;
  assign new_n30442_ = ~new_n30254_ & new_n30273_;
  assign new_n30443_ = ~new_n30269_ & new_n30442_;
  assign new_n30444_ = ~new_n30270_ & ~new_n30273_;
  assign new_n30445_ = ~new_n30443_ & ~new_n30444_;
  assign new_n30446_ = ~new_n30340_ & ~new_n30445_;
  assign new_n30447_ = ~new_n30245_ & ~new_n30339_;
  assign new_n30448_ = ~new_n30338_ & new_n30447_;
  assign new_n30449_ = ~new_n30446_ & ~new_n30448_;
  assign new_n30450_ = ~\b[4]  & ~new_n30449_;
  assign new_n30451_ = ~new_n30264_ & new_n30268_;
  assign new_n30452_ = ~new_n30263_ & new_n30451_;
  assign new_n30453_ = ~new_n30265_ & ~new_n30268_;
  assign new_n30454_ = ~new_n30452_ & ~new_n30453_;
  assign new_n30455_ = ~new_n30340_ & ~new_n30454_;
  assign new_n30456_ = ~new_n30253_ & ~new_n30339_;
  assign new_n30457_ = ~new_n30338_ & new_n30456_;
  assign new_n30458_ = ~new_n30455_ & ~new_n30457_;
  assign new_n30459_ = ~\b[3]  & ~new_n30458_;
  assign new_n30460_ = new_n1942_ & ~new_n30261_;
  assign new_n30461_ = ~new_n30259_ & new_n30460_;
  assign new_n30462_ = ~new_n30263_ & ~new_n30461_;
  assign new_n30463_ = ~new_n30340_ & new_n30462_;
  assign new_n30464_ = ~new_n30258_ & ~new_n30339_;
  assign new_n30465_ = ~new_n30338_ & new_n30464_;
  assign new_n30466_ = ~new_n30463_ & ~new_n30465_;
  assign new_n30467_ = ~\b[2]  & ~new_n30466_;
  assign new_n30468_ = \b[0]  & ~new_n30340_;
  assign new_n30469_ = \a[49]  & ~new_n30468_;
  assign new_n30470_ = new_n1942_ & ~new_n30340_;
  assign new_n30471_ = ~new_n30469_ & ~new_n30470_;
  assign new_n30472_ = \b[1]  & ~new_n30471_;
  assign new_n30473_ = ~\b[1]  & ~new_n30470_;
  assign new_n30474_ = ~new_n30469_ & new_n30473_;
  assign new_n30475_ = ~new_n30472_ & ~new_n30474_;
  assign new_n30476_ = ~new_n2159_ & ~new_n30475_;
  assign new_n30477_ = ~\b[1]  & ~new_n30471_;
  assign new_n30478_ = ~new_n30476_ & ~new_n30477_;
  assign new_n30479_ = \b[2]  & ~new_n30465_;
  assign new_n30480_ = ~new_n30463_ & new_n30479_;
  assign new_n30481_ = ~new_n30467_ & ~new_n30480_;
  assign new_n30482_ = ~new_n30478_ & new_n30481_;
  assign new_n30483_ = ~new_n30467_ & ~new_n30482_;
  assign new_n30484_ = \b[3]  & ~new_n30457_;
  assign new_n30485_ = ~new_n30455_ & new_n30484_;
  assign new_n30486_ = ~new_n30459_ & ~new_n30485_;
  assign new_n30487_ = ~new_n30483_ & new_n30486_;
  assign new_n30488_ = ~new_n30459_ & ~new_n30487_;
  assign new_n30489_ = \b[4]  & ~new_n30448_;
  assign new_n30490_ = ~new_n30446_ & new_n30489_;
  assign new_n30491_ = ~new_n30450_ & ~new_n30490_;
  assign new_n30492_ = ~new_n30488_ & new_n30491_;
  assign new_n30493_ = ~new_n30450_ & ~new_n30492_;
  assign new_n30494_ = \b[5]  & ~new_n30439_;
  assign new_n30495_ = ~new_n30437_ & new_n30494_;
  assign new_n30496_ = ~new_n30441_ & ~new_n30495_;
  assign new_n30497_ = ~new_n30493_ & new_n30496_;
  assign new_n30498_ = ~new_n30441_ & ~new_n30497_;
  assign new_n30499_ = \b[6]  & ~new_n30430_;
  assign new_n30500_ = ~new_n30428_ & new_n30499_;
  assign new_n30501_ = ~new_n30432_ & ~new_n30500_;
  assign new_n30502_ = ~new_n30498_ & new_n30501_;
  assign new_n30503_ = ~new_n30432_ & ~new_n30502_;
  assign new_n30504_ = \b[7]  & ~new_n30421_;
  assign new_n30505_ = ~new_n30419_ & new_n30504_;
  assign new_n30506_ = ~new_n30423_ & ~new_n30505_;
  assign new_n30507_ = ~new_n30503_ & new_n30506_;
  assign new_n30508_ = ~new_n30423_ & ~new_n30507_;
  assign new_n30509_ = \b[8]  & ~new_n30412_;
  assign new_n30510_ = ~new_n30410_ & new_n30509_;
  assign new_n30511_ = ~new_n30414_ & ~new_n30510_;
  assign new_n30512_ = ~new_n30508_ & new_n30511_;
  assign new_n30513_ = ~new_n30414_ & ~new_n30512_;
  assign new_n30514_ = \b[9]  & ~new_n30403_;
  assign new_n30515_ = ~new_n30401_ & new_n30514_;
  assign new_n30516_ = ~new_n30405_ & ~new_n30515_;
  assign new_n30517_ = ~new_n30513_ & new_n30516_;
  assign new_n30518_ = ~new_n30405_ & ~new_n30517_;
  assign new_n30519_ = \b[10]  & ~new_n30394_;
  assign new_n30520_ = ~new_n30392_ & new_n30519_;
  assign new_n30521_ = ~new_n30396_ & ~new_n30520_;
  assign new_n30522_ = ~new_n30518_ & new_n30521_;
  assign new_n30523_ = ~new_n30396_ & ~new_n30522_;
  assign new_n30524_ = \b[11]  & ~new_n30385_;
  assign new_n30525_ = ~new_n30383_ & new_n30524_;
  assign new_n30526_ = ~new_n30387_ & ~new_n30525_;
  assign new_n30527_ = ~new_n30523_ & new_n30526_;
  assign new_n30528_ = ~new_n30387_ & ~new_n30527_;
  assign new_n30529_ = \b[12]  & ~new_n30376_;
  assign new_n30530_ = ~new_n30374_ & new_n30529_;
  assign new_n30531_ = ~new_n30378_ & ~new_n30530_;
  assign new_n30532_ = ~new_n30528_ & new_n30531_;
  assign new_n30533_ = ~new_n30378_ & ~new_n30532_;
  assign new_n30534_ = \b[13]  & ~new_n30367_;
  assign new_n30535_ = ~new_n30365_ & new_n30534_;
  assign new_n30536_ = ~new_n30369_ & ~new_n30535_;
  assign new_n30537_ = ~new_n30533_ & new_n30536_;
  assign new_n30538_ = ~new_n30369_ & ~new_n30537_;
  assign new_n30539_ = \b[14]  & ~new_n30347_;
  assign new_n30540_ = ~new_n30345_ & new_n30539_;
  assign new_n30541_ = ~new_n30360_ & ~new_n30540_;
  assign new_n30542_ = ~new_n30538_ & new_n30541_;
  assign new_n30543_ = ~new_n30360_ & ~new_n30542_;
  assign new_n30544_ = \b[15]  & ~new_n30357_;
  assign new_n30545_ = ~new_n30355_ & new_n30544_;
  assign new_n30546_ = ~new_n30359_ & ~new_n30545_;
  assign new_n30547_ = ~new_n30543_ & new_n30546_;
  assign new_n30548_ = ~new_n30359_ & ~new_n30547_;
  assign new_n30549_ = new_n346_ & ~new_n30548_;
  assign new_n30550_ = ~new_n30348_ & ~new_n30549_;
  assign new_n30551_ = ~new_n30369_ & new_n30541_;
  assign new_n30552_ = ~new_n30537_ & new_n30551_;
  assign new_n30553_ = ~new_n30538_ & ~new_n30541_;
  assign new_n30554_ = ~new_n30552_ & ~new_n30553_;
  assign new_n30555_ = new_n346_ & ~new_n30554_;
  assign new_n30556_ = ~new_n30548_ & new_n30555_;
  assign new_n30557_ = ~new_n30550_ & ~new_n30556_;
  assign new_n30558_ = ~new_n30358_ & ~new_n30549_;
  assign new_n30559_ = ~new_n30360_ & new_n30546_;
  assign new_n30560_ = ~new_n30542_ & new_n30559_;
  assign new_n30561_ = ~new_n30543_ & ~new_n30546_;
  assign new_n30562_ = ~new_n30560_ & ~new_n30561_;
  assign new_n30563_ = new_n30549_ & ~new_n30562_;
  assign new_n30564_ = ~new_n30558_ & ~new_n30563_;
  assign new_n30565_ = ~\b[16]  & ~new_n30564_;
  assign new_n30566_ = ~\b[15]  & ~new_n30557_;
  assign new_n30567_ = ~new_n30368_ & ~new_n30549_;
  assign new_n30568_ = ~new_n30378_ & new_n30536_;
  assign new_n30569_ = ~new_n30532_ & new_n30568_;
  assign new_n30570_ = ~new_n30533_ & ~new_n30536_;
  assign new_n30571_ = ~new_n30569_ & ~new_n30570_;
  assign new_n30572_ = new_n346_ & ~new_n30571_;
  assign new_n30573_ = ~new_n30548_ & new_n30572_;
  assign new_n30574_ = ~new_n30567_ & ~new_n30573_;
  assign new_n30575_ = ~\b[14]  & ~new_n30574_;
  assign new_n30576_ = ~new_n30377_ & ~new_n30549_;
  assign new_n30577_ = ~new_n30387_ & new_n30531_;
  assign new_n30578_ = ~new_n30527_ & new_n30577_;
  assign new_n30579_ = ~new_n30528_ & ~new_n30531_;
  assign new_n30580_ = ~new_n30578_ & ~new_n30579_;
  assign new_n30581_ = new_n346_ & ~new_n30580_;
  assign new_n30582_ = ~new_n30548_ & new_n30581_;
  assign new_n30583_ = ~new_n30576_ & ~new_n30582_;
  assign new_n30584_ = ~\b[13]  & ~new_n30583_;
  assign new_n30585_ = ~new_n30386_ & ~new_n30549_;
  assign new_n30586_ = ~new_n30396_ & new_n30526_;
  assign new_n30587_ = ~new_n30522_ & new_n30586_;
  assign new_n30588_ = ~new_n30523_ & ~new_n30526_;
  assign new_n30589_ = ~new_n30587_ & ~new_n30588_;
  assign new_n30590_ = new_n346_ & ~new_n30589_;
  assign new_n30591_ = ~new_n30548_ & new_n30590_;
  assign new_n30592_ = ~new_n30585_ & ~new_n30591_;
  assign new_n30593_ = ~\b[12]  & ~new_n30592_;
  assign new_n30594_ = ~new_n30395_ & ~new_n30549_;
  assign new_n30595_ = ~new_n30405_ & new_n30521_;
  assign new_n30596_ = ~new_n30517_ & new_n30595_;
  assign new_n30597_ = ~new_n30518_ & ~new_n30521_;
  assign new_n30598_ = ~new_n30596_ & ~new_n30597_;
  assign new_n30599_ = new_n346_ & ~new_n30598_;
  assign new_n30600_ = ~new_n30548_ & new_n30599_;
  assign new_n30601_ = ~new_n30594_ & ~new_n30600_;
  assign new_n30602_ = ~\b[11]  & ~new_n30601_;
  assign new_n30603_ = ~new_n30404_ & ~new_n30549_;
  assign new_n30604_ = ~new_n30414_ & new_n30516_;
  assign new_n30605_ = ~new_n30512_ & new_n30604_;
  assign new_n30606_ = ~new_n30513_ & ~new_n30516_;
  assign new_n30607_ = ~new_n30605_ & ~new_n30606_;
  assign new_n30608_ = new_n346_ & ~new_n30607_;
  assign new_n30609_ = ~new_n30548_ & new_n30608_;
  assign new_n30610_ = ~new_n30603_ & ~new_n30609_;
  assign new_n30611_ = ~\b[10]  & ~new_n30610_;
  assign new_n30612_ = ~new_n30413_ & ~new_n30549_;
  assign new_n30613_ = ~new_n30423_ & new_n30511_;
  assign new_n30614_ = ~new_n30507_ & new_n30613_;
  assign new_n30615_ = ~new_n30508_ & ~new_n30511_;
  assign new_n30616_ = ~new_n30614_ & ~new_n30615_;
  assign new_n30617_ = new_n346_ & ~new_n30616_;
  assign new_n30618_ = ~new_n30548_ & new_n30617_;
  assign new_n30619_ = ~new_n30612_ & ~new_n30618_;
  assign new_n30620_ = ~\b[9]  & ~new_n30619_;
  assign new_n30621_ = ~new_n30422_ & ~new_n30549_;
  assign new_n30622_ = ~new_n30432_ & new_n30506_;
  assign new_n30623_ = ~new_n30502_ & new_n30622_;
  assign new_n30624_ = ~new_n30503_ & ~new_n30506_;
  assign new_n30625_ = ~new_n30623_ & ~new_n30624_;
  assign new_n30626_ = new_n346_ & ~new_n30625_;
  assign new_n30627_ = ~new_n30548_ & new_n30626_;
  assign new_n30628_ = ~new_n30621_ & ~new_n30627_;
  assign new_n30629_ = ~\b[8]  & ~new_n30628_;
  assign new_n30630_ = ~new_n30431_ & ~new_n30549_;
  assign new_n30631_ = ~new_n30441_ & new_n30501_;
  assign new_n30632_ = ~new_n30497_ & new_n30631_;
  assign new_n30633_ = ~new_n30498_ & ~new_n30501_;
  assign new_n30634_ = ~new_n30632_ & ~new_n30633_;
  assign new_n30635_ = new_n346_ & ~new_n30634_;
  assign new_n30636_ = ~new_n30548_ & new_n30635_;
  assign new_n30637_ = ~new_n30630_ & ~new_n30636_;
  assign new_n30638_ = ~\b[7]  & ~new_n30637_;
  assign new_n30639_ = ~new_n30440_ & ~new_n30549_;
  assign new_n30640_ = ~new_n30450_ & new_n30496_;
  assign new_n30641_ = ~new_n30492_ & new_n30640_;
  assign new_n30642_ = ~new_n30493_ & ~new_n30496_;
  assign new_n30643_ = ~new_n30641_ & ~new_n30642_;
  assign new_n30644_ = new_n346_ & ~new_n30643_;
  assign new_n30645_ = ~new_n30548_ & new_n30644_;
  assign new_n30646_ = ~new_n30639_ & ~new_n30645_;
  assign new_n30647_ = ~\b[6]  & ~new_n30646_;
  assign new_n30648_ = ~new_n30449_ & ~new_n30549_;
  assign new_n30649_ = ~new_n30459_ & new_n30491_;
  assign new_n30650_ = ~new_n30487_ & new_n30649_;
  assign new_n30651_ = ~new_n30488_ & ~new_n30491_;
  assign new_n30652_ = ~new_n30650_ & ~new_n30651_;
  assign new_n30653_ = new_n346_ & ~new_n30652_;
  assign new_n30654_ = ~new_n30548_ & new_n30653_;
  assign new_n30655_ = ~new_n30648_ & ~new_n30654_;
  assign new_n30656_ = ~\b[5]  & ~new_n30655_;
  assign new_n30657_ = ~new_n30458_ & ~new_n30549_;
  assign new_n30658_ = ~new_n30467_ & new_n30486_;
  assign new_n30659_ = ~new_n30482_ & new_n30658_;
  assign new_n30660_ = ~new_n30483_ & ~new_n30486_;
  assign new_n30661_ = ~new_n30659_ & ~new_n30660_;
  assign new_n30662_ = new_n346_ & ~new_n30661_;
  assign new_n30663_ = ~new_n30548_ & new_n30662_;
  assign new_n30664_ = ~new_n30657_ & ~new_n30663_;
  assign new_n30665_ = ~\b[4]  & ~new_n30664_;
  assign new_n30666_ = ~new_n30466_ & ~new_n30549_;
  assign new_n30667_ = ~new_n30477_ & new_n30481_;
  assign new_n30668_ = ~new_n30476_ & new_n30667_;
  assign new_n30669_ = ~new_n30478_ & ~new_n30481_;
  assign new_n30670_ = ~new_n30668_ & ~new_n30669_;
  assign new_n30671_ = new_n346_ & ~new_n30670_;
  assign new_n30672_ = ~new_n30548_ & new_n30671_;
  assign new_n30673_ = ~new_n30666_ & ~new_n30672_;
  assign new_n30674_ = ~\b[3]  & ~new_n30673_;
  assign new_n30675_ = ~new_n30471_ & ~new_n30549_;
  assign new_n30676_ = new_n2159_ & ~new_n30474_;
  assign new_n30677_ = ~new_n30472_ & new_n30676_;
  assign new_n30678_ = new_n346_ & ~new_n30677_;
  assign new_n30679_ = ~new_n30476_ & new_n30678_;
  assign new_n30680_ = ~new_n30548_ & new_n30679_;
  assign new_n30681_ = ~new_n30675_ & ~new_n30680_;
  assign new_n30682_ = ~\b[2]  & ~new_n30681_;
  assign new_n30683_ = new_n2370_ & ~new_n30548_;
  assign new_n30684_ = \a[48]  & ~new_n30683_;
  assign new_n30685_ = new_n2375_ & ~new_n30548_;
  assign new_n30686_ = ~new_n30684_ & ~new_n30685_;
  assign new_n30687_ = \b[1]  & ~new_n30686_;
  assign new_n30688_ = ~\b[1]  & ~new_n30685_;
  assign new_n30689_ = ~new_n30684_ & new_n30688_;
  assign new_n30690_ = ~new_n30687_ & ~new_n30689_;
  assign new_n30691_ = ~new_n2382_ & ~new_n30690_;
  assign new_n30692_ = ~\b[1]  & ~new_n30686_;
  assign new_n30693_ = ~new_n30691_ & ~new_n30692_;
  assign new_n30694_ = \b[2]  & ~new_n30680_;
  assign new_n30695_ = ~new_n30675_ & new_n30694_;
  assign new_n30696_ = ~new_n30682_ & ~new_n30695_;
  assign new_n30697_ = ~new_n30693_ & new_n30696_;
  assign new_n30698_ = ~new_n30682_ & ~new_n30697_;
  assign new_n30699_ = \b[3]  & ~new_n30672_;
  assign new_n30700_ = ~new_n30666_ & new_n30699_;
  assign new_n30701_ = ~new_n30674_ & ~new_n30700_;
  assign new_n30702_ = ~new_n30698_ & new_n30701_;
  assign new_n30703_ = ~new_n30674_ & ~new_n30702_;
  assign new_n30704_ = \b[4]  & ~new_n30663_;
  assign new_n30705_ = ~new_n30657_ & new_n30704_;
  assign new_n30706_ = ~new_n30665_ & ~new_n30705_;
  assign new_n30707_ = ~new_n30703_ & new_n30706_;
  assign new_n30708_ = ~new_n30665_ & ~new_n30707_;
  assign new_n30709_ = \b[5]  & ~new_n30654_;
  assign new_n30710_ = ~new_n30648_ & new_n30709_;
  assign new_n30711_ = ~new_n30656_ & ~new_n30710_;
  assign new_n30712_ = ~new_n30708_ & new_n30711_;
  assign new_n30713_ = ~new_n30656_ & ~new_n30712_;
  assign new_n30714_ = \b[6]  & ~new_n30645_;
  assign new_n30715_ = ~new_n30639_ & new_n30714_;
  assign new_n30716_ = ~new_n30647_ & ~new_n30715_;
  assign new_n30717_ = ~new_n30713_ & new_n30716_;
  assign new_n30718_ = ~new_n30647_ & ~new_n30717_;
  assign new_n30719_ = \b[7]  & ~new_n30636_;
  assign new_n30720_ = ~new_n30630_ & new_n30719_;
  assign new_n30721_ = ~new_n30638_ & ~new_n30720_;
  assign new_n30722_ = ~new_n30718_ & new_n30721_;
  assign new_n30723_ = ~new_n30638_ & ~new_n30722_;
  assign new_n30724_ = \b[8]  & ~new_n30627_;
  assign new_n30725_ = ~new_n30621_ & new_n30724_;
  assign new_n30726_ = ~new_n30629_ & ~new_n30725_;
  assign new_n30727_ = ~new_n30723_ & new_n30726_;
  assign new_n30728_ = ~new_n30629_ & ~new_n30727_;
  assign new_n30729_ = \b[9]  & ~new_n30618_;
  assign new_n30730_ = ~new_n30612_ & new_n30729_;
  assign new_n30731_ = ~new_n30620_ & ~new_n30730_;
  assign new_n30732_ = ~new_n30728_ & new_n30731_;
  assign new_n30733_ = ~new_n30620_ & ~new_n30732_;
  assign new_n30734_ = \b[10]  & ~new_n30609_;
  assign new_n30735_ = ~new_n30603_ & new_n30734_;
  assign new_n30736_ = ~new_n30611_ & ~new_n30735_;
  assign new_n30737_ = ~new_n30733_ & new_n30736_;
  assign new_n30738_ = ~new_n30611_ & ~new_n30737_;
  assign new_n30739_ = \b[11]  & ~new_n30600_;
  assign new_n30740_ = ~new_n30594_ & new_n30739_;
  assign new_n30741_ = ~new_n30602_ & ~new_n30740_;
  assign new_n30742_ = ~new_n30738_ & new_n30741_;
  assign new_n30743_ = ~new_n30602_ & ~new_n30742_;
  assign new_n30744_ = \b[12]  & ~new_n30591_;
  assign new_n30745_ = ~new_n30585_ & new_n30744_;
  assign new_n30746_ = ~new_n30593_ & ~new_n30745_;
  assign new_n30747_ = ~new_n30743_ & new_n30746_;
  assign new_n30748_ = ~new_n30593_ & ~new_n30747_;
  assign new_n30749_ = \b[13]  & ~new_n30582_;
  assign new_n30750_ = ~new_n30576_ & new_n30749_;
  assign new_n30751_ = ~new_n30584_ & ~new_n30750_;
  assign new_n30752_ = ~new_n30748_ & new_n30751_;
  assign new_n30753_ = ~new_n30584_ & ~new_n30752_;
  assign new_n30754_ = \b[14]  & ~new_n30573_;
  assign new_n30755_ = ~new_n30567_ & new_n30754_;
  assign new_n30756_ = ~new_n30575_ & ~new_n30755_;
  assign new_n30757_ = ~new_n30753_ & new_n30756_;
  assign new_n30758_ = ~new_n30575_ & ~new_n30757_;
  assign new_n30759_ = \b[15]  & ~new_n30556_;
  assign new_n30760_ = ~new_n30550_ & new_n30759_;
  assign new_n30761_ = ~new_n30566_ & ~new_n30760_;
  assign new_n30762_ = ~new_n30758_ & new_n30761_;
  assign new_n30763_ = ~new_n30566_ & ~new_n30762_;
  assign new_n30764_ = \b[16]  & ~new_n30558_;
  assign new_n30765_ = ~new_n30563_ & new_n30764_;
  assign new_n30766_ = ~new_n30565_ & ~new_n30765_;
  assign new_n30767_ = ~new_n30763_ & new_n30766_;
  assign new_n30768_ = ~new_n30565_ & ~new_n30767_;
  assign new_n30769_ = new_n475_ & ~new_n30768_;
  assign new_n30770_ = ~new_n30557_ & ~new_n30769_;
  assign new_n30771_ = ~new_n30575_ & new_n30761_;
  assign new_n30772_ = ~new_n30757_ & new_n30771_;
  assign new_n30773_ = ~new_n30758_ & ~new_n30761_;
  assign new_n30774_ = ~new_n30772_ & ~new_n30773_;
  assign new_n30775_ = new_n475_ & ~new_n30774_;
  assign new_n30776_ = ~new_n30768_ & new_n30775_;
  assign new_n30777_ = ~new_n30770_ & ~new_n30776_;
  assign new_n30778_ = ~\b[16]  & ~new_n30777_;
  assign new_n30779_ = ~new_n30574_ & ~new_n30769_;
  assign new_n30780_ = ~new_n30584_ & new_n30756_;
  assign new_n30781_ = ~new_n30752_ & new_n30780_;
  assign new_n30782_ = ~new_n30753_ & ~new_n30756_;
  assign new_n30783_ = ~new_n30781_ & ~new_n30782_;
  assign new_n30784_ = new_n475_ & ~new_n30783_;
  assign new_n30785_ = ~new_n30768_ & new_n30784_;
  assign new_n30786_ = ~new_n30779_ & ~new_n30785_;
  assign new_n30787_ = ~\b[15]  & ~new_n30786_;
  assign new_n30788_ = ~new_n30583_ & ~new_n30769_;
  assign new_n30789_ = ~new_n30593_ & new_n30751_;
  assign new_n30790_ = ~new_n30747_ & new_n30789_;
  assign new_n30791_ = ~new_n30748_ & ~new_n30751_;
  assign new_n30792_ = ~new_n30790_ & ~new_n30791_;
  assign new_n30793_ = new_n475_ & ~new_n30792_;
  assign new_n30794_ = ~new_n30768_ & new_n30793_;
  assign new_n30795_ = ~new_n30788_ & ~new_n30794_;
  assign new_n30796_ = ~\b[14]  & ~new_n30795_;
  assign new_n30797_ = ~new_n30592_ & ~new_n30769_;
  assign new_n30798_ = ~new_n30602_ & new_n30746_;
  assign new_n30799_ = ~new_n30742_ & new_n30798_;
  assign new_n30800_ = ~new_n30743_ & ~new_n30746_;
  assign new_n30801_ = ~new_n30799_ & ~new_n30800_;
  assign new_n30802_ = new_n475_ & ~new_n30801_;
  assign new_n30803_ = ~new_n30768_ & new_n30802_;
  assign new_n30804_ = ~new_n30797_ & ~new_n30803_;
  assign new_n30805_ = ~\b[13]  & ~new_n30804_;
  assign new_n30806_ = ~new_n30601_ & ~new_n30769_;
  assign new_n30807_ = ~new_n30611_ & new_n30741_;
  assign new_n30808_ = ~new_n30737_ & new_n30807_;
  assign new_n30809_ = ~new_n30738_ & ~new_n30741_;
  assign new_n30810_ = ~new_n30808_ & ~new_n30809_;
  assign new_n30811_ = new_n475_ & ~new_n30810_;
  assign new_n30812_ = ~new_n30768_ & new_n30811_;
  assign new_n30813_ = ~new_n30806_ & ~new_n30812_;
  assign new_n30814_ = ~\b[12]  & ~new_n30813_;
  assign new_n30815_ = ~new_n30610_ & ~new_n30769_;
  assign new_n30816_ = ~new_n30620_ & new_n30736_;
  assign new_n30817_ = ~new_n30732_ & new_n30816_;
  assign new_n30818_ = ~new_n30733_ & ~new_n30736_;
  assign new_n30819_ = ~new_n30817_ & ~new_n30818_;
  assign new_n30820_ = new_n475_ & ~new_n30819_;
  assign new_n30821_ = ~new_n30768_ & new_n30820_;
  assign new_n30822_ = ~new_n30815_ & ~new_n30821_;
  assign new_n30823_ = ~\b[11]  & ~new_n30822_;
  assign new_n30824_ = ~new_n30619_ & ~new_n30769_;
  assign new_n30825_ = ~new_n30629_ & new_n30731_;
  assign new_n30826_ = ~new_n30727_ & new_n30825_;
  assign new_n30827_ = ~new_n30728_ & ~new_n30731_;
  assign new_n30828_ = ~new_n30826_ & ~new_n30827_;
  assign new_n30829_ = new_n475_ & ~new_n30828_;
  assign new_n30830_ = ~new_n30768_ & new_n30829_;
  assign new_n30831_ = ~new_n30824_ & ~new_n30830_;
  assign new_n30832_ = ~\b[10]  & ~new_n30831_;
  assign new_n30833_ = ~new_n30628_ & ~new_n30769_;
  assign new_n30834_ = ~new_n30638_ & new_n30726_;
  assign new_n30835_ = ~new_n30722_ & new_n30834_;
  assign new_n30836_ = ~new_n30723_ & ~new_n30726_;
  assign new_n30837_ = ~new_n30835_ & ~new_n30836_;
  assign new_n30838_ = new_n475_ & ~new_n30837_;
  assign new_n30839_ = ~new_n30768_ & new_n30838_;
  assign new_n30840_ = ~new_n30833_ & ~new_n30839_;
  assign new_n30841_ = ~\b[9]  & ~new_n30840_;
  assign new_n30842_ = ~new_n30637_ & ~new_n30769_;
  assign new_n30843_ = ~new_n30647_ & new_n30721_;
  assign new_n30844_ = ~new_n30717_ & new_n30843_;
  assign new_n30845_ = ~new_n30718_ & ~new_n30721_;
  assign new_n30846_ = ~new_n30844_ & ~new_n30845_;
  assign new_n30847_ = new_n475_ & ~new_n30846_;
  assign new_n30848_ = ~new_n30768_ & new_n30847_;
  assign new_n30849_ = ~new_n30842_ & ~new_n30848_;
  assign new_n30850_ = ~\b[8]  & ~new_n30849_;
  assign new_n30851_ = ~new_n30646_ & ~new_n30769_;
  assign new_n30852_ = ~new_n30656_ & new_n30716_;
  assign new_n30853_ = ~new_n30712_ & new_n30852_;
  assign new_n30854_ = ~new_n30713_ & ~new_n30716_;
  assign new_n30855_ = ~new_n30853_ & ~new_n30854_;
  assign new_n30856_ = new_n475_ & ~new_n30855_;
  assign new_n30857_ = ~new_n30768_ & new_n30856_;
  assign new_n30858_ = ~new_n30851_ & ~new_n30857_;
  assign new_n30859_ = ~\b[7]  & ~new_n30858_;
  assign new_n30860_ = ~new_n30655_ & ~new_n30769_;
  assign new_n30861_ = ~new_n30665_ & new_n30711_;
  assign new_n30862_ = ~new_n30707_ & new_n30861_;
  assign new_n30863_ = ~new_n30708_ & ~new_n30711_;
  assign new_n30864_ = ~new_n30862_ & ~new_n30863_;
  assign new_n30865_ = new_n475_ & ~new_n30864_;
  assign new_n30866_ = ~new_n30768_ & new_n30865_;
  assign new_n30867_ = ~new_n30860_ & ~new_n30866_;
  assign new_n30868_ = ~\b[6]  & ~new_n30867_;
  assign new_n30869_ = ~new_n30664_ & ~new_n30769_;
  assign new_n30870_ = ~new_n30674_ & new_n30706_;
  assign new_n30871_ = ~new_n30702_ & new_n30870_;
  assign new_n30872_ = ~new_n30703_ & ~new_n30706_;
  assign new_n30873_ = ~new_n30871_ & ~new_n30872_;
  assign new_n30874_ = new_n475_ & ~new_n30873_;
  assign new_n30875_ = ~new_n30768_ & new_n30874_;
  assign new_n30876_ = ~new_n30869_ & ~new_n30875_;
  assign new_n30877_ = ~\b[5]  & ~new_n30876_;
  assign new_n30878_ = ~new_n30673_ & ~new_n30769_;
  assign new_n30879_ = ~new_n30682_ & new_n30701_;
  assign new_n30880_ = ~new_n30697_ & new_n30879_;
  assign new_n30881_ = ~new_n30698_ & ~new_n30701_;
  assign new_n30882_ = ~new_n30880_ & ~new_n30881_;
  assign new_n30883_ = new_n475_ & ~new_n30882_;
  assign new_n30884_ = ~new_n30768_ & new_n30883_;
  assign new_n30885_ = ~new_n30878_ & ~new_n30884_;
  assign new_n30886_ = ~\b[4]  & ~new_n30885_;
  assign new_n30887_ = ~new_n30681_ & ~new_n30769_;
  assign new_n30888_ = ~new_n30692_ & new_n30696_;
  assign new_n30889_ = ~new_n30691_ & new_n30888_;
  assign new_n30890_ = ~new_n30693_ & ~new_n30696_;
  assign new_n30891_ = ~new_n30889_ & ~new_n30890_;
  assign new_n30892_ = new_n475_ & ~new_n30891_;
  assign new_n30893_ = ~new_n30768_ & new_n30892_;
  assign new_n30894_ = ~new_n30887_ & ~new_n30893_;
  assign new_n30895_ = ~\b[3]  & ~new_n30894_;
  assign new_n30896_ = ~new_n30686_ & ~new_n30769_;
  assign new_n30897_ = new_n2382_ & ~new_n30689_;
  assign new_n30898_ = ~new_n30687_ & new_n30897_;
  assign new_n30899_ = new_n475_ & ~new_n30898_;
  assign new_n30900_ = ~new_n30691_ & new_n30899_;
  assign new_n30901_ = ~new_n30768_ & new_n30900_;
  assign new_n30902_ = ~new_n30896_ & ~new_n30901_;
  assign new_n30903_ = ~\b[2]  & ~new_n30902_;
  assign new_n30904_ = new_n2601_ & ~new_n30768_;
  assign new_n30905_ = \a[47]  & ~new_n30904_;
  assign new_n30906_ = new_n2606_ & ~new_n30768_;
  assign new_n30907_ = ~new_n30905_ & ~new_n30906_;
  assign new_n30908_ = \b[1]  & ~new_n30907_;
  assign new_n30909_ = ~\b[1]  & ~new_n30906_;
  assign new_n30910_ = ~new_n30905_ & new_n30909_;
  assign new_n30911_ = ~new_n30908_ & ~new_n30910_;
  assign new_n30912_ = ~new_n2613_ & ~new_n30911_;
  assign new_n30913_ = ~\b[1]  & ~new_n30907_;
  assign new_n30914_ = ~new_n30912_ & ~new_n30913_;
  assign new_n30915_ = \b[2]  & ~new_n30901_;
  assign new_n30916_ = ~new_n30896_ & new_n30915_;
  assign new_n30917_ = ~new_n30903_ & ~new_n30916_;
  assign new_n30918_ = ~new_n30914_ & new_n30917_;
  assign new_n30919_ = ~new_n30903_ & ~new_n30918_;
  assign new_n30920_ = \b[3]  & ~new_n30893_;
  assign new_n30921_ = ~new_n30887_ & new_n30920_;
  assign new_n30922_ = ~new_n30895_ & ~new_n30921_;
  assign new_n30923_ = ~new_n30919_ & new_n30922_;
  assign new_n30924_ = ~new_n30895_ & ~new_n30923_;
  assign new_n30925_ = \b[4]  & ~new_n30884_;
  assign new_n30926_ = ~new_n30878_ & new_n30925_;
  assign new_n30927_ = ~new_n30886_ & ~new_n30926_;
  assign new_n30928_ = ~new_n30924_ & new_n30927_;
  assign new_n30929_ = ~new_n30886_ & ~new_n30928_;
  assign new_n30930_ = \b[5]  & ~new_n30875_;
  assign new_n30931_ = ~new_n30869_ & new_n30930_;
  assign new_n30932_ = ~new_n30877_ & ~new_n30931_;
  assign new_n30933_ = ~new_n30929_ & new_n30932_;
  assign new_n30934_ = ~new_n30877_ & ~new_n30933_;
  assign new_n30935_ = \b[6]  & ~new_n30866_;
  assign new_n30936_ = ~new_n30860_ & new_n30935_;
  assign new_n30937_ = ~new_n30868_ & ~new_n30936_;
  assign new_n30938_ = ~new_n30934_ & new_n30937_;
  assign new_n30939_ = ~new_n30868_ & ~new_n30938_;
  assign new_n30940_ = \b[7]  & ~new_n30857_;
  assign new_n30941_ = ~new_n30851_ & new_n30940_;
  assign new_n30942_ = ~new_n30859_ & ~new_n30941_;
  assign new_n30943_ = ~new_n30939_ & new_n30942_;
  assign new_n30944_ = ~new_n30859_ & ~new_n30943_;
  assign new_n30945_ = \b[8]  & ~new_n30848_;
  assign new_n30946_ = ~new_n30842_ & new_n30945_;
  assign new_n30947_ = ~new_n30850_ & ~new_n30946_;
  assign new_n30948_ = ~new_n30944_ & new_n30947_;
  assign new_n30949_ = ~new_n30850_ & ~new_n30948_;
  assign new_n30950_ = \b[9]  & ~new_n30839_;
  assign new_n30951_ = ~new_n30833_ & new_n30950_;
  assign new_n30952_ = ~new_n30841_ & ~new_n30951_;
  assign new_n30953_ = ~new_n30949_ & new_n30952_;
  assign new_n30954_ = ~new_n30841_ & ~new_n30953_;
  assign new_n30955_ = \b[10]  & ~new_n30830_;
  assign new_n30956_ = ~new_n30824_ & new_n30955_;
  assign new_n30957_ = ~new_n30832_ & ~new_n30956_;
  assign new_n30958_ = ~new_n30954_ & new_n30957_;
  assign new_n30959_ = ~new_n30832_ & ~new_n30958_;
  assign new_n30960_ = \b[11]  & ~new_n30821_;
  assign new_n30961_ = ~new_n30815_ & new_n30960_;
  assign new_n30962_ = ~new_n30823_ & ~new_n30961_;
  assign new_n30963_ = ~new_n30959_ & new_n30962_;
  assign new_n30964_ = ~new_n30823_ & ~new_n30963_;
  assign new_n30965_ = \b[12]  & ~new_n30812_;
  assign new_n30966_ = ~new_n30806_ & new_n30965_;
  assign new_n30967_ = ~new_n30814_ & ~new_n30966_;
  assign new_n30968_ = ~new_n30964_ & new_n30967_;
  assign new_n30969_ = ~new_n30814_ & ~new_n30968_;
  assign new_n30970_ = \b[13]  & ~new_n30803_;
  assign new_n30971_ = ~new_n30797_ & new_n30970_;
  assign new_n30972_ = ~new_n30805_ & ~new_n30971_;
  assign new_n30973_ = ~new_n30969_ & new_n30972_;
  assign new_n30974_ = ~new_n30805_ & ~new_n30973_;
  assign new_n30975_ = \b[14]  & ~new_n30794_;
  assign new_n30976_ = ~new_n30788_ & new_n30975_;
  assign new_n30977_ = ~new_n30796_ & ~new_n30976_;
  assign new_n30978_ = ~new_n30974_ & new_n30977_;
  assign new_n30979_ = ~new_n30796_ & ~new_n30978_;
  assign new_n30980_ = \b[15]  & ~new_n30785_;
  assign new_n30981_ = ~new_n30779_ & new_n30980_;
  assign new_n30982_ = ~new_n30787_ & ~new_n30981_;
  assign new_n30983_ = ~new_n30979_ & new_n30982_;
  assign new_n30984_ = ~new_n30787_ & ~new_n30983_;
  assign new_n30985_ = \b[16]  & ~new_n30776_;
  assign new_n30986_ = ~new_n30770_ & new_n30985_;
  assign new_n30987_ = ~new_n30778_ & ~new_n30986_;
  assign new_n30988_ = ~new_n30984_ & new_n30987_;
  assign new_n30989_ = ~new_n30778_ & ~new_n30988_;
  assign new_n30990_ = ~new_n30564_ & ~new_n30769_;
  assign new_n30991_ = ~new_n30566_ & new_n30766_;
  assign new_n30992_ = ~new_n30762_ & new_n30991_;
  assign new_n30993_ = ~new_n30763_ & ~new_n30766_;
  assign new_n30994_ = ~new_n30992_ & ~new_n30993_;
  assign new_n30995_ = new_n30769_ & ~new_n30994_;
  assign new_n30996_ = ~new_n30990_ & ~new_n30995_;
  assign new_n30997_ = ~\b[17]  & ~new_n30996_;
  assign new_n30998_ = \b[17]  & ~new_n30990_;
  assign new_n30999_ = ~new_n30995_ & new_n30998_;
  assign new_n31000_ = new_n2705_ & ~new_n30999_;
  assign new_n31001_ = ~new_n30997_ & new_n31000_;
  assign new_n31002_ = ~new_n30989_ & new_n31001_;
  assign new_n31003_ = new_n475_ & ~new_n30996_;
  assign new_n31004_ = ~new_n31002_ & ~new_n31003_;
  assign new_n31005_ = ~new_n30787_ & new_n30987_;
  assign new_n31006_ = ~new_n30983_ & new_n31005_;
  assign new_n31007_ = ~new_n30984_ & ~new_n30987_;
  assign new_n31008_ = ~new_n31006_ & ~new_n31007_;
  assign new_n31009_ = ~new_n31004_ & ~new_n31008_;
  assign new_n31010_ = ~new_n30777_ & ~new_n31003_;
  assign new_n31011_ = ~new_n31002_ & new_n31010_;
  assign new_n31012_ = ~new_n31009_ & ~new_n31011_;
  assign new_n31013_ = ~new_n30778_ & ~new_n30999_;
  assign new_n31014_ = ~new_n30997_ & new_n31013_;
  assign new_n31015_ = ~new_n30988_ & new_n31014_;
  assign new_n31016_ = ~new_n30997_ & ~new_n30999_;
  assign new_n31017_ = ~new_n30989_ & ~new_n31016_;
  assign new_n31018_ = ~new_n31015_ & ~new_n31017_;
  assign new_n31019_ = ~new_n31004_ & ~new_n31018_;
  assign new_n31020_ = ~new_n30996_ & ~new_n31003_;
  assign new_n31021_ = ~new_n31002_ & new_n31020_;
  assign new_n31022_ = ~new_n31019_ & ~new_n31021_;
  assign new_n31023_ = ~\b[18]  & ~new_n31022_;
  assign new_n31024_ = ~\b[17]  & ~new_n31012_;
  assign new_n31025_ = ~new_n30796_ & new_n30982_;
  assign new_n31026_ = ~new_n30978_ & new_n31025_;
  assign new_n31027_ = ~new_n30979_ & ~new_n30982_;
  assign new_n31028_ = ~new_n31026_ & ~new_n31027_;
  assign new_n31029_ = ~new_n31004_ & ~new_n31028_;
  assign new_n31030_ = ~new_n30786_ & ~new_n31003_;
  assign new_n31031_ = ~new_n31002_ & new_n31030_;
  assign new_n31032_ = ~new_n31029_ & ~new_n31031_;
  assign new_n31033_ = ~\b[16]  & ~new_n31032_;
  assign new_n31034_ = ~new_n30805_ & new_n30977_;
  assign new_n31035_ = ~new_n30973_ & new_n31034_;
  assign new_n31036_ = ~new_n30974_ & ~new_n30977_;
  assign new_n31037_ = ~new_n31035_ & ~new_n31036_;
  assign new_n31038_ = ~new_n31004_ & ~new_n31037_;
  assign new_n31039_ = ~new_n30795_ & ~new_n31003_;
  assign new_n31040_ = ~new_n31002_ & new_n31039_;
  assign new_n31041_ = ~new_n31038_ & ~new_n31040_;
  assign new_n31042_ = ~\b[15]  & ~new_n31041_;
  assign new_n31043_ = ~new_n30814_ & new_n30972_;
  assign new_n31044_ = ~new_n30968_ & new_n31043_;
  assign new_n31045_ = ~new_n30969_ & ~new_n30972_;
  assign new_n31046_ = ~new_n31044_ & ~new_n31045_;
  assign new_n31047_ = ~new_n31004_ & ~new_n31046_;
  assign new_n31048_ = ~new_n30804_ & ~new_n31003_;
  assign new_n31049_ = ~new_n31002_ & new_n31048_;
  assign new_n31050_ = ~new_n31047_ & ~new_n31049_;
  assign new_n31051_ = ~\b[14]  & ~new_n31050_;
  assign new_n31052_ = ~new_n30823_ & new_n30967_;
  assign new_n31053_ = ~new_n30963_ & new_n31052_;
  assign new_n31054_ = ~new_n30964_ & ~new_n30967_;
  assign new_n31055_ = ~new_n31053_ & ~new_n31054_;
  assign new_n31056_ = ~new_n31004_ & ~new_n31055_;
  assign new_n31057_ = ~new_n30813_ & ~new_n31003_;
  assign new_n31058_ = ~new_n31002_ & new_n31057_;
  assign new_n31059_ = ~new_n31056_ & ~new_n31058_;
  assign new_n31060_ = ~\b[13]  & ~new_n31059_;
  assign new_n31061_ = ~new_n30832_ & new_n30962_;
  assign new_n31062_ = ~new_n30958_ & new_n31061_;
  assign new_n31063_ = ~new_n30959_ & ~new_n30962_;
  assign new_n31064_ = ~new_n31062_ & ~new_n31063_;
  assign new_n31065_ = ~new_n31004_ & ~new_n31064_;
  assign new_n31066_ = ~new_n30822_ & ~new_n31003_;
  assign new_n31067_ = ~new_n31002_ & new_n31066_;
  assign new_n31068_ = ~new_n31065_ & ~new_n31067_;
  assign new_n31069_ = ~\b[12]  & ~new_n31068_;
  assign new_n31070_ = ~new_n30841_ & new_n30957_;
  assign new_n31071_ = ~new_n30953_ & new_n31070_;
  assign new_n31072_ = ~new_n30954_ & ~new_n30957_;
  assign new_n31073_ = ~new_n31071_ & ~new_n31072_;
  assign new_n31074_ = ~new_n31004_ & ~new_n31073_;
  assign new_n31075_ = ~new_n30831_ & ~new_n31003_;
  assign new_n31076_ = ~new_n31002_ & new_n31075_;
  assign new_n31077_ = ~new_n31074_ & ~new_n31076_;
  assign new_n31078_ = ~\b[11]  & ~new_n31077_;
  assign new_n31079_ = ~new_n30850_ & new_n30952_;
  assign new_n31080_ = ~new_n30948_ & new_n31079_;
  assign new_n31081_ = ~new_n30949_ & ~new_n30952_;
  assign new_n31082_ = ~new_n31080_ & ~new_n31081_;
  assign new_n31083_ = ~new_n31004_ & ~new_n31082_;
  assign new_n31084_ = ~new_n30840_ & ~new_n31003_;
  assign new_n31085_ = ~new_n31002_ & new_n31084_;
  assign new_n31086_ = ~new_n31083_ & ~new_n31085_;
  assign new_n31087_ = ~\b[10]  & ~new_n31086_;
  assign new_n31088_ = ~new_n30859_ & new_n30947_;
  assign new_n31089_ = ~new_n30943_ & new_n31088_;
  assign new_n31090_ = ~new_n30944_ & ~new_n30947_;
  assign new_n31091_ = ~new_n31089_ & ~new_n31090_;
  assign new_n31092_ = ~new_n31004_ & ~new_n31091_;
  assign new_n31093_ = ~new_n30849_ & ~new_n31003_;
  assign new_n31094_ = ~new_n31002_ & new_n31093_;
  assign new_n31095_ = ~new_n31092_ & ~new_n31094_;
  assign new_n31096_ = ~\b[9]  & ~new_n31095_;
  assign new_n31097_ = ~new_n30868_ & new_n30942_;
  assign new_n31098_ = ~new_n30938_ & new_n31097_;
  assign new_n31099_ = ~new_n30939_ & ~new_n30942_;
  assign new_n31100_ = ~new_n31098_ & ~new_n31099_;
  assign new_n31101_ = ~new_n31004_ & ~new_n31100_;
  assign new_n31102_ = ~new_n30858_ & ~new_n31003_;
  assign new_n31103_ = ~new_n31002_ & new_n31102_;
  assign new_n31104_ = ~new_n31101_ & ~new_n31103_;
  assign new_n31105_ = ~\b[8]  & ~new_n31104_;
  assign new_n31106_ = ~new_n30877_ & new_n30937_;
  assign new_n31107_ = ~new_n30933_ & new_n31106_;
  assign new_n31108_ = ~new_n30934_ & ~new_n30937_;
  assign new_n31109_ = ~new_n31107_ & ~new_n31108_;
  assign new_n31110_ = ~new_n31004_ & ~new_n31109_;
  assign new_n31111_ = ~new_n30867_ & ~new_n31003_;
  assign new_n31112_ = ~new_n31002_ & new_n31111_;
  assign new_n31113_ = ~new_n31110_ & ~new_n31112_;
  assign new_n31114_ = ~\b[7]  & ~new_n31113_;
  assign new_n31115_ = ~new_n30886_ & new_n30932_;
  assign new_n31116_ = ~new_n30928_ & new_n31115_;
  assign new_n31117_ = ~new_n30929_ & ~new_n30932_;
  assign new_n31118_ = ~new_n31116_ & ~new_n31117_;
  assign new_n31119_ = ~new_n31004_ & ~new_n31118_;
  assign new_n31120_ = ~new_n30876_ & ~new_n31003_;
  assign new_n31121_ = ~new_n31002_ & new_n31120_;
  assign new_n31122_ = ~new_n31119_ & ~new_n31121_;
  assign new_n31123_ = ~\b[6]  & ~new_n31122_;
  assign new_n31124_ = ~new_n30895_ & new_n30927_;
  assign new_n31125_ = ~new_n30923_ & new_n31124_;
  assign new_n31126_ = ~new_n30924_ & ~new_n30927_;
  assign new_n31127_ = ~new_n31125_ & ~new_n31126_;
  assign new_n31128_ = ~new_n31004_ & ~new_n31127_;
  assign new_n31129_ = ~new_n30885_ & ~new_n31003_;
  assign new_n31130_ = ~new_n31002_ & new_n31129_;
  assign new_n31131_ = ~new_n31128_ & ~new_n31130_;
  assign new_n31132_ = ~\b[5]  & ~new_n31131_;
  assign new_n31133_ = ~new_n30903_ & new_n30922_;
  assign new_n31134_ = ~new_n30918_ & new_n31133_;
  assign new_n31135_ = ~new_n30919_ & ~new_n30922_;
  assign new_n31136_ = ~new_n31134_ & ~new_n31135_;
  assign new_n31137_ = ~new_n31004_ & ~new_n31136_;
  assign new_n31138_ = ~new_n30894_ & ~new_n31003_;
  assign new_n31139_ = ~new_n31002_ & new_n31138_;
  assign new_n31140_ = ~new_n31137_ & ~new_n31139_;
  assign new_n31141_ = ~\b[4]  & ~new_n31140_;
  assign new_n31142_ = ~new_n30913_ & new_n30917_;
  assign new_n31143_ = ~new_n30912_ & new_n31142_;
  assign new_n31144_ = ~new_n30914_ & ~new_n30917_;
  assign new_n31145_ = ~new_n31143_ & ~new_n31144_;
  assign new_n31146_ = ~new_n31004_ & ~new_n31145_;
  assign new_n31147_ = ~new_n30902_ & ~new_n31003_;
  assign new_n31148_ = ~new_n31002_ & new_n31147_;
  assign new_n31149_ = ~new_n31146_ & ~new_n31148_;
  assign new_n31150_ = ~\b[3]  & ~new_n31149_;
  assign new_n31151_ = new_n2613_ & ~new_n30910_;
  assign new_n31152_ = ~new_n30908_ & new_n31151_;
  assign new_n31153_ = ~new_n30912_ & ~new_n31152_;
  assign new_n31154_ = ~new_n31004_ & new_n31153_;
  assign new_n31155_ = ~new_n30907_ & ~new_n31003_;
  assign new_n31156_ = ~new_n31002_ & new_n31155_;
  assign new_n31157_ = ~new_n31154_ & ~new_n31156_;
  assign new_n31158_ = ~\b[2]  & ~new_n31157_;
  assign new_n31159_ = \b[0]  & ~new_n31004_;
  assign new_n31160_ = \a[46]  & ~new_n31159_;
  assign new_n31161_ = new_n2613_ & ~new_n31004_;
  assign new_n31162_ = ~new_n31160_ & ~new_n31161_;
  assign new_n31163_ = \b[1]  & ~new_n31162_;
  assign new_n31164_ = ~\b[1]  & ~new_n31161_;
  assign new_n31165_ = ~new_n31160_ & new_n31164_;
  assign new_n31166_ = ~new_n31163_ & ~new_n31165_;
  assign new_n31167_ = ~new_n2873_ & ~new_n31166_;
  assign new_n31168_ = ~\b[1]  & ~new_n31162_;
  assign new_n31169_ = ~new_n31167_ & ~new_n31168_;
  assign new_n31170_ = \b[2]  & ~new_n31156_;
  assign new_n31171_ = ~new_n31154_ & new_n31170_;
  assign new_n31172_ = ~new_n31158_ & ~new_n31171_;
  assign new_n31173_ = ~new_n31169_ & new_n31172_;
  assign new_n31174_ = ~new_n31158_ & ~new_n31173_;
  assign new_n31175_ = \b[3]  & ~new_n31148_;
  assign new_n31176_ = ~new_n31146_ & new_n31175_;
  assign new_n31177_ = ~new_n31150_ & ~new_n31176_;
  assign new_n31178_ = ~new_n31174_ & new_n31177_;
  assign new_n31179_ = ~new_n31150_ & ~new_n31178_;
  assign new_n31180_ = \b[4]  & ~new_n31139_;
  assign new_n31181_ = ~new_n31137_ & new_n31180_;
  assign new_n31182_ = ~new_n31141_ & ~new_n31181_;
  assign new_n31183_ = ~new_n31179_ & new_n31182_;
  assign new_n31184_ = ~new_n31141_ & ~new_n31183_;
  assign new_n31185_ = \b[5]  & ~new_n31130_;
  assign new_n31186_ = ~new_n31128_ & new_n31185_;
  assign new_n31187_ = ~new_n31132_ & ~new_n31186_;
  assign new_n31188_ = ~new_n31184_ & new_n31187_;
  assign new_n31189_ = ~new_n31132_ & ~new_n31188_;
  assign new_n31190_ = \b[6]  & ~new_n31121_;
  assign new_n31191_ = ~new_n31119_ & new_n31190_;
  assign new_n31192_ = ~new_n31123_ & ~new_n31191_;
  assign new_n31193_ = ~new_n31189_ & new_n31192_;
  assign new_n31194_ = ~new_n31123_ & ~new_n31193_;
  assign new_n31195_ = \b[7]  & ~new_n31112_;
  assign new_n31196_ = ~new_n31110_ & new_n31195_;
  assign new_n31197_ = ~new_n31114_ & ~new_n31196_;
  assign new_n31198_ = ~new_n31194_ & new_n31197_;
  assign new_n31199_ = ~new_n31114_ & ~new_n31198_;
  assign new_n31200_ = \b[8]  & ~new_n31103_;
  assign new_n31201_ = ~new_n31101_ & new_n31200_;
  assign new_n31202_ = ~new_n31105_ & ~new_n31201_;
  assign new_n31203_ = ~new_n31199_ & new_n31202_;
  assign new_n31204_ = ~new_n31105_ & ~new_n31203_;
  assign new_n31205_ = \b[9]  & ~new_n31094_;
  assign new_n31206_ = ~new_n31092_ & new_n31205_;
  assign new_n31207_ = ~new_n31096_ & ~new_n31206_;
  assign new_n31208_ = ~new_n31204_ & new_n31207_;
  assign new_n31209_ = ~new_n31096_ & ~new_n31208_;
  assign new_n31210_ = \b[10]  & ~new_n31085_;
  assign new_n31211_ = ~new_n31083_ & new_n31210_;
  assign new_n31212_ = ~new_n31087_ & ~new_n31211_;
  assign new_n31213_ = ~new_n31209_ & new_n31212_;
  assign new_n31214_ = ~new_n31087_ & ~new_n31213_;
  assign new_n31215_ = \b[11]  & ~new_n31076_;
  assign new_n31216_ = ~new_n31074_ & new_n31215_;
  assign new_n31217_ = ~new_n31078_ & ~new_n31216_;
  assign new_n31218_ = ~new_n31214_ & new_n31217_;
  assign new_n31219_ = ~new_n31078_ & ~new_n31218_;
  assign new_n31220_ = \b[12]  & ~new_n31067_;
  assign new_n31221_ = ~new_n31065_ & new_n31220_;
  assign new_n31222_ = ~new_n31069_ & ~new_n31221_;
  assign new_n31223_ = ~new_n31219_ & new_n31222_;
  assign new_n31224_ = ~new_n31069_ & ~new_n31223_;
  assign new_n31225_ = \b[13]  & ~new_n31058_;
  assign new_n31226_ = ~new_n31056_ & new_n31225_;
  assign new_n31227_ = ~new_n31060_ & ~new_n31226_;
  assign new_n31228_ = ~new_n31224_ & new_n31227_;
  assign new_n31229_ = ~new_n31060_ & ~new_n31228_;
  assign new_n31230_ = \b[14]  & ~new_n31049_;
  assign new_n31231_ = ~new_n31047_ & new_n31230_;
  assign new_n31232_ = ~new_n31051_ & ~new_n31231_;
  assign new_n31233_ = ~new_n31229_ & new_n31232_;
  assign new_n31234_ = ~new_n31051_ & ~new_n31233_;
  assign new_n31235_ = \b[15]  & ~new_n31040_;
  assign new_n31236_ = ~new_n31038_ & new_n31235_;
  assign new_n31237_ = ~new_n31042_ & ~new_n31236_;
  assign new_n31238_ = ~new_n31234_ & new_n31237_;
  assign new_n31239_ = ~new_n31042_ & ~new_n31238_;
  assign new_n31240_ = \b[16]  & ~new_n31031_;
  assign new_n31241_ = ~new_n31029_ & new_n31240_;
  assign new_n31242_ = ~new_n31033_ & ~new_n31241_;
  assign new_n31243_ = ~new_n31239_ & new_n31242_;
  assign new_n31244_ = ~new_n31033_ & ~new_n31243_;
  assign new_n31245_ = \b[17]  & ~new_n31011_;
  assign new_n31246_ = ~new_n31009_ & new_n31245_;
  assign new_n31247_ = ~new_n31024_ & ~new_n31246_;
  assign new_n31248_ = ~new_n31244_ & new_n31247_;
  assign new_n31249_ = ~new_n31024_ & ~new_n31248_;
  assign new_n31250_ = \b[18]  & ~new_n31021_;
  assign new_n31251_ = ~new_n31019_ & new_n31250_;
  assign new_n31252_ = ~new_n31023_ & ~new_n31251_;
  assign new_n31253_ = ~new_n31249_ & new_n31252_;
  assign new_n31254_ = ~new_n31023_ & ~new_n31253_;
  assign new_n31255_ = new_n2965_ & ~new_n31254_;
  assign new_n31256_ = ~new_n31012_ & ~new_n31255_;
  assign new_n31257_ = ~new_n31033_ & new_n31247_;
  assign new_n31258_ = ~new_n31243_ & new_n31257_;
  assign new_n31259_ = ~new_n31244_ & ~new_n31247_;
  assign new_n31260_ = ~new_n31258_ & ~new_n31259_;
  assign new_n31261_ = new_n2965_ & ~new_n31260_;
  assign new_n31262_ = ~new_n31254_ & new_n31261_;
  assign new_n31263_ = ~new_n31256_ & ~new_n31262_;
  assign new_n31264_ = ~new_n31022_ & ~new_n31255_;
  assign new_n31265_ = ~new_n31024_ & new_n31252_;
  assign new_n31266_ = ~new_n31248_ & new_n31265_;
  assign new_n31267_ = ~new_n31249_ & ~new_n31252_;
  assign new_n31268_ = ~new_n31266_ & ~new_n31267_;
  assign new_n31269_ = new_n31255_ & ~new_n31268_;
  assign new_n31270_ = ~new_n31264_ & ~new_n31269_;
  assign new_n31271_ = ~\b[19]  & ~new_n31270_;
  assign new_n31272_ = ~\b[18]  & ~new_n31263_;
  assign new_n31273_ = ~new_n31032_ & ~new_n31255_;
  assign new_n31274_ = ~new_n31042_ & new_n31242_;
  assign new_n31275_ = ~new_n31238_ & new_n31274_;
  assign new_n31276_ = ~new_n31239_ & ~new_n31242_;
  assign new_n31277_ = ~new_n31275_ & ~new_n31276_;
  assign new_n31278_ = new_n2965_ & ~new_n31277_;
  assign new_n31279_ = ~new_n31254_ & new_n31278_;
  assign new_n31280_ = ~new_n31273_ & ~new_n31279_;
  assign new_n31281_ = ~\b[17]  & ~new_n31280_;
  assign new_n31282_ = ~new_n31041_ & ~new_n31255_;
  assign new_n31283_ = ~new_n31051_ & new_n31237_;
  assign new_n31284_ = ~new_n31233_ & new_n31283_;
  assign new_n31285_ = ~new_n31234_ & ~new_n31237_;
  assign new_n31286_ = ~new_n31284_ & ~new_n31285_;
  assign new_n31287_ = new_n2965_ & ~new_n31286_;
  assign new_n31288_ = ~new_n31254_ & new_n31287_;
  assign new_n31289_ = ~new_n31282_ & ~new_n31288_;
  assign new_n31290_ = ~\b[16]  & ~new_n31289_;
  assign new_n31291_ = ~new_n31050_ & ~new_n31255_;
  assign new_n31292_ = ~new_n31060_ & new_n31232_;
  assign new_n31293_ = ~new_n31228_ & new_n31292_;
  assign new_n31294_ = ~new_n31229_ & ~new_n31232_;
  assign new_n31295_ = ~new_n31293_ & ~new_n31294_;
  assign new_n31296_ = new_n2965_ & ~new_n31295_;
  assign new_n31297_ = ~new_n31254_ & new_n31296_;
  assign new_n31298_ = ~new_n31291_ & ~new_n31297_;
  assign new_n31299_ = ~\b[15]  & ~new_n31298_;
  assign new_n31300_ = ~new_n31059_ & ~new_n31255_;
  assign new_n31301_ = ~new_n31069_ & new_n31227_;
  assign new_n31302_ = ~new_n31223_ & new_n31301_;
  assign new_n31303_ = ~new_n31224_ & ~new_n31227_;
  assign new_n31304_ = ~new_n31302_ & ~new_n31303_;
  assign new_n31305_ = new_n2965_ & ~new_n31304_;
  assign new_n31306_ = ~new_n31254_ & new_n31305_;
  assign new_n31307_ = ~new_n31300_ & ~new_n31306_;
  assign new_n31308_ = ~\b[14]  & ~new_n31307_;
  assign new_n31309_ = ~new_n31068_ & ~new_n31255_;
  assign new_n31310_ = ~new_n31078_ & new_n31222_;
  assign new_n31311_ = ~new_n31218_ & new_n31310_;
  assign new_n31312_ = ~new_n31219_ & ~new_n31222_;
  assign new_n31313_ = ~new_n31311_ & ~new_n31312_;
  assign new_n31314_ = new_n2965_ & ~new_n31313_;
  assign new_n31315_ = ~new_n31254_ & new_n31314_;
  assign new_n31316_ = ~new_n31309_ & ~new_n31315_;
  assign new_n31317_ = ~\b[13]  & ~new_n31316_;
  assign new_n31318_ = ~new_n31077_ & ~new_n31255_;
  assign new_n31319_ = ~new_n31087_ & new_n31217_;
  assign new_n31320_ = ~new_n31213_ & new_n31319_;
  assign new_n31321_ = ~new_n31214_ & ~new_n31217_;
  assign new_n31322_ = ~new_n31320_ & ~new_n31321_;
  assign new_n31323_ = new_n2965_ & ~new_n31322_;
  assign new_n31324_ = ~new_n31254_ & new_n31323_;
  assign new_n31325_ = ~new_n31318_ & ~new_n31324_;
  assign new_n31326_ = ~\b[12]  & ~new_n31325_;
  assign new_n31327_ = ~new_n31086_ & ~new_n31255_;
  assign new_n31328_ = ~new_n31096_ & new_n31212_;
  assign new_n31329_ = ~new_n31208_ & new_n31328_;
  assign new_n31330_ = ~new_n31209_ & ~new_n31212_;
  assign new_n31331_ = ~new_n31329_ & ~new_n31330_;
  assign new_n31332_ = new_n2965_ & ~new_n31331_;
  assign new_n31333_ = ~new_n31254_ & new_n31332_;
  assign new_n31334_ = ~new_n31327_ & ~new_n31333_;
  assign new_n31335_ = ~\b[11]  & ~new_n31334_;
  assign new_n31336_ = ~new_n31095_ & ~new_n31255_;
  assign new_n31337_ = ~new_n31105_ & new_n31207_;
  assign new_n31338_ = ~new_n31203_ & new_n31337_;
  assign new_n31339_ = ~new_n31204_ & ~new_n31207_;
  assign new_n31340_ = ~new_n31338_ & ~new_n31339_;
  assign new_n31341_ = new_n2965_ & ~new_n31340_;
  assign new_n31342_ = ~new_n31254_ & new_n31341_;
  assign new_n31343_ = ~new_n31336_ & ~new_n31342_;
  assign new_n31344_ = ~\b[10]  & ~new_n31343_;
  assign new_n31345_ = ~new_n31104_ & ~new_n31255_;
  assign new_n31346_ = ~new_n31114_ & new_n31202_;
  assign new_n31347_ = ~new_n31198_ & new_n31346_;
  assign new_n31348_ = ~new_n31199_ & ~new_n31202_;
  assign new_n31349_ = ~new_n31347_ & ~new_n31348_;
  assign new_n31350_ = new_n2965_ & ~new_n31349_;
  assign new_n31351_ = ~new_n31254_ & new_n31350_;
  assign new_n31352_ = ~new_n31345_ & ~new_n31351_;
  assign new_n31353_ = ~\b[9]  & ~new_n31352_;
  assign new_n31354_ = ~new_n31113_ & ~new_n31255_;
  assign new_n31355_ = ~new_n31123_ & new_n31197_;
  assign new_n31356_ = ~new_n31193_ & new_n31355_;
  assign new_n31357_ = ~new_n31194_ & ~new_n31197_;
  assign new_n31358_ = ~new_n31356_ & ~new_n31357_;
  assign new_n31359_ = new_n2965_ & ~new_n31358_;
  assign new_n31360_ = ~new_n31254_ & new_n31359_;
  assign new_n31361_ = ~new_n31354_ & ~new_n31360_;
  assign new_n31362_ = ~\b[8]  & ~new_n31361_;
  assign new_n31363_ = ~new_n31122_ & ~new_n31255_;
  assign new_n31364_ = ~new_n31132_ & new_n31192_;
  assign new_n31365_ = ~new_n31188_ & new_n31364_;
  assign new_n31366_ = ~new_n31189_ & ~new_n31192_;
  assign new_n31367_ = ~new_n31365_ & ~new_n31366_;
  assign new_n31368_ = new_n2965_ & ~new_n31367_;
  assign new_n31369_ = ~new_n31254_ & new_n31368_;
  assign new_n31370_ = ~new_n31363_ & ~new_n31369_;
  assign new_n31371_ = ~\b[7]  & ~new_n31370_;
  assign new_n31372_ = ~new_n31131_ & ~new_n31255_;
  assign new_n31373_ = ~new_n31141_ & new_n31187_;
  assign new_n31374_ = ~new_n31183_ & new_n31373_;
  assign new_n31375_ = ~new_n31184_ & ~new_n31187_;
  assign new_n31376_ = ~new_n31374_ & ~new_n31375_;
  assign new_n31377_ = new_n2965_ & ~new_n31376_;
  assign new_n31378_ = ~new_n31254_ & new_n31377_;
  assign new_n31379_ = ~new_n31372_ & ~new_n31378_;
  assign new_n31380_ = ~\b[6]  & ~new_n31379_;
  assign new_n31381_ = ~new_n31140_ & ~new_n31255_;
  assign new_n31382_ = ~new_n31150_ & new_n31182_;
  assign new_n31383_ = ~new_n31178_ & new_n31382_;
  assign new_n31384_ = ~new_n31179_ & ~new_n31182_;
  assign new_n31385_ = ~new_n31383_ & ~new_n31384_;
  assign new_n31386_ = new_n2965_ & ~new_n31385_;
  assign new_n31387_ = ~new_n31254_ & new_n31386_;
  assign new_n31388_ = ~new_n31381_ & ~new_n31387_;
  assign new_n31389_ = ~\b[5]  & ~new_n31388_;
  assign new_n31390_ = ~new_n31149_ & ~new_n31255_;
  assign new_n31391_ = ~new_n31158_ & new_n31177_;
  assign new_n31392_ = ~new_n31173_ & new_n31391_;
  assign new_n31393_ = ~new_n31174_ & ~new_n31177_;
  assign new_n31394_ = ~new_n31392_ & ~new_n31393_;
  assign new_n31395_ = new_n2965_ & ~new_n31394_;
  assign new_n31396_ = ~new_n31254_ & new_n31395_;
  assign new_n31397_ = ~new_n31390_ & ~new_n31396_;
  assign new_n31398_ = ~\b[4]  & ~new_n31397_;
  assign new_n31399_ = ~new_n31157_ & ~new_n31255_;
  assign new_n31400_ = ~new_n31168_ & new_n31172_;
  assign new_n31401_ = ~new_n31167_ & new_n31400_;
  assign new_n31402_ = ~new_n31169_ & ~new_n31172_;
  assign new_n31403_ = ~new_n31401_ & ~new_n31402_;
  assign new_n31404_ = new_n2965_ & ~new_n31403_;
  assign new_n31405_ = ~new_n31254_ & new_n31404_;
  assign new_n31406_ = ~new_n31399_ & ~new_n31405_;
  assign new_n31407_ = ~\b[3]  & ~new_n31406_;
  assign new_n31408_ = ~new_n31162_ & ~new_n31255_;
  assign new_n31409_ = new_n2873_ & ~new_n31165_;
  assign new_n31410_ = ~new_n31163_ & new_n31409_;
  assign new_n31411_ = new_n2965_ & ~new_n31410_;
  assign new_n31412_ = ~new_n31167_ & new_n31411_;
  assign new_n31413_ = ~new_n31254_ & new_n31412_;
  assign new_n31414_ = ~new_n31408_ & ~new_n31413_;
  assign new_n31415_ = ~\b[2]  & ~new_n31414_;
  assign new_n31416_ = new_n3131_ & ~new_n31254_;
  assign new_n31417_ = \a[45]  & ~new_n31416_;
  assign new_n31418_ = new_n3138_ & ~new_n31254_;
  assign new_n31419_ = ~new_n31417_ & ~new_n31418_;
  assign new_n31420_ = \b[1]  & ~new_n31419_;
  assign new_n31421_ = ~\b[1]  & ~new_n31418_;
  assign new_n31422_ = ~new_n31417_ & new_n31421_;
  assign new_n31423_ = ~new_n31420_ & ~new_n31422_;
  assign new_n31424_ = ~new_n3145_ & ~new_n31423_;
  assign new_n31425_ = ~\b[1]  & ~new_n31419_;
  assign new_n31426_ = ~new_n31424_ & ~new_n31425_;
  assign new_n31427_ = \b[2]  & ~new_n31413_;
  assign new_n31428_ = ~new_n31408_ & new_n31427_;
  assign new_n31429_ = ~new_n31415_ & ~new_n31428_;
  assign new_n31430_ = ~new_n31426_ & new_n31429_;
  assign new_n31431_ = ~new_n31415_ & ~new_n31430_;
  assign new_n31432_ = \b[3]  & ~new_n31405_;
  assign new_n31433_ = ~new_n31399_ & new_n31432_;
  assign new_n31434_ = ~new_n31407_ & ~new_n31433_;
  assign new_n31435_ = ~new_n31431_ & new_n31434_;
  assign new_n31436_ = ~new_n31407_ & ~new_n31435_;
  assign new_n31437_ = \b[4]  & ~new_n31396_;
  assign new_n31438_ = ~new_n31390_ & new_n31437_;
  assign new_n31439_ = ~new_n31398_ & ~new_n31438_;
  assign new_n31440_ = ~new_n31436_ & new_n31439_;
  assign new_n31441_ = ~new_n31398_ & ~new_n31440_;
  assign new_n31442_ = \b[5]  & ~new_n31387_;
  assign new_n31443_ = ~new_n31381_ & new_n31442_;
  assign new_n31444_ = ~new_n31389_ & ~new_n31443_;
  assign new_n31445_ = ~new_n31441_ & new_n31444_;
  assign new_n31446_ = ~new_n31389_ & ~new_n31445_;
  assign new_n31447_ = \b[6]  & ~new_n31378_;
  assign new_n31448_ = ~new_n31372_ & new_n31447_;
  assign new_n31449_ = ~new_n31380_ & ~new_n31448_;
  assign new_n31450_ = ~new_n31446_ & new_n31449_;
  assign new_n31451_ = ~new_n31380_ & ~new_n31450_;
  assign new_n31452_ = \b[7]  & ~new_n31369_;
  assign new_n31453_ = ~new_n31363_ & new_n31452_;
  assign new_n31454_ = ~new_n31371_ & ~new_n31453_;
  assign new_n31455_ = ~new_n31451_ & new_n31454_;
  assign new_n31456_ = ~new_n31371_ & ~new_n31455_;
  assign new_n31457_ = \b[8]  & ~new_n31360_;
  assign new_n31458_ = ~new_n31354_ & new_n31457_;
  assign new_n31459_ = ~new_n31362_ & ~new_n31458_;
  assign new_n31460_ = ~new_n31456_ & new_n31459_;
  assign new_n31461_ = ~new_n31362_ & ~new_n31460_;
  assign new_n31462_ = \b[9]  & ~new_n31351_;
  assign new_n31463_ = ~new_n31345_ & new_n31462_;
  assign new_n31464_ = ~new_n31353_ & ~new_n31463_;
  assign new_n31465_ = ~new_n31461_ & new_n31464_;
  assign new_n31466_ = ~new_n31353_ & ~new_n31465_;
  assign new_n31467_ = \b[10]  & ~new_n31342_;
  assign new_n31468_ = ~new_n31336_ & new_n31467_;
  assign new_n31469_ = ~new_n31344_ & ~new_n31468_;
  assign new_n31470_ = ~new_n31466_ & new_n31469_;
  assign new_n31471_ = ~new_n31344_ & ~new_n31470_;
  assign new_n31472_ = \b[11]  & ~new_n31333_;
  assign new_n31473_ = ~new_n31327_ & new_n31472_;
  assign new_n31474_ = ~new_n31335_ & ~new_n31473_;
  assign new_n31475_ = ~new_n31471_ & new_n31474_;
  assign new_n31476_ = ~new_n31335_ & ~new_n31475_;
  assign new_n31477_ = \b[12]  & ~new_n31324_;
  assign new_n31478_ = ~new_n31318_ & new_n31477_;
  assign new_n31479_ = ~new_n31326_ & ~new_n31478_;
  assign new_n31480_ = ~new_n31476_ & new_n31479_;
  assign new_n31481_ = ~new_n31326_ & ~new_n31480_;
  assign new_n31482_ = \b[13]  & ~new_n31315_;
  assign new_n31483_ = ~new_n31309_ & new_n31482_;
  assign new_n31484_ = ~new_n31317_ & ~new_n31483_;
  assign new_n31485_ = ~new_n31481_ & new_n31484_;
  assign new_n31486_ = ~new_n31317_ & ~new_n31485_;
  assign new_n31487_ = \b[14]  & ~new_n31306_;
  assign new_n31488_ = ~new_n31300_ & new_n31487_;
  assign new_n31489_ = ~new_n31308_ & ~new_n31488_;
  assign new_n31490_ = ~new_n31486_ & new_n31489_;
  assign new_n31491_ = ~new_n31308_ & ~new_n31490_;
  assign new_n31492_ = \b[15]  & ~new_n31297_;
  assign new_n31493_ = ~new_n31291_ & new_n31492_;
  assign new_n31494_ = ~new_n31299_ & ~new_n31493_;
  assign new_n31495_ = ~new_n31491_ & new_n31494_;
  assign new_n31496_ = ~new_n31299_ & ~new_n31495_;
  assign new_n31497_ = \b[16]  & ~new_n31288_;
  assign new_n31498_ = ~new_n31282_ & new_n31497_;
  assign new_n31499_ = ~new_n31290_ & ~new_n31498_;
  assign new_n31500_ = ~new_n31496_ & new_n31499_;
  assign new_n31501_ = ~new_n31290_ & ~new_n31500_;
  assign new_n31502_ = \b[17]  & ~new_n31279_;
  assign new_n31503_ = ~new_n31273_ & new_n31502_;
  assign new_n31504_ = ~new_n31281_ & ~new_n31503_;
  assign new_n31505_ = ~new_n31501_ & new_n31504_;
  assign new_n31506_ = ~new_n31281_ & ~new_n31505_;
  assign new_n31507_ = \b[18]  & ~new_n31262_;
  assign new_n31508_ = ~new_n31256_ & new_n31507_;
  assign new_n31509_ = ~new_n31272_ & ~new_n31508_;
  assign new_n31510_ = ~new_n31506_ & new_n31509_;
  assign new_n31511_ = ~new_n31272_ & ~new_n31510_;
  assign new_n31512_ = \b[19]  & ~new_n31264_;
  assign new_n31513_ = ~new_n31269_ & new_n31512_;
  assign new_n31514_ = ~new_n31271_ & ~new_n31513_;
  assign new_n31515_ = ~new_n31511_ & new_n31514_;
  assign new_n31516_ = ~new_n31271_ & ~new_n31515_;
  assign new_n31517_ = new_n320_ & ~new_n31516_;
  assign new_n31518_ = ~new_n31263_ & ~new_n31517_;
  assign new_n31519_ = ~new_n31281_ & new_n31509_;
  assign new_n31520_ = ~new_n31505_ & new_n31519_;
  assign new_n31521_ = ~new_n31506_ & ~new_n31509_;
  assign new_n31522_ = ~new_n31520_ & ~new_n31521_;
  assign new_n31523_ = new_n320_ & ~new_n31522_;
  assign new_n31524_ = ~new_n31516_ & new_n31523_;
  assign new_n31525_ = ~new_n31518_ & ~new_n31524_;
  assign new_n31526_ = ~\b[19]  & ~new_n31525_;
  assign new_n31527_ = ~new_n31280_ & ~new_n31517_;
  assign new_n31528_ = ~new_n31290_ & new_n31504_;
  assign new_n31529_ = ~new_n31500_ & new_n31528_;
  assign new_n31530_ = ~new_n31501_ & ~new_n31504_;
  assign new_n31531_ = ~new_n31529_ & ~new_n31530_;
  assign new_n31532_ = new_n320_ & ~new_n31531_;
  assign new_n31533_ = ~new_n31516_ & new_n31532_;
  assign new_n31534_ = ~new_n31527_ & ~new_n31533_;
  assign new_n31535_ = ~\b[18]  & ~new_n31534_;
  assign new_n31536_ = ~new_n31289_ & ~new_n31517_;
  assign new_n31537_ = ~new_n31299_ & new_n31499_;
  assign new_n31538_ = ~new_n31495_ & new_n31537_;
  assign new_n31539_ = ~new_n31496_ & ~new_n31499_;
  assign new_n31540_ = ~new_n31538_ & ~new_n31539_;
  assign new_n31541_ = new_n320_ & ~new_n31540_;
  assign new_n31542_ = ~new_n31516_ & new_n31541_;
  assign new_n31543_ = ~new_n31536_ & ~new_n31542_;
  assign new_n31544_ = ~\b[17]  & ~new_n31543_;
  assign new_n31545_ = ~new_n31298_ & ~new_n31517_;
  assign new_n31546_ = ~new_n31308_ & new_n31494_;
  assign new_n31547_ = ~new_n31490_ & new_n31546_;
  assign new_n31548_ = ~new_n31491_ & ~new_n31494_;
  assign new_n31549_ = ~new_n31547_ & ~new_n31548_;
  assign new_n31550_ = new_n320_ & ~new_n31549_;
  assign new_n31551_ = ~new_n31516_ & new_n31550_;
  assign new_n31552_ = ~new_n31545_ & ~new_n31551_;
  assign new_n31553_ = ~\b[16]  & ~new_n31552_;
  assign new_n31554_ = ~new_n31307_ & ~new_n31517_;
  assign new_n31555_ = ~new_n31317_ & new_n31489_;
  assign new_n31556_ = ~new_n31485_ & new_n31555_;
  assign new_n31557_ = ~new_n31486_ & ~new_n31489_;
  assign new_n31558_ = ~new_n31556_ & ~new_n31557_;
  assign new_n31559_ = new_n320_ & ~new_n31558_;
  assign new_n31560_ = ~new_n31516_ & new_n31559_;
  assign new_n31561_ = ~new_n31554_ & ~new_n31560_;
  assign new_n31562_ = ~\b[15]  & ~new_n31561_;
  assign new_n31563_ = ~new_n31316_ & ~new_n31517_;
  assign new_n31564_ = ~new_n31326_ & new_n31484_;
  assign new_n31565_ = ~new_n31480_ & new_n31564_;
  assign new_n31566_ = ~new_n31481_ & ~new_n31484_;
  assign new_n31567_ = ~new_n31565_ & ~new_n31566_;
  assign new_n31568_ = new_n320_ & ~new_n31567_;
  assign new_n31569_ = ~new_n31516_ & new_n31568_;
  assign new_n31570_ = ~new_n31563_ & ~new_n31569_;
  assign new_n31571_ = ~\b[14]  & ~new_n31570_;
  assign new_n31572_ = ~new_n31325_ & ~new_n31517_;
  assign new_n31573_ = ~new_n31335_ & new_n31479_;
  assign new_n31574_ = ~new_n31475_ & new_n31573_;
  assign new_n31575_ = ~new_n31476_ & ~new_n31479_;
  assign new_n31576_ = ~new_n31574_ & ~new_n31575_;
  assign new_n31577_ = new_n320_ & ~new_n31576_;
  assign new_n31578_ = ~new_n31516_ & new_n31577_;
  assign new_n31579_ = ~new_n31572_ & ~new_n31578_;
  assign new_n31580_ = ~\b[13]  & ~new_n31579_;
  assign new_n31581_ = ~new_n31334_ & ~new_n31517_;
  assign new_n31582_ = ~new_n31344_ & new_n31474_;
  assign new_n31583_ = ~new_n31470_ & new_n31582_;
  assign new_n31584_ = ~new_n31471_ & ~new_n31474_;
  assign new_n31585_ = ~new_n31583_ & ~new_n31584_;
  assign new_n31586_ = new_n320_ & ~new_n31585_;
  assign new_n31587_ = ~new_n31516_ & new_n31586_;
  assign new_n31588_ = ~new_n31581_ & ~new_n31587_;
  assign new_n31589_ = ~\b[12]  & ~new_n31588_;
  assign new_n31590_ = ~new_n31343_ & ~new_n31517_;
  assign new_n31591_ = ~new_n31353_ & new_n31469_;
  assign new_n31592_ = ~new_n31465_ & new_n31591_;
  assign new_n31593_ = ~new_n31466_ & ~new_n31469_;
  assign new_n31594_ = ~new_n31592_ & ~new_n31593_;
  assign new_n31595_ = new_n320_ & ~new_n31594_;
  assign new_n31596_ = ~new_n31516_ & new_n31595_;
  assign new_n31597_ = ~new_n31590_ & ~new_n31596_;
  assign new_n31598_ = ~\b[11]  & ~new_n31597_;
  assign new_n31599_ = ~new_n31352_ & ~new_n31517_;
  assign new_n31600_ = ~new_n31362_ & new_n31464_;
  assign new_n31601_ = ~new_n31460_ & new_n31600_;
  assign new_n31602_ = ~new_n31461_ & ~new_n31464_;
  assign new_n31603_ = ~new_n31601_ & ~new_n31602_;
  assign new_n31604_ = new_n320_ & ~new_n31603_;
  assign new_n31605_ = ~new_n31516_ & new_n31604_;
  assign new_n31606_ = ~new_n31599_ & ~new_n31605_;
  assign new_n31607_ = ~\b[10]  & ~new_n31606_;
  assign new_n31608_ = ~new_n31361_ & ~new_n31517_;
  assign new_n31609_ = ~new_n31371_ & new_n31459_;
  assign new_n31610_ = ~new_n31455_ & new_n31609_;
  assign new_n31611_ = ~new_n31456_ & ~new_n31459_;
  assign new_n31612_ = ~new_n31610_ & ~new_n31611_;
  assign new_n31613_ = new_n320_ & ~new_n31612_;
  assign new_n31614_ = ~new_n31516_ & new_n31613_;
  assign new_n31615_ = ~new_n31608_ & ~new_n31614_;
  assign new_n31616_ = ~\b[9]  & ~new_n31615_;
  assign new_n31617_ = ~new_n31370_ & ~new_n31517_;
  assign new_n31618_ = ~new_n31380_ & new_n31454_;
  assign new_n31619_ = ~new_n31450_ & new_n31618_;
  assign new_n31620_ = ~new_n31451_ & ~new_n31454_;
  assign new_n31621_ = ~new_n31619_ & ~new_n31620_;
  assign new_n31622_ = new_n320_ & ~new_n31621_;
  assign new_n31623_ = ~new_n31516_ & new_n31622_;
  assign new_n31624_ = ~new_n31617_ & ~new_n31623_;
  assign new_n31625_ = ~\b[8]  & ~new_n31624_;
  assign new_n31626_ = ~new_n31379_ & ~new_n31517_;
  assign new_n31627_ = ~new_n31389_ & new_n31449_;
  assign new_n31628_ = ~new_n31445_ & new_n31627_;
  assign new_n31629_ = ~new_n31446_ & ~new_n31449_;
  assign new_n31630_ = ~new_n31628_ & ~new_n31629_;
  assign new_n31631_ = new_n320_ & ~new_n31630_;
  assign new_n31632_ = ~new_n31516_ & new_n31631_;
  assign new_n31633_ = ~new_n31626_ & ~new_n31632_;
  assign new_n31634_ = ~\b[7]  & ~new_n31633_;
  assign new_n31635_ = ~new_n31388_ & ~new_n31517_;
  assign new_n31636_ = ~new_n31398_ & new_n31444_;
  assign new_n31637_ = ~new_n31440_ & new_n31636_;
  assign new_n31638_ = ~new_n31441_ & ~new_n31444_;
  assign new_n31639_ = ~new_n31637_ & ~new_n31638_;
  assign new_n31640_ = new_n320_ & ~new_n31639_;
  assign new_n31641_ = ~new_n31516_ & new_n31640_;
  assign new_n31642_ = ~new_n31635_ & ~new_n31641_;
  assign new_n31643_ = ~\b[6]  & ~new_n31642_;
  assign new_n31644_ = ~new_n31397_ & ~new_n31517_;
  assign new_n31645_ = ~new_n31407_ & new_n31439_;
  assign new_n31646_ = ~new_n31435_ & new_n31645_;
  assign new_n31647_ = ~new_n31436_ & ~new_n31439_;
  assign new_n31648_ = ~new_n31646_ & ~new_n31647_;
  assign new_n31649_ = new_n320_ & ~new_n31648_;
  assign new_n31650_ = ~new_n31516_ & new_n31649_;
  assign new_n31651_ = ~new_n31644_ & ~new_n31650_;
  assign new_n31652_ = ~\b[5]  & ~new_n31651_;
  assign new_n31653_ = ~new_n31406_ & ~new_n31517_;
  assign new_n31654_ = ~new_n31415_ & new_n31434_;
  assign new_n31655_ = ~new_n31430_ & new_n31654_;
  assign new_n31656_ = ~new_n31431_ & ~new_n31434_;
  assign new_n31657_ = ~new_n31655_ & ~new_n31656_;
  assign new_n31658_ = new_n320_ & ~new_n31657_;
  assign new_n31659_ = ~new_n31516_ & new_n31658_;
  assign new_n31660_ = ~new_n31653_ & ~new_n31659_;
  assign new_n31661_ = ~\b[4]  & ~new_n31660_;
  assign new_n31662_ = ~new_n31414_ & ~new_n31517_;
  assign new_n31663_ = ~new_n31425_ & new_n31429_;
  assign new_n31664_ = ~new_n31424_ & new_n31663_;
  assign new_n31665_ = ~new_n31426_ & ~new_n31429_;
  assign new_n31666_ = ~new_n31664_ & ~new_n31665_;
  assign new_n31667_ = new_n320_ & ~new_n31666_;
  assign new_n31668_ = ~new_n31516_ & new_n31667_;
  assign new_n31669_ = ~new_n31662_ & ~new_n31668_;
  assign new_n31670_ = ~\b[3]  & ~new_n31669_;
  assign new_n31671_ = ~new_n31419_ & ~new_n31517_;
  assign new_n31672_ = new_n3145_ & ~new_n31422_;
  assign new_n31673_ = ~new_n31420_ & new_n31672_;
  assign new_n31674_ = new_n320_ & ~new_n31673_;
  assign new_n31675_ = ~new_n31424_ & new_n31674_;
  assign new_n31676_ = ~new_n31516_ & new_n31675_;
  assign new_n31677_ = ~new_n31671_ & ~new_n31676_;
  assign new_n31678_ = ~\b[2]  & ~new_n31677_;
  assign new_n31679_ = new_n3405_ & ~new_n31516_;
  assign new_n31680_ = \a[44]  & ~new_n31679_;
  assign new_n31681_ = new_n3411_ & ~new_n31516_;
  assign new_n31682_ = ~new_n31680_ & ~new_n31681_;
  assign new_n31683_ = \b[1]  & ~new_n31682_;
  assign new_n31684_ = ~\b[1]  & ~new_n31681_;
  assign new_n31685_ = ~new_n31680_ & new_n31684_;
  assign new_n31686_ = ~new_n31683_ & ~new_n31685_;
  assign new_n31687_ = ~new_n3418_ & ~new_n31686_;
  assign new_n31688_ = ~\b[1]  & ~new_n31682_;
  assign new_n31689_ = ~new_n31687_ & ~new_n31688_;
  assign new_n31690_ = \b[2]  & ~new_n31676_;
  assign new_n31691_ = ~new_n31671_ & new_n31690_;
  assign new_n31692_ = ~new_n31678_ & ~new_n31691_;
  assign new_n31693_ = ~new_n31689_ & new_n31692_;
  assign new_n31694_ = ~new_n31678_ & ~new_n31693_;
  assign new_n31695_ = \b[3]  & ~new_n31668_;
  assign new_n31696_ = ~new_n31662_ & new_n31695_;
  assign new_n31697_ = ~new_n31670_ & ~new_n31696_;
  assign new_n31698_ = ~new_n31694_ & new_n31697_;
  assign new_n31699_ = ~new_n31670_ & ~new_n31698_;
  assign new_n31700_ = \b[4]  & ~new_n31659_;
  assign new_n31701_ = ~new_n31653_ & new_n31700_;
  assign new_n31702_ = ~new_n31661_ & ~new_n31701_;
  assign new_n31703_ = ~new_n31699_ & new_n31702_;
  assign new_n31704_ = ~new_n31661_ & ~new_n31703_;
  assign new_n31705_ = \b[5]  & ~new_n31650_;
  assign new_n31706_ = ~new_n31644_ & new_n31705_;
  assign new_n31707_ = ~new_n31652_ & ~new_n31706_;
  assign new_n31708_ = ~new_n31704_ & new_n31707_;
  assign new_n31709_ = ~new_n31652_ & ~new_n31708_;
  assign new_n31710_ = \b[6]  & ~new_n31641_;
  assign new_n31711_ = ~new_n31635_ & new_n31710_;
  assign new_n31712_ = ~new_n31643_ & ~new_n31711_;
  assign new_n31713_ = ~new_n31709_ & new_n31712_;
  assign new_n31714_ = ~new_n31643_ & ~new_n31713_;
  assign new_n31715_ = \b[7]  & ~new_n31632_;
  assign new_n31716_ = ~new_n31626_ & new_n31715_;
  assign new_n31717_ = ~new_n31634_ & ~new_n31716_;
  assign new_n31718_ = ~new_n31714_ & new_n31717_;
  assign new_n31719_ = ~new_n31634_ & ~new_n31718_;
  assign new_n31720_ = \b[8]  & ~new_n31623_;
  assign new_n31721_ = ~new_n31617_ & new_n31720_;
  assign new_n31722_ = ~new_n31625_ & ~new_n31721_;
  assign new_n31723_ = ~new_n31719_ & new_n31722_;
  assign new_n31724_ = ~new_n31625_ & ~new_n31723_;
  assign new_n31725_ = \b[9]  & ~new_n31614_;
  assign new_n31726_ = ~new_n31608_ & new_n31725_;
  assign new_n31727_ = ~new_n31616_ & ~new_n31726_;
  assign new_n31728_ = ~new_n31724_ & new_n31727_;
  assign new_n31729_ = ~new_n31616_ & ~new_n31728_;
  assign new_n31730_ = \b[10]  & ~new_n31605_;
  assign new_n31731_ = ~new_n31599_ & new_n31730_;
  assign new_n31732_ = ~new_n31607_ & ~new_n31731_;
  assign new_n31733_ = ~new_n31729_ & new_n31732_;
  assign new_n31734_ = ~new_n31607_ & ~new_n31733_;
  assign new_n31735_ = \b[11]  & ~new_n31596_;
  assign new_n31736_ = ~new_n31590_ & new_n31735_;
  assign new_n31737_ = ~new_n31598_ & ~new_n31736_;
  assign new_n31738_ = ~new_n31734_ & new_n31737_;
  assign new_n31739_ = ~new_n31598_ & ~new_n31738_;
  assign new_n31740_ = \b[12]  & ~new_n31587_;
  assign new_n31741_ = ~new_n31581_ & new_n31740_;
  assign new_n31742_ = ~new_n31589_ & ~new_n31741_;
  assign new_n31743_ = ~new_n31739_ & new_n31742_;
  assign new_n31744_ = ~new_n31589_ & ~new_n31743_;
  assign new_n31745_ = \b[13]  & ~new_n31578_;
  assign new_n31746_ = ~new_n31572_ & new_n31745_;
  assign new_n31747_ = ~new_n31580_ & ~new_n31746_;
  assign new_n31748_ = ~new_n31744_ & new_n31747_;
  assign new_n31749_ = ~new_n31580_ & ~new_n31748_;
  assign new_n31750_ = \b[14]  & ~new_n31569_;
  assign new_n31751_ = ~new_n31563_ & new_n31750_;
  assign new_n31752_ = ~new_n31571_ & ~new_n31751_;
  assign new_n31753_ = ~new_n31749_ & new_n31752_;
  assign new_n31754_ = ~new_n31571_ & ~new_n31753_;
  assign new_n31755_ = \b[15]  & ~new_n31560_;
  assign new_n31756_ = ~new_n31554_ & new_n31755_;
  assign new_n31757_ = ~new_n31562_ & ~new_n31756_;
  assign new_n31758_ = ~new_n31754_ & new_n31757_;
  assign new_n31759_ = ~new_n31562_ & ~new_n31758_;
  assign new_n31760_ = \b[16]  & ~new_n31551_;
  assign new_n31761_ = ~new_n31545_ & new_n31760_;
  assign new_n31762_ = ~new_n31553_ & ~new_n31761_;
  assign new_n31763_ = ~new_n31759_ & new_n31762_;
  assign new_n31764_ = ~new_n31553_ & ~new_n31763_;
  assign new_n31765_ = \b[17]  & ~new_n31542_;
  assign new_n31766_ = ~new_n31536_ & new_n31765_;
  assign new_n31767_ = ~new_n31544_ & ~new_n31766_;
  assign new_n31768_ = ~new_n31764_ & new_n31767_;
  assign new_n31769_ = ~new_n31544_ & ~new_n31768_;
  assign new_n31770_ = \b[18]  & ~new_n31533_;
  assign new_n31771_ = ~new_n31527_ & new_n31770_;
  assign new_n31772_ = ~new_n31535_ & ~new_n31771_;
  assign new_n31773_ = ~new_n31769_ & new_n31772_;
  assign new_n31774_ = ~new_n31535_ & ~new_n31773_;
  assign new_n31775_ = \b[19]  & ~new_n31524_;
  assign new_n31776_ = ~new_n31518_ & new_n31775_;
  assign new_n31777_ = ~new_n31526_ & ~new_n31776_;
  assign new_n31778_ = ~new_n31774_ & new_n31777_;
  assign new_n31779_ = ~new_n31526_ & ~new_n31778_;
  assign new_n31780_ = ~new_n31270_ & ~new_n31517_;
  assign new_n31781_ = ~new_n31272_ & new_n31514_;
  assign new_n31782_ = ~new_n31510_ & new_n31781_;
  assign new_n31783_ = ~new_n31511_ & ~new_n31514_;
  assign new_n31784_ = ~new_n31782_ & ~new_n31783_;
  assign new_n31785_ = new_n31517_ & ~new_n31784_;
  assign new_n31786_ = ~new_n31780_ & ~new_n31785_;
  assign new_n31787_ = ~\b[20]  & ~new_n31786_;
  assign new_n31788_ = \b[20]  & ~new_n31780_;
  assign new_n31789_ = ~new_n31785_ & new_n31788_;
  assign new_n31790_ = new_n643_ & ~new_n31789_;
  assign new_n31791_ = ~new_n31787_ & new_n31790_;
  assign new_n31792_ = ~new_n31779_ & new_n31791_;
  assign new_n31793_ = new_n320_ & ~new_n31786_;
  assign new_n31794_ = ~new_n31792_ & ~new_n31793_;
  assign new_n31795_ = ~new_n31535_ & new_n31777_;
  assign new_n31796_ = ~new_n31773_ & new_n31795_;
  assign new_n31797_ = ~new_n31774_ & ~new_n31777_;
  assign new_n31798_ = ~new_n31796_ & ~new_n31797_;
  assign new_n31799_ = ~new_n31794_ & ~new_n31798_;
  assign new_n31800_ = ~new_n31525_ & ~new_n31793_;
  assign new_n31801_ = ~new_n31792_ & new_n31800_;
  assign new_n31802_ = ~new_n31799_ & ~new_n31801_;
  assign new_n31803_ = ~new_n31526_ & ~new_n31789_;
  assign new_n31804_ = ~new_n31787_ & new_n31803_;
  assign new_n31805_ = ~new_n31778_ & new_n31804_;
  assign new_n31806_ = ~new_n31787_ & ~new_n31789_;
  assign new_n31807_ = ~new_n31779_ & ~new_n31806_;
  assign new_n31808_ = ~new_n31805_ & ~new_n31807_;
  assign new_n31809_ = ~new_n31794_ & ~new_n31808_;
  assign new_n31810_ = ~new_n31786_ & ~new_n31793_;
  assign new_n31811_ = ~new_n31792_ & new_n31810_;
  assign new_n31812_ = ~new_n31809_ & ~new_n31811_;
  assign new_n31813_ = ~\b[21]  & ~new_n31812_;
  assign new_n31814_ = ~\b[20]  & ~new_n31802_;
  assign new_n31815_ = ~new_n31544_ & new_n31772_;
  assign new_n31816_ = ~new_n31768_ & new_n31815_;
  assign new_n31817_ = ~new_n31769_ & ~new_n31772_;
  assign new_n31818_ = ~new_n31816_ & ~new_n31817_;
  assign new_n31819_ = ~new_n31794_ & ~new_n31818_;
  assign new_n31820_ = ~new_n31534_ & ~new_n31793_;
  assign new_n31821_ = ~new_n31792_ & new_n31820_;
  assign new_n31822_ = ~new_n31819_ & ~new_n31821_;
  assign new_n31823_ = ~\b[19]  & ~new_n31822_;
  assign new_n31824_ = ~new_n31553_ & new_n31767_;
  assign new_n31825_ = ~new_n31763_ & new_n31824_;
  assign new_n31826_ = ~new_n31764_ & ~new_n31767_;
  assign new_n31827_ = ~new_n31825_ & ~new_n31826_;
  assign new_n31828_ = ~new_n31794_ & ~new_n31827_;
  assign new_n31829_ = ~new_n31543_ & ~new_n31793_;
  assign new_n31830_ = ~new_n31792_ & new_n31829_;
  assign new_n31831_ = ~new_n31828_ & ~new_n31830_;
  assign new_n31832_ = ~\b[18]  & ~new_n31831_;
  assign new_n31833_ = ~new_n31562_ & new_n31762_;
  assign new_n31834_ = ~new_n31758_ & new_n31833_;
  assign new_n31835_ = ~new_n31759_ & ~new_n31762_;
  assign new_n31836_ = ~new_n31834_ & ~new_n31835_;
  assign new_n31837_ = ~new_n31794_ & ~new_n31836_;
  assign new_n31838_ = ~new_n31552_ & ~new_n31793_;
  assign new_n31839_ = ~new_n31792_ & new_n31838_;
  assign new_n31840_ = ~new_n31837_ & ~new_n31839_;
  assign new_n31841_ = ~\b[17]  & ~new_n31840_;
  assign new_n31842_ = ~new_n31571_ & new_n31757_;
  assign new_n31843_ = ~new_n31753_ & new_n31842_;
  assign new_n31844_ = ~new_n31754_ & ~new_n31757_;
  assign new_n31845_ = ~new_n31843_ & ~new_n31844_;
  assign new_n31846_ = ~new_n31794_ & ~new_n31845_;
  assign new_n31847_ = ~new_n31561_ & ~new_n31793_;
  assign new_n31848_ = ~new_n31792_ & new_n31847_;
  assign new_n31849_ = ~new_n31846_ & ~new_n31848_;
  assign new_n31850_ = ~\b[16]  & ~new_n31849_;
  assign new_n31851_ = ~new_n31580_ & new_n31752_;
  assign new_n31852_ = ~new_n31748_ & new_n31851_;
  assign new_n31853_ = ~new_n31749_ & ~new_n31752_;
  assign new_n31854_ = ~new_n31852_ & ~new_n31853_;
  assign new_n31855_ = ~new_n31794_ & ~new_n31854_;
  assign new_n31856_ = ~new_n31570_ & ~new_n31793_;
  assign new_n31857_ = ~new_n31792_ & new_n31856_;
  assign new_n31858_ = ~new_n31855_ & ~new_n31857_;
  assign new_n31859_ = ~\b[15]  & ~new_n31858_;
  assign new_n31860_ = ~new_n31589_ & new_n31747_;
  assign new_n31861_ = ~new_n31743_ & new_n31860_;
  assign new_n31862_ = ~new_n31744_ & ~new_n31747_;
  assign new_n31863_ = ~new_n31861_ & ~new_n31862_;
  assign new_n31864_ = ~new_n31794_ & ~new_n31863_;
  assign new_n31865_ = ~new_n31579_ & ~new_n31793_;
  assign new_n31866_ = ~new_n31792_ & new_n31865_;
  assign new_n31867_ = ~new_n31864_ & ~new_n31866_;
  assign new_n31868_ = ~\b[14]  & ~new_n31867_;
  assign new_n31869_ = ~new_n31598_ & new_n31742_;
  assign new_n31870_ = ~new_n31738_ & new_n31869_;
  assign new_n31871_ = ~new_n31739_ & ~new_n31742_;
  assign new_n31872_ = ~new_n31870_ & ~new_n31871_;
  assign new_n31873_ = ~new_n31794_ & ~new_n31872_;
  assign new_n31874_ = ~new_n31588_ & ~new_n31793_;
  assign new_n31875_ = ~new_n31792_ & new_n31874_;
  assign new_n31876_ = ~new_n31873_ & ~new_n31875_;
  assign new_n31877_ = ~\b[13]  & ~new_n31876_;
  assign new_n31878_ = ~new_n31607_ & new_n31737_;
  assign new_n31879_ = ~new_n31733_ & new_n31878_;
  assign new_n31880_ = ~new_n31734_ & ~new_n31737_;
  assign new_n31881_ = ~new_n31879_ & ~new_n31880_;
  assign new_n31882_ = ~new_n31794_ & ~new_n31881_;
  assign new_n31883_ = ~new_n31597_ & ~new_n31793_;
  assign new_n31884_ = ~new_n31792_ & new_n31883_;
  assign new_n31885_ = ~new_n31882_ & ~new_n31884_;
  assign new_n31886_ = ~\b[12]  & ~new_n31885_;
  assign new_n31887_ = ~new_n31616_ & new_n31732_;
  assign new_n31888_ = ~new_n31728_ & new_n31887_;
  assign new_n31889_ = ~new_n31729_ & ~new_n31732_;
  assign new_n31890_ = ~new_n31888_ & ~new_n31889_;
  assign new_n31891_ = ~new_n31794_ & ~new_n31890_;
  assign new_n31892_ = ~new_n31606_ & ~new_n31793_;
  assign new_n31893_ = ~new_n31792_ & new_n31892_;
  assign new_n31894_ = ~new_n31891_ & ~new_n31893_;
  assign new_n31895_ = ~\b[11]  & ~new_n31894_;
  assign new_n31896_ = ~new_n31625_ & new_n31727_;
  assign new_n31897_ = ~new_n31723_ & new_n31896_;
  assign new_n31898_ = ~new_n31724_ & ~new_n31727_;
  assign new_n31899_ = ~new_n31897_ & ~new_n31898_;
  assign new_n31900_ = ~new_n31794_ & ~new_n31899_;
  assign new_n31901_ = ~new_n31615_ & ~new_n31793_;
  assign new_n31902_ = ~new_n31792_ & new_n31901_;
  assign new_n31903_ = ~new_n31900_ & ~new_n31902_;
  assign new_n31904_ = ~\b[10]  & ~new_n31903_;
  assign new_n31905_ = ~new_n31634_ & new_n31722_;
  assign new_n31906_ = ~new_n31718_ & new_n31905_;
  assign new_n31907_ = ~new_n31719_ & ~new_n31722_;
  assign new_n31908_ = ~new_n31906_ & ~new_n31907_;
  assign new_n31909_ = ~new_n31794_ & ~new_n31908_;
  assign new_n31910_ = ~new_n31624_ & ~new_n31793_;
  assign new_n31911_ = ~new_n31792_ & new_n31910_;
  assign new_n31912_ = ~new_n31909_ & ~new_n31911_;
  assign new_n31913_ = ~\b[9]  & ~new_n31912_;
  assign new_n31914_ = ~new_n31643_ & new_n31717_;
  assign new_n31915_ = ~new_n31713_ & new_n31914_;
  assign new_n31916_ = ~new_n31714_ & ~new_n31717_;
  assign new_n31917_ = ~new_n31915_ & ~new_n31916_;
  assign new_n31918_ = ~new_n31794_ & ~new_n31917_;
  assign new_n31919_ = ~new_n31633_ & ~new_n31793_;
  assign new_n31920_ = ~new_n31792_ & new_n31919_;
  assign new_n31921_ = ~new_n31918_ & ~new_n31920_;
  assign new_n31922_ = ~\b[8]  & ~new_n31921_;
  assign new_n31923_ = ~new_n31652_ & new_n31712_;
  assign new_n31924_ = ~new_n31708_ & new_n31923_;
  assign new_n31925_ = ~new_n31709_ & ~new_n31712_;
  assign new_n31926_ = ~new_n31924_ & ~new_n31925_;
  assign new_n31927_ = ~new_n31794_ & ~new_n31926_;
  assign new_n31928_ = ~new_n31642_ & ~new_n31793_;
  assign new_n31929_ = ~new_n31792_ & new_n31928_;
  assign new_n31930_ = ~new_n31927_ & ~new_n31929_;
  assign new_n31931_ = ~\b[7]  & ~new_n31930_;
  assign new_n31932_ = ~new_n31661_ & new_n31707_;
  assign new_n31933_ = ~new_n31703_ & new_n31932_;
  assign new_n31934_ = ~new_n31704_ & ~new_n31707_;
  assign new_n31935_ = ~new_n31933_ & ~new_n31934_;
  assign new_n31936_ = ~new_n31794_ & ~new_n31935_;
  assign new_n31937_ = ~new_n31651_ & ~new_n31793_;
  assign new_n31938_ = ~new_n31792_ & new_n31937_;
  assign new_n31939_ = ~new_n31936_ & ~new_n31938_;
  assign new_n31940_ = ~\b[6]  & ~new_n31939_;
  assign new_n31941_ = ~new_n31670_ & new_n31702_;
  assign new_n31942_ = ~new_n31698_ & new_n31941_;
  assign new_n31943_ = ~new_n31699_ & ~new_n31702_;
  assign new_n31944_ = ~new_n31942_ & ~new_n31943_;
  assign new_n31945_ = ~new_n31794_ & ~new_n31944_;
  assign new_n31946_ = ~new_n31660_ & ~new_n31793_;
  assign new_n31947_ = ~new_n31792_ & new_n31946_;
  assign new_n31948_ = ~new_n31945_ & ~new_n31947_;
  assign new_n31949_ = ~\b[5]  & ~new_n31948_;
  assign new_n31950_ = ~new_n31678_ & new_n31697_;
  assign new_n31951_ = ~new_n31693_ & new_n31950_;
  assign new_n31952_ = ~new_n31694_ & ~new_n31697_;
  assign new_n31953_ = ~new_n31951_ & ~new_n31952_;
  assign new_n31954_ = ~new_n31794_ & ~new_n31953_;
  assign new_n31955_ = ~new_n31669_ & ~new_n31793_;
  assign new_n31956_ = ~new_n31792_ & new_n31955_;
  assign new_n31957_ = ~new_n31954_ & ~new_n31956_;
  assign new_n31958_ = ~\b[4]  & ~new_n31957_;
  assign new_n31959_ = ~new_n31688_ & new_n31692_;
  assign new_n31960_ = ~new_n31687_ & new_n31959_;
  assign new_n31961_ = ~new_n31689_ & ~new_n31692_;
  assign new_n31962_ = ~new_n31960_ & ~new_n31961_;
  assign new_n31963_ = ~new_n31794_ & ~new_n31962_;
  assign new_n31964_ = ~new_n31677_ & ~new_n31793_;
  assign new_n31965_ = ~new_n31792_ & new_n31964_;
  assign new_n31966_ = ~new_n31963_ & ~new_n31965_;
  assign new_n31967_ = ~\b[3]  & ~new_n31966_;
  assign new_n31968_ = new_n3418_ & ~new_n31685_;
  assign new_n31969_ = ~new_n31683_ & new_n31968_;
  assign new_n31970_ = ~new_n31687_ & ~new_n31969_;
  assign new_n31971_ = ~new_n31794_ & new_n31970_;
  assign new_n31972_ = ~new_n31682_ & ~new_n31793_;
  assign new_n31973_ = ~new_n31792_ & new_n31972_;
  assign new_n31974_ = ~new_n31971_ & ~new_n31973_;
  assign new_n31975_ = ~\b[2]  & ~new_n31974_;
  assign new_n31976_ = \b[0]  & ~new_n31794_;
  assign new_n31977_ = \a[43]  & ~new_n31976_;
  assign new_n31978_ = new_n3418_ & ~new_n31794_;
  assign new_n31979_ = ~new_n31977_ & ~new_n31978_;
  assign new_n31980_ = \b[1]  & ~new_n31979_;
  assign new_n31981_ = ~\b[1]  & ~new_n31978_;
  assign new_n31982_ = ~new_n31977_ & new_n31981_;
  assign new_n31983_ = ~new_n31980_ & ~new_n31982_;
  assign new_n31984_ = ~new_n3716_ & ~new_n31983_;
  assign new_n31985_ = ~\b[1]  & ~new_n31979_;
  assign new_n31986_ = ~new_n31984_ & ~new_n31985_;
  assign new_n31987_ = \b[2]  & ~new_n31973_;
  assign new_n31988_ = ~new_n31971_ & new_n31987_;
  assign new_n31989_ = ~new_n31975_ & ~new_n31988_;
  assign new_n31990_ = ~new_n31986_ & new_n31989_;
  assign new_n31991_ = ~new_n31975_ & ~new_n31990_;
  assign new_n31992_ = \b[3]  & ~new_n31965_;
  assign new_n31993_ = ~new_n31963_ & new_n31992_;
  assign new_n31994_ = ~new_n31967_ & ~new_n31993_;
  assign new_n31995_ = ~new_n31991_ & new_n31994_;
  assign new_n31996_ = ~new_n31967_ & ~new_n31995_;
  assign new_n31997_ = \b[4]  & ~new_n31956_;
  assign new_n31998_ = ~new_n31954_ & new_n31997_;
  assign new_n31999_ = ~new_n31958_ & ~new_n31998_;
  assign new_n32000_ = ~new_n31996_ & new_n31999_;
  assign new_n32001_ = ~new_n31958_ & ~new_n32000_;
  assign new_n32002_ = \b[5]  & ~new_n31947_;
  assign new_n32003_ = ~new_n31945_ & new_n32002_;
  assign new_n32004_ = ~new_n31949_ & ~new_n32003_;
  assign new_n32005_ = ~new_n32001_ & new_n32004_;
  assign new_n32006_ = ~new_n31949_ & ~new_n32005_;
  assign new_n32007_ = \b[6]  & ~new_n31938_;
  assign new_n32008_ = ~new_n31936_ & new_n32007_;
  assign new_n32009_ = ~new_n31940_ & ~new_n32008_;
  assign new_n32010_ = ~new_n32006_ & new_n32009_;
  assign new_n32011_ = ~new_n31940_ & ~new_n32010_;
  assign new_n32012_ = \b[7]  & ~new_n31929_;
  assign new_n32013_ = ~new_n31927_ & new_n32012_;
  assign new_n32014_ = ~new_n31931_ & ~new_n32013_;
  assign new_n32015_ = ~new_n32011_ & new_n32014_;
  assign new_n32016_ = ~new_n31931_ & ~new_n32015_;
  assign new_n32017_ = \b[8]  & ~new_n31920_;
  assign new_n32018_ = ~new_n31918_ & new_n32017_;
  assign new_n32019_ = ~new_n31922_ & ~new_n32018_;
  assign new_n32020_ = ~new_n32016_ & new_n32019_;
  assign new_n32021_ = ~new_n31922_ & ~new_n32020_;
  assign new_n32022_ = \b[9]  & ~new_n31911_;
  assign new_n32023_ = ~new_n31909_ & new_n32022_;
  assign new_n32024_ = ~new_n31913_ & ~new_n32023_;
  assign new_n32025_ = ~new_n32021_ & new_n32024_;
  assign new_n32026_ = ~new_n31913_ & ~new_n32025_;
  assign new_n32027_ = \b[10]  & ~new_n31902_;
  assign new_n32028_ = ~new_n31900_ & new_n32027_;
  assign new_n32029_ = ~new_n31904_ & ~new_n32028_;
  assign new_n32030_ = ~new_n32026_ & new_n32029_;
  assign new_n32031_ = ~new_n31904_ & ~new_n32030_;
  assign new_n32032_ = \b[11]  & ~new_n31893_;
  assign new_n32033_ = ~new_n31891_ & new_n32032_;
  assign new_n32034_ = ~new_n31895_ & ~new_n32033_;
  assign new_n32035_ = ~new_n32031_ & new_n32034_;
  assign new_n32036_ = ~new_n31895_ & ~new_n32035_;
  assign new_n32037_ = \b[12]  & ~new_n31884_;
  assign new_n32038_ = ~new_n31882_ & new_n32037_;
  assign new_n32039_ = ~new_n31886_ & ~new_n32038_;
  assign new_n32040_ = ~new_n32036_ & new_n32039_;
  assign new_n32041_ = ~new_n31886_ & ~new_n32040_;
  assign new_n32042_ = \b[13]  & ~new_n31875_;
  assign new_n32043_ = ~new_n31873_ & new_n32042_;
  assign new_n32044_ = ~new_n31877_ & ~new_n32043_;
  assign new_n32045_ = ~new_n32041_ & new_n32044_;
  assign new_n32046_ = ~new_n31877_ & ~new_n32045_;
  assign new_n32047_ = \b[14]  & ~new_n31866_;
  assign new_n32048_ = ~new_n31864_ & new_n32047_;
  assign new_n32049_ = ~new_n31868_ & ~new_n32048_;
  assign new_n32050_ = ~new_n32046_ & new_n32049_;
  assign new_n32051_ = ~new_n31868_ & ~new_n32050_;
  assign new_n32052_ = \b[15]  & ~new_n31857_;
  assign new_n32053_ = ~new_n31855_ & new_n32052_;
  assign new_n32054_ = ~new_n31859_ & ~new_n32053_;
  assign new_n32055_ = ~new_n32051_ & new_n32054_;
  assign new_n32056_ = ~new_n31859_ & ~new_n32055_;
  assign new_n32057_ = \b[16]  & ~new_n31848_;
  assign new_n32058_ = ~new_n31846_ & new_n32057_;
  assign new_n32059_ = ~new_n31850_ & ~new_n32058_;
  assign new_n32060_ = ~new_n32056_ & new_n32059_;
  assign new_n32061_ = ~new_n31850_ & ~new_n32060_;
  assign new_n32062_ = \b[17]  & ~new_n31839_;
  assign new_n32063_ = ~new_n31837_ & new_n32062_;
  assign new_n32064_ = ~new_n31841_ & ~new_n32063_;
  assign new_n32065_ = ~new_n32061_ & new_n32064_;
  assign new_n32066_ = ~new_n31841_ & ~new_n32065_;
  assign new_n32067_ = \b[18]  & ~new_n31830_;
  assign new_n32068_ = ~new_n31828_ & new_n32067_;
  assign new_n32069_ = ~new_n31832_ & ~new_n32068_;
  assign new_n32070_ = ~new_n32066_ & new_n32069_;
  assign new_n32071_ = ~new_n31832_ & ~new_n32070_;
  assign new_n32072_ = \b[19]  & ~new_n31821_;
  assign new_n32073_ = ~new_n31819_ & new_n32072_;
  assign new_n32074_ = ~new_n31823_ & ~new_n32073_;
  assign new_n32075_ = ~new_n32071_ & new_n32074_;
  assign new_n32076_ = ~new_n31823_ & ~new_n32075_;
  assign new_n32077_ = \b[20]  & ~new_n31801_;
  assign new_n32078_ = ~new_n31799_ & new_n32077_;
  assign new_n32079_ = ~new_n31814_ & ~new_n32078_;
  assign new_n32080_ = ~new_n32076_ & new_n32079_;
  assign new_n32081_ = ~new_n31814_ & ~new_n32080_;
  assign new_n32082_ = \b[21]  & ~new_n31811_;
  assign new_n32083_ = ~new_n31809_ & new_n32082_;
  assign new_n32084_ = ~new_n31813_ & ~new_n32083_;
  assign new_n32085_ = ~new_n32081_ & new_n32084_;
  assign new_n32086_ = ~new_n31813_ & ~new_n32085_;
  assign new_n32087_ = new_n3823_ & ~new_n32086_;
  assign new_n32088_ = ~new_n31802_ & ~new_n32087_;
  assign new_n32089_ = ~new_n31823_ & new_n32079_;
  assign new_n32090_ = ~new_n32075_ & new_n32089_;
  assign new_n32091_ = ~new_n32076_ & ~new_n32079_;
  assign new_n32092_ = ~new_n32090_ & ~new_n32091_;
  assign new_n32093_ = new_n3823_ & ~new_n32092_;
  assign new_n32094_ = ~new_n32086_ & new_n32093_;
  assign new_n32095_ = ~new_n32088_ & ~new_n32094_;
  assign new_n32096_ = ~new_n31812_ & ~new_n32087_;
  assign new_n32097_ = ~new_n31814_ & new_n32084_;
  assign new_n32098_ = ~new_n32080_ & new_n32097_;
  assign new_n32099_ = ~new_n32081_ & ~new_n32084_;
  assign new_n32100_ = ~new_n32098_ & ~new_n32099_;
  assign new_n32101_ = new_n32087_ & ~new_n32100_;
  assign new_n32102_ = ~new_n32096_ & ~new_n32101_;
  assign new_n32103_ = ~\b[22]  & ~new_n32102_;
  assign new_n32104_ = ~\b[21]  & ~new_n32095_;
  assign new_n32105_ = ~new_n31822_ & ~new_n32087_;
  assign new_n32106_ = ~new_n31832_ & new_n32074_;
  assign new_n32107_ = ~new_n32070_ & new_n32106_;
  assign new_n32108_ = ~new_n32071_ & ~new_n32074_;
  assign new_n32109_ = ~new_n32107_ & ~new_n32108_;
  assign new_n32110_ = new_n3823_ & ~new_n32109_;
  assign new_n32111_ = ~new_n32086_ & new_n32110_;
  assign new_n32112_ = ~new_n32105_ & ~new_n32111_;
  assign new_n32113_ = ~\b[20]  & ~new_n32112_;
  assign new_n32114_ = ~new_n31831_ & ~new_n32087_;
  assign new_n32115_ = ~new_n31841_ & new_n32069_;
  assign new_n32116_ = ~new_n32065_ & new_n32115_;
  assign new_n32117_ = ~new_n32066_ & ~new_n32069_;
  assign new_n32118_ = ~new_n32116_ & ~new_n32117_;
  assign new_n32119_ = new_n3823_ & ~new_n32118_;
  assign new_n32120_ = ~new_n32086_ & new_n32119_;
  assign new_n32121_ = ~new_n32114_ & ~new_n32120_;
  assign new_n32122_ = ~\b[19]  & ~new_n32121_;
  assign new_n32123_ = ~new_n31840_ & ~new_n32087_;
  assign new_n32124_ = ~new_n31850_ & new_n32064_;
  assign new_n32125_ = ~new_n32060_ & new_n32124_;
  assign new_n32126_ = ~new_n32061_ & ~new_n32064_;
  assign new_n32127_ = ~new_n32125_ & ~new_n32126_;
  assign new_n32128_ = new_n3823_ & ~new_n32127_;
  assign new_n32129_ = ~new_n32086_ & new_n32128_;
  assign new_n32130_ = ~new_n32123_ & ~new_n32129_;
  assign new_n32131_ = ~\b[18]  & ~new_n32130_;
  assign new_n32132_ = ~new_n31849_ & ~new_n32087_;
  assign new_n32133_ = ~new_n31859_ & new_n32059_;
  assign new_n32134_ = ~new_n32055_ & new_n32133_;
  assign new_n32135_ = ~new_n32056_ & ~new_n32059_;
  assign new_n32136_ = ~new_n32134_ & ~new_n32135_;
  assign new_n32137_ = new_n3823_ & ~new_n32136_;
  assign new_n32138_ = ~new_n32086_ & new_n32137_;
  assign new_n32139_ = ~new_n32132_ & ~new_n32138_;
  assign new_n32140_ = ~\b[17]  & ~new_n32139_;
  assign new_n32141_ = ~new_n31858_ & ~new_n32087_;
  assign new_n32142_ = ~new_n31868_ & new_n32054_;
  assign new_n32143_ = ~new_n32050_ & new_n32142_;
  assign new_n32144_ = ~new_n32051_ & ~new_n32054_;
  assign new_n32145_ = ~new_n32143_ & ~new_n32144_;
  assign new_n32146_ = new_n3823_ & ~new_n32145_;
  assign new_n32147_ = ~new_n32086_ & new_n32146_;
  assign new_n32148_ = ~new_n32141_ & ~new_n32147_;
  assign new_n32149_ = ~\b[16]  & ~new_n32148_;
  assign new_n32150_ = ~new_n31867_ & ~new_n32087_;
  assign new_n32151_ = ~new_n31877_ & new_n32049_;
  assign new_n32152_ = ~new_n32045_ & new_n32151_;
  assign new_n32153_ = ~new_n32046_ & ~new_n32049_;
  assign new_n32154_ = ~new_n32152_ & ~new_n32153_;
  assign new_n32155_ = new_n3823_ & ~new_n32154_;
  assign new_n32156_ = ~new_n32086_ & new_n32155_;
  assign new_n32157_ = ~new_n32150_ & ~new_n32156_;
  assign new_n32158_ = ~\b[15]  & ~new_n32157_;
  assign new_n32159_ = ~new_n31876_ & ~new_n32087_;
  assign new_n32160_ = ~new_n31886_ & new_n32044_;
  assign new_n32161_ = ~new_n32040_ & new_n32160_;
  assign new_n32162_ = ~new_n32041_ & ~new_n32044_;
  assign new_n32163_ = ~new_n32161_ & ~new_n32162_;
  assign new_n32164_ = new_n3823_ & ~new_n32163_;
  assign new_n32165_ = ~new_n32086_ & new_n32164_;
  assign new_n32166_ = ~new_n32159_ & ~new_n32165_;
  assign new_n32167_ = ~\b[14]  & ~new_n32166_;
  assign new_n32168_ = ~new_n31885_ & ~new_n32087_;
  assign new_n32169_ = ~new_n31895_ & new_n32039_;
  assign new_n32170_ = ~new_n32035_ & new_n32169_;
  assign new_n32171_ = ~new_n32036_ & ~new_n32039_;
  assign new_n32172_ = ~new_n32170_ & ~new_n32171_;
  assign new_n32173_ = new_n3823_ & ~new_n32172_;
  assign new_n32174_ = ~new_n32086_ & new_n32173_;
  assign new_n32175_ = ~new_n32168_ & ~new_n32174_;
  assign new_n32176_ = ~\b[13]  & ~new_n32175_;
  assign new_n32177_ = ~new_n31894_ & ~new_n32087_;
  assign new_n32178_ = ~new_n31904_ & new_n32034_;
  assign new_n32179_ = ~new_n32030_ & new_n32178_;
  assign new_n32180_ = ~new_n32031_ & ~new_n32034_;
  assign new_n32181_ = ~new_n32179_ & ~new_n32180_;
  assign new_n32182_ = new_n3823_ & ~new_n32181_;
  assign new_n32183_ = ~new_n32086_ & new_n32182_;
  assign new_n32184_ = ~new_n32177_ & ~new_n32183_;
  assign new_n32185_ = ~\b[12]  & ~new_n32184_;
  assign new_n32186_ = ~new_n31903_ & ~new_n32087_;
  assign new_n32187_ = ~new_n31913_ & new_n32029_;
  assign new_n32188_ = ~new_n32025_ & new_n32187_;
  assign new_n32189_ = ~new_n32026_ & ~new_n32029_;
  assign new_n32190_ = ~new_n32188_ & ~new_n32189_;
  assign new_n32191_ = new_n3823_ & ~new_n32190_;
  assign new_n32192_ = ~new_n32086_ & new_n32191_;
  assign new_n32193_ = ~new_n32186_ & ~new_n32192_;
  assign new_n32194_ = ~\b[11]  & ~new_n32193_;
  assign new_n32195_ = ~new_n31912_ & ~new_n32087_;
  assign new_n32196_ = ~new_n31922_ & new_n32024_;
  assign new_n32197_ = ~new_n32020_ & new_n32196_;
  assign new_n32198_ = ~new_n32021_ & ~new_n32024_;
  assign new_n32199_ = ~new_n32197_ & ~new_n32198_;
  assign new_n32200_ = new_n3823_ & ~new_n32199_;
  assign new_n32201_ = ~new_n32086_ & new_n32200_;
  assign new_n32202_ = ~new_n32195_ & ~new_n32201_;
  assign new_n32203_ = ~\b[10]  & ~new_n32202_;
  assign new_n32204_ = ~new_n31921_ & ~new_n32087_;
  assign new_n32205_ = ~new_n31931_ & new_n32019_;
  assign new_n32206_ = ~new_n32015_ & new_n32205_;
  assign new_n32207_ = ~new_n32016_ & ~new_n32019_;
  assign new_n32208_ = ~new_n32206_ & ~new_n32207_;
  assign new_n32209_ = new_n3823_ & ~new_n32208_;
  assign new_n32210_ = ~new_n32086_ & new_n32209_;
  assign new_n32211_ = ~new_n32204_ & ~new_n32210_;
  assign new_n32212_ = ~\b[9]  & ~new_n32211_;
  assign new_n32213_ = ~new_n31930_ & ~new_n32087_;
  assign new_n32214_ = ~new_n31940_ & new_n32014_;
  assign new_n32215_ = ~new_n32010_ & new_n32214_;
  assign new_n32216_ = ~new_n32011_ & ~new_n32014_;
  assign new_n32217_ = ~new_n32215_ & ~new_n32216_;
  assign new_n32218_ = new_n3823_ & ~new_n32217_;
  assign new_n32219_ = ~new_n32086_ & new_n32218_;
  assign new_n32220_ = ~new_n32213_ & ~new_n32219_;
  assign new_n32221_ = ~\b[8]  & ~new_n32220_;
  assign new_n32222_ = ~new_n31939_ & ~new_n32087_;
  assign new_n32223_ = ~new_n31949_ & new_n32009_;
  assign new_n32224_ = ~new_n32005_ & new_n32223_;
  assign new_n32225_ = ~new_n32006_ & ~new_n32009_;
  assign new_n32226_ = ~new_n32224_ & ~new_n32225_;
  assign new_n32227_ = new_n3823_ & ~new_n32226_;
  assign new_n32228_ = ~new_n32086_ & new_n32227_;
  assign new_n32229_ = ~new_n32222_ & ~new_n32228_;
  assign new_n32230_ = ~\b[7]  & ~new_n32229_;
  assign new_n32231_ = ~new_n31948_ & ~new_n32087_;
  assign new_n32232_ = ~new_n31958_ & new_n32004_;
  assign new_n32233_ = ~new_n32000_ & new_n32232_;
  assign new_n32234_ = ~new_n32001_ & ~new_n32004_;
  assign new_n32235_ = ~new_n32233_ & ~new_n32234_;
  assign new_n32236_ = new_n3823_ & ~new_n32235_;
  assign new_n32237_ = ~new_n32086_ & new_n32236_;
  assign new_n32238_ = ~new_n32231_ & ~new_n32237_;
  assign new_n32239_ = ~\b[6]  & ~new_n32238_;
  assign new_n32240_ = ~new_n31957_ & ~new_n32087_;
  assign new_n32241_ = ~new_n31967_ & new_n31999_;
  assign new_n32242_ = ~new_n31995_ & new_n32241_;
  assign new_n32243_ = ~new_n31996_ & ~new_n31999_;
  assign new_n32244_ = ~new_n32242_ & ~new_n32243_;
  assign new_n32245_ = new_n3823_ & ~new_n32244_;
  assign new_n32246_ = ~new_n32086_ & new_n32245_;
  assign new_n32247_ = ~new_n32240_ & ~new_n32246_;
  assign new_n32248_ = ~\b[5]  & ~new_n32247_;
  assign new_n32249_ = ~new_n31966_ & ~new_n32087_;
  assign new_n32250_ = ~new_n31975_ & new_n31994_;
  assign new_n32251_ = ~new_n31990_ & new_n32250_;
  assign new_n32252_ = ~new_n31991_ & ~new_n31994_;
  assign new_n32253_ = ~new_n32251_ & ~new_n32252_;
  assign new_n32254_ = new_n3823_ & ~new_n32253_;
  assign new_n32255_ = ~new_n32086_ & new_n32254_;
  assign new_n32256_ = ~new_n32249_ & ~new_n32255_;
  assign new_n32257_ = ~\b[4]  & ~new_n32256_;
  assign new_n32258_ = ~new_n31974_ & ~new_n32087_;
  assign new_n32259_ = ~new_n31985_ & new_n31989_;
  assign new_n32260_ = ~new_n31984_ & new_n32259_;
  assign new_n32261_ = ~new_n31986_ & ~new_n31989_;
  assign new_n32262_ = ~new_n32260_ & ~new_n32261_;
  assign new_n32263_ = new_n3823_ & ~new_n32262_;
  assign new_n32264_ = ~new_n32086_ & new_n32263_;
  assign new_n32265_ = ~new_n32258_ & ~new_n32264_;
  assign new_n32266_ = ~\b[3]  & ~new_n32265_;
  assign new_n32267_ = ~new_n31979_ & ~new_n32087_;
  assign new_n32268_ = new_n3716_ & ~new_n31982_;
  assign new_n32269_ = ~new_n31980_ & new_n32268_;
  assign new_n32270_ = new_n3823_ & ~new_n32269_;
  assign new_n32271_ = ~new_n31984_ & new_n32270_;
  assign new_n32272_ = ~new_n32086_ & new_n32271_;
  assign new_n32273_ = ~new_n32267_ & ~new_n32272_;
  assign new_n32274_ = ~\b[2]  & ~new_n32273_;
  assign new_n32275_ = new_n4017_ & ~new_n32086_;
  assign new_n32276_ = \a[42]  & ~new_n32275_;
  assign new_n32277_ = new_n4024_ & ~new_n32086_;
  assign new_n32278_ = ~new_n32276_ & ~new_n32277_;
  assign new_n32279_ = \b[1]  & ~new_n32278_;
  assign new_n32280_ = ~\b[1]  & ~new_n32277_;
  assign new_n32281_ = ~new_n32276_ & new_n32280_;
  assign new_n32282_ = ~new_n32279_ & ~new_n32281_;
  assign new_n32283_ = ~new_n4031_ & ~new_n32282_;
  assign new_n32284_ = ~\b[1]  & ~new_n32278_;
  assign new_n32285_ = ~new_n32283_ & ~new_n32284_;
  assign new_n32286_ = \b[2]  & ~new_n32272_;
  assign new_n32287_ = ~new_n32267_ & new_n32286_;
  assign new_n32288_ = ~new_n32274_ & ~new_n32287_;
  assign new_n32289_ = ~new_n32285_ & new_n32288_;
  assign new_n32290_ = ~new_n32274_ & ~new_n32289_;
  assign new_n32291_ = \b[3]  & ~new_n32264_;
  assign new_n32292_ = ~new_n32258_ & new_n32291_;
  assign new_n32293_ = ~new_n32266_ & ~new_n32292_;
  assign new_n32294_ = ~new_n32290_ & new_n32293_;
  assign new_n32295_ = ~new_n32266_ & ~new_n32294_;
  assign new_n32296_ = \b[4]  & ~new_n32255_;
  assign new_n32297_ = ~new_n32249_ & new_n32296_;
  assign new_n32298_ = ~new_n32257_ & ~new_n32297_;
  assign new_n32299_ = ~new_n32295_ & new_n32298_;
  assign new_n32300_ = ~new_n32257_ & ~new_n32299_;
  assign new_n32301_ = \b[5]  & ~new_n32246_;
  assign new_n32302_ = ~new_n32240_ & new_n32301_;
  assign new_n32303_ = ~new_n32248_ & ~new_n32302_;
  assign new_n32304_ = ~new_n32300_ & new_n32303_;
  assign new_n32305_ = ~new_n32248_ & ~new_n32304_;
  assign new_n32306_ = \b[6]  & ~new_n32237_;
  assign new_n32307_ = ~new_n32231_ & new_n32306_;
  assign new_n32308_ = ~new_n32239_ & ~new_n32307_;
  assign new_n32309_ = ~new_n32305_ & new_n32308_;
  assign new_n32310_ = ~new_n32239_ & ~new_n32309_;
  assign new_n32311_ = \b[7]  & ~new_n32228_;
  assign new_n32312_ = ~new_n32222_ & new_n32311_;
  assign new_n32313_ = ~new_n32230_ & ~new_n32312_;
  assign new_n32314_ = ~new_n32310_ & new_n32313_;
  assign new_n32315_ = ~new_n32230_ & ~new_n32314_;
  assign new_n32316_ = \b[8]  & ~new_n32219_;
  assign new_n32317_ = ~new_n32213_ & new_n32316_;
  assign new_n32318_ = ~new_n32221_ & ~new_n32317_;
  assign new_n32319_ = ~new_n32315_ & new_n32318_;
  assign new_n32320_ = ~new_n32221_ & ~new_n32319_;
  assign new_n32321_ = \b[9]  & ~new_n32210_;
  assign new_n32322_ = ~new_n32204_ & new_n32321_;
  assign new_n32323_ = ~new_n32212_ & ~new_n32322_;
  assign new_n32324_ = ~new_n32320_ & new_n32323_;
  assign new_n32325_ = ~new_n32212_ & ~new_n32324_;
  assign new_n32326_ = \b[10]  & ~new_n32201_;
  assign new_n32327_ = ~new_n32195_ & new_n32326_;
  assign new_n32328_ = ~new_n32203_ & ~new_n32327_;
  assign new_n32329_ = ~new_n32325_ & new_n32328_;
  assign new_n32330_ = ~new_n32203_ & ~new_n32329_;
  assign new_n32331_ = \b[11]  & ~new_n32192_;
  assign new_n32332_ = ~new_n32186_ & new_n32331_;
  assign new_n32333_ = ~new_n32194_ & ~new_n32332_;
  assign new_n32334_ = ~new_n32330_ & new_n32333_;
  assign new_n32335_ = ~new_n32194_ & ~new_n32334_;
  assign new_n32336_ = \b[12]  & ~new_n32183_;
  assign new_n32337_ = ~new_n32177_ & new_n32336_;
  assign new_n32338_ = ~new_n32185_ & ~new_n32337_;
  assign new_n32339_ = ~new_n32335_ & new_n32338_;
  assign new_n32340_ = ~new_n32185_ & ~new_n32339_;
  assign new_n32341_ = \b[13]  & ~new_n32174_;
  assign new_n32342_ = ~new_n32168_ & new_n32341_;
  assign new_n32343_ = ~new_n32176_ & ~new_n32342_;
  assign new_n32344_ = ~new_n32340_ & new_n32343_;
  assign new_n32345_ = ~new_n32176_ & ~new_n32344_;
  assign new_n32346_ = \b[14]  & ~new_n32165_;
  assign new_n32347_ = ~new_n32159_ & new_n32346_;
  assign new_n32348_ = ~new_n32167_ & ~new_n32347_;
  assign new_n32349_ = ~new_n32345_ & new_n32348_;
  assign new_n32350_ = ~new_n32167_ & ~new_n32349_;
  assign new_n32351_ = \b[15]  & ~new_n32156_;
  assign new_n32352_ = ~new_n32150_ & new_n32351_;
  assign new_n32353_ = ~new_n32158_ & ~new_n32352_;
  assign new_n32354_ = ~new_n32350_ & new_n32353_;
  assign new_n32355_ = ~new_n32158_ & ~new_n32354_;
  assign new_n32356_ = \b[16]  & ~new_n32147_;
  assign new_n32357_ = ~new_n32141_ & new_n32356_;
  assign new_n32358_ = ~new_n32149_ & ~new_n32357_;
  assign new_n32359_ = ~new_n32355_ & new_n32358_;
  assign new_n32360_ = ~new_n32149_ & ~new_n32359_;
  assign new_n32361_ = \b[17]  & ~new_n32138_;
  assign new_n32362_ = ~new_n32132_ & new_n32361_;
  assign new_n32363_ = ~new_n32140_ & ~new_n32362_;
  assign new_n32364_ = ~new_n32360_ & new_n32363_;
  assign new_n32365_ = ~new_n32140_ & ~new_n32364_;
  assign new_n32366_ = \b[18]  & ~new_n32129_;
  assign new_n32367_ = ~new_n32123_ & new_n32366_;
  assign new_n32368_ = ~new_n32131_ & ~new_n32367_;
  assign new_n32369_ = ~new_n32365_ & new_n32368_;
  assign new_n32370_ = ~new_n32131_ & ~new_n32369_;
  assign new_n32371_ = \b[19]  & ~new_n32120_;
  assign new_n32372_ = ~new_n32114_ & new_n32371_;
  assign new_n32373_ = ~new_n32122_ & ~new_n32372_;
  assign new_n32374_ = ~new_n32370_ & new_n32373_;
  assign new_n32375_ = ~new_n32122_ & ~new_n32374_;
  assign new_n32376_ = \b[20]  & ~new_n32111_;
  assign new_n32377_ = ~new_n32105_ & new_n32376_;
  assign new_n32378_ = ~new_n32113_ & ~new_n32377_;
  assign new_n32379_ = ~new_n32375_ & new_n32378_;
  assign new_n32380_ = ~new_n32113_ & ~new_n32379_;
  assign new_n32381_ = \b[21]  & ~new_n32094_;
  assign new_n32382_ = ~new_n32088_ & new_n32381_;
  assign new_n32383_ = ~new_n32104_ & ~new_n32382_;
  assign new_n32384_ = ~new_n32380_ & new_n32383_;
  assign new_n32385_ = ~new_n32104_ & ~new_n32384_;
  assign new_n32386_ = \b[22]  & ~new_n32096_;
  assign new_n32387_ = ~new_n32101_ & new_n32386_;
  assign new_n32388_ = ~new_n32103_ & ~new_n32387_;
  assign new_n32389_ = ~new_n32385_ & new_n32388_;
  assign new_n32390_ = ~new_n32103_ & ~new_n32389_;
  assign new_n32391_ = new_n4143_ & ~new_n32390_;
  assign new_n32392_ = ~new_n32095_ & ~new_n32391_;
  assign new_n32393_ = ~new_n32113_ & new_n32383_;
  assign new_n32394_ = ~new_n32379_ & new_n32393_;
  assign new_n32395_ = ~new_n32380_ & ~new_n32383_;
  assign new_n32396_ = ~new_n32394_ & ~new_n32395_;
  assign new_n32397_ = new_n4143_ & ~new_n32396_;
  assign new_n32398_ = ~new_n32390_ & new_n32397_;
  assign new_n32399_ = ~new_n32392_ & ~new_n32398_;
  assign new_n32400_ = ~\b[22]  & ~new_n32399_;
  assign new_n32401_ = ~new_n32112_ & ~new_n32391_;
  assign new_n32402_ = ~new_n32122_ & new_n32378_;
  assign new_n32403_ = ~new_n32374_ & new_n32402_;
  assign new_n32404_ = ~new_n32375_ & ~new_n32378_;
  assign new_n32405_ = ~new_n32403_ & ~new_n32404_;
  assign new_n32406_ = new_n4143_ & ~new_n32405_;
  assign new_n32407_ = ~new_n32390_ & new_n32406_;
  assign new_n32408_ = ~new_n32401_ & ~new_n32407_;
  assign new_n32409_ = ~\b[21]  & ~new_n32408_;
  assign new_n32410_ = ~new_n32121_ & ~new_n32391_;
  assign new_n32411_ = ~new_n32131_ & new_n32373_;
  assign new_n32412_ = ~new_n32369_ & new_n32411_;
  assign new_n32413_ = ~new_n32370_ & ~new_n32373_;
  assign new_n32414_ = ~new_n32412_ & ~new_n32413_;
  assign new_n32415_ = new_n4143_ & ~new_n32414_;
  assign new_n32416_ = ~new_n32390_ & new_n32415_;
  assign new_n32417_ = ~new_n32410_ & ~new_n32416_;
  assign new_n32418_ = ~\b[20]  & ~new_n32417_;
  assign new_n32419_ = ~new_n32130_ & ~new_n32391_;
  assign new_n32420_ = ~new_n32140_ & new_n32368_;
  assign new_n32421_ = ~new_n32364_ & new_n32420_;
  assign new_n32422_ = ~new_n32365_ & ~new_n32368_;
  assign new_n32423_ = ~new_n32421_ & ~new_n32422_;
  assign new_n32424_ = new_n4143_ & ~new_n32423_;
  assign new_n32425_ = ~new_n32390_ & new_n32424_;
  assign new_n32426_ = ~new_n32419_ & ~new_n32425_;
  assign new_n32427_ = ~\b[19]  & ~new_n32426_;
  assign new_n32428_ = ~new_n32139_ & ~new_n32391_;
  assign new_n32429_ = ~new_n32149_ & new_n32363_;
  assign new_n32430_ = ~new_n32359_ & new_n32429_;
  assign new_n32431_ = ~new_n32360_ & ~new_n32363_;
  assign new_n32432_ = ~new_n32430_ & ~new_n32431_;
  assign new_n32433_ = new_n4143_ & ~new_n32432_;
  assign new_n32434_ = ~new_n32390_ & new_n32433_;
  assign new_n32435_ = ~new_n32428_ & ~new_n32434_;
  assign new_n32436_ = ~\b[18]  & ~new_n32435_;
  assign new_n32437_ = ~new_n32148_ & ~new_n32391_;
  assign new_n32438_ = ~new_n32158_ & new_n32358_;
  assign new_n32439_ = ~new_n32354_ & new_n32438_;
  assign new_n32440_ = ~new_n32355_ & ~new_n32358_;
  assign new_n32441_ = ~new_n32439_ & ~new_n32440_;
  assign new_n32442_ = new_n4143_ & ~new_n32441_;
  assign new_n32443_ = ~new_n32390_ & new_n32442_;
  assign new_n32444_ = ~new_n32437_ & ~new_n32443_;
  assign new_n32445_ = ~\b[17]  & ~new_n32444_;
  assign new_n32446_ = ~new_n32157_ & ~new_n32391_;
  assign new_n32447_ = ~new_n32167_ & new_n32353_;
  assign new_n32448_ = ~new_n32349_ & new_n32447_;
  assign new_n32449_ = ~new_n32350_ & ~new_n32353_;
  assign new_n32450_ = ~new_n32448_ & ~new_n32449_;
  assign new_n32451_ = new_n4143_ & ~new_n32450_;
  assign new_n32452_ = ~new_n32390_ & new_n32451_;
  assign new_n32453_ = ~new_n32446_ & ~new_n32452_;
  assign new_n32454_ = ~\b[16]  & ~new_n32453_;
  assign new_n32455_ = ~new_n32166_ & ~new_n32391_;
  assign new_n32456_ = ~new_n32176_ & new_n32348_;
  assign new_n32457_ = ~new_n32344_ & new_n32456_;
  assign new_n32458_ = ~new_n32345_ & ~new_n32348_;
  assign new_n32459_ = ~new_n32457_ & ~new_n32458_;
  assign new_n32460_ = new_n4143_ & ~new_n32459_;
  assign new_n32461_ = ~new_n32390_ & new_n32460_;
  assign new_n32462_ = ~new_n32455_ & ~new_n32461_;
  assign new_n32463_ = ~\b[15]  & ~new_n32462_;
  assign new_n32464_ = ~new_n32175_ & ~new_n32391_;
  assign new_n32465_ = ~new_n32185_ & new_n32343_;
  assign new_n32466_ = ~new_n32339_ & new_n32465_;
  assign new_n32467_ = ~new_n32340_ & ~new_n32343_;
  assign new_n32468_ = ~new_n32466_ & ~new_n32467_;
  assign new_n32469_ = new_n4143_ & ~new_n32468_;
  assign new_n32470_ = ~new_n32390_ & new_n32469_;
  assign new_n32471_ = ~new_n32464_ & ~new_n32470_;
  assign new_n32472_ = ~\b[14]  & ~new_n32471_;
  assign new_n32473_ = ~new_n32184_ & ~new_n32391_;
  assign new_n32474_ = ~new_n32194_ & new_n32338_;
  assign new_n32475_ = ~new_n32334_ & new_n32474_;
  assign new_n32476_ = ~new_n32335_ & ~new_n32338_;
  assign new_n32477_ = ~new_n32475_ & ~new_n32476_;
  assign new_n32478_ = new_n4143_ & ~new_n32477_;
  assign new_n32479_ = ~new_n32390_ & new_n32478_;
  assign new_n32480_ = ~new_n32473_ & ~new_n32479_;
  assign new_n32481_ = ~\b[13]  & ~new_n32480_;
  assign new_n32482_ = ~new_n32193_ & ~new_n32391_;
  assign new_n32483_ = ~new_n32203_ & new_n32333_;
  assign new_n32484_ = ~new_n32329_ & new_n32483_;
  assign new_n32485_ = ~new_n32330_ & ~new_n32333_;
  assign new_n32486_ = ~new_n32484_ & ~new_n32485_;
  assign new_n32487_ = new_n4143_ & ~new_n32486_;
  assign new_n32488_ = ~new_n32390_ & new_n32487_;
  assign new_n32489_ = ~new_n32482_ & ~new_n32488_;
  assign new_n32490_ = ~\b[12]  & ~new_n32489_;
  assign new_n32491_ = ~new_n32202_ & ~new_n32391_;
  assign new_n32492_ = ~new_n32212_ & new_n32328_;
  assign new_n32493_ = ~new_n32324_ & new_n32492_;
  assign new_n32494_ = ~new_n32325_ & ~new_n32328_;
  assign new_n32495_ = ~new_n32493_ & ~new_n32494_;
  assign new_n32496_ = new_n4143_ & ~new_n32495_;
  assign new_n32497_ = ~new_n32390_ & new_n32496_;
  assign new_n32498_ = ~new_n32491_ & ~new_n32497_;
  assign new_n32499_ = ~\b[11]  & ~new_n32498_;
  assign new_n32500_ = ~new_n32211_ & ~new_n32391_;
  assign new_n32501_ = ~new_n32221_ & new_n32323_;
  assign new_n32502_ = ~new_n32319_ & new_n32501_;
  assign new_n32503_ = ~new_n32320_ & ~new_n32323_;
  assign new_n32504_ = ~new_n32502_ & ~new_n32503_;
  assign new_n32505_ = new_n4143_ & ~new_n32504_;
  assign new_n32506_ = ~new_n32390_ & new_n32505_;
  assign new_n32507_ = ~new_n32500_ & ~new_n32506_;
  assign new_n32508_ = ~\b[10]  & ~new_n32507_;
  assign new_n32509_ = ~new_n32220_ & ~new_n32391_;
  assign new_n32510_ = ~new_n32230_ & new_n32318_;
  assign new_n32511_ = ~new_n32314_ & new_n32510_;
  assign new_n32512_ = ~new_n32315_ & ~new_n32318_;
  assign new_n32513_ = ~new_n32511_ & ~new_n32512_;
  assign new_n32514_ = new_n4143_ & ~new_n32513_;
  assign new_n32515_ = ~new_n32390_ & new_n32514_;
  assign new_n32516_ = ~new_n32509_ & ~new_n32515_;
  assign new_n32517_ = ~\b[9]  & ~new_n32516_;
  assign new_n32518_ = ~new_n32229_ & ~new_n32391_;
  assign new_n32519_ = ~new_n32239_ & new_n32313_;
  assign new_n32520_ = ~new_n32309_ & new_n32519_;
  assign new_n32521_ = ~new_n32310_ & ~new_n32313_;
  assign new_n32522_ = ~new_n32520_ & ~new_n32521_;
  assign new_n32523_ = new_n4143_ & ~new_n32522_;
  assign new_n32524_ = ~new_n32390_ & new_n32523_;
  assign new_n32525_ = ~new_n32518_ & ~new_n32524_;
  assign new_n32526_ = ~\b[8]  & ~new_n32525_;
  assign new_n32527_ = ~new_n32238_ & ~new_n32391_;
  assign new_n32528_ = ~new_n32248_ & new_n32308_;
  assign new_n32529_ = ~new_n32304_ & new_n32528_;
  assign new_n32530_ = ~new_n32305_ & ~new_n32308_;
  assign new_n32531_ = ~new_n32529_ & ~new_n32530_;
  assign new_n32532_ = new_n4143_ & ~new_n32531_;
  assign new_n32533_ = ~new_n32390_ & new_n32532_;
  assign new_n32534_ = ~new_n32527_ & ~new_n32533_;
  assign new_n32535_ = ~\b[7]  & ~new_n32534_;
  assign new_n32536_ = ~new_n32247_ & ~new_n32391_;
  assign new_n32537_ = ~new_n32257_ & new_n32303_;
  assign new_n32538_ = ~new_n32299_ & new_n32537_;
  assign new_n32539_ = ~new_n32300_ & ~new_n32303_;
  assign new_n32540_ = ~new_n32538_ & ~new_n32539_;
  assign new_n32541_ = new_n4143_ & ~new_n32540_;
  assign new_n32542_ = ~new_n32390_ & new_n32541_;
  assign new_n32543_ = ~new_n32536_ & ~new_n32542_;
  assign new_n32544_ = ~\b[6]  & ~new_n32543_;
  assign new_n32545_ = ~new_n32256_ & ~new_n32391_;
  assign new_n32546_ = ~new_n32266_ & new_n32298_;
  assign new_n32547_ = ~new_n32294_ & new_n32546_;
  assign new_n32548_ = ~new_n32295_ & ~new_n32298_;
  assign new_n32549_ = ~new_n32547_ & ~new_n32548_;
  assign new_n32550_ = new_n4143_ & ~new_n32549_;
  assign new_n32551_ = ~new_n32390_ & new_n32550_;
  assign new_n32552_ = ~new_n32545_ & ~new_n32551_;
  assign new_n32553_ = ~\b[5]  & ~new_n32552_;
  assign new_n32554_ = ~new_n32265_ & ~new_n32391_;
  assign new_n32555_ = ~new_n32274_ & new_n32293_;
  assign new_n32556_ = ~new_n32289_ & new_n32555_;
  assign new_n32557_ = ~new_n32290_ & ~new_n32293_;
  assign new_n32558_ = ~new_n32556_ & ~new_n32557_;
  assign new_n32559_ = new_n4143_ & ~new_n32558_;
  assign new_n32560_ = ~new_n32390_ & new_n32559_;
  assign new_n32561_ = ~new_n32554_ & ~new_n32560_;
  assign new_n32562_ = ~\b[4]  & ~new_n32561_;
  assign new_n32563_ = ~new_n32273_ & ~new_n32391_;
  assign new_n32564_ = ~new_n32284_ & new_n32288_;
  assign new_n32565_ = ~new_n32283_ & new_n32564_;
  assign new_n32566_ = ~new_n32285_ & ~new_n32288_;
  assign new_n32567_ = ~new_n32565_ & ~new_n32566_;
  assign new_n32568_ = new_n4143_ & ~new_n32567_;
  assign new_n32569_ = ~new_n32390_ & new_n32568_;
  assign new_n32570_ = ~new_n32563_ & ~new_n32569_;
  assign new_n32571_ = ~\b[3]  & ~new_n32570_;
  assign new_n32572_ = ~new_n32278_ & ~new_n32391_;
  assign new_n32573_ = new_n4031_ & ~new_n32281_;
  assign new_n32574_ = ~new_n32279_ & new_n32573_;
  assign new_n32575_ = new_n4143_ & ~new_n32574_;
  assign new_n32576_ = ~new_n32283_ & new_n32575_;
  assign new_n32577_ = ~new_n32390_ & new_n32576_;
  assign new_n32578_ = ~new_n32572_ & ~new_n32577_;
  assign new_n32579_ = ~\b[2]  & ~new_n32578_;
  assign new_n32580_ = new_n4337_ & ~new_n32390_;
  assign new_n32581_ = \a[41]  & ~new_n32580_;
  assign new_n32582_ = new_n4344_ & ~new_n32390_;
  assign new_n32583_ = ~new_n32581_ & ~new_n32582_;
  assign new_n32584_ = \b[1]  & ~new_n32583_;
  assign new_n32585_ = ~\b[1]  & ~new_n32582_;
  assign new_n32586_ = ~new_n32581_ & new_n32585_;
  assign new_n32587_ = ~new_n32584_ & ~new_n32586_;
  assign new_n32588_ = ~new_n4351_ & ~new_n32587_;
  assign new_n32589_ = ~\b[1]  & ~new_n32583_;
  assign new_n32590_ = ~new_n32588_ & ~new_n32589_;
  assign new_n32591_ = \b[2]  & ~new_n32577_;
  assign new_n32592_ = ~new_n32572_ & new_n32591_;
  assign new_n32593_ = ~new_n32579_ & ~new_n32592_;
  assign new_n32594_ = ~new_n32590_ & new_n32593_;
  assign new_n32595_ = ~new_n32579_ & ~new_n32594_;
  assign new_n32596_ = \b[3]  & ~new_n32569_;
  assign new_n32597_ = ~new_n32563_ & new_n32596_;
  assign new_n32598_ = ~new_n32571_ & ~new_n32597_;
  assign new_n32599_ = ~new_n32595_ & new_n32598_;
  assign new_n32600_ = ~new_n32571_ & ~new_n32599_;
  assign new_n32601_ = \b[4]  & ~new_n32560_;
  assign new_n32602_ = ~new_n32554_ & new_n32601_;
  assign new_n32603_ = ~new_n32562_ & ~new_n32602_;
  assign new_n32604_ = ~new_n32600_ & new_n32603_;
  assign new_n32605_ = ~new_n32562_ & ~new_n32604_;
  assign new_n32606_ = \b[5]  & ~new_n32551_;
  assign new_n32607_ = ~new_n32545_ & new_n32606_;
  assign new_n32608_ = ~new_n32553_ & ~new_n32607_;
  assign new_n32609_ = ~new_n32605_ & new_n32608_;
  assign new_n32610_ = ~new_n32553_ & ~new_n32609_;
  assign new_n32611_ = \b[6]  & ~new_n32542_;
  assign new_n32612_ = ~new_n32536_ & new_n32611_;
  assign new_n32613_ = ~new_n32544_ & ~new_n32612_;
  assign new_n32614_ = ~new_n32610_ & new_n32613_;
  assign new_n32615_ = ~new_n32544_ & ~new_n32614_;
  assign new_n32616_ = \b[7]  & ~new_n32533_;
  assign new_n32617_ = ~new_n32527_ & new_n32616_;
  assign new_n32618_ = ~new_n32535_ & ~new_n32617_;
  assign new_n32619_ = ~new_n32615_ & new_n32618_;
  assign new_n32620_ = ~new_n32535_ & ~new_n32619_;
  assign new_n32621_ = \b[8]  & ~new_n32524_;
  assign new_n32622_ = ~new_n32518_ & new_n32621_;
  assign new_n32623_ = ~new_n32526_ & ~new_n32622_;
  assign new_n32624_ = ~new_n32620_ & new_n32623_;
  assign new_n32625_ = ~new_n32526_ & ~new_n32624_;
  assign new_n32626_ = \b[9]  & ~new_n32515_;
  assign new_n32627_ = ~new_n32509_ & new_n32626_;
  assign new_n32628_ = ~new_n32517_ & ~new_n32627_;
  assign new_n32629_ = ~new_n32625_ & new_n32628_;
  assign new_n32630_ = ~new_n32517_ & ~new_n32629_;
  assign new_n32631_ = \b[10]  & ~new_n32506_;
  assign new_n32632_ = ~new_n32500_ & new_n32631_;
  assign new_n32633_ = ~new_n32508_ & ~new_n32632_;
  assign new_n32634_ = ~new_n32630_ & new_n32633_;
  assign new_n32635_ = ~new_n32508_ & ~new_n32634_;
  assign new_n32636_ = \b[11]  & ~new_n32497_;
  assign new_n32637_ = ~new_n32491_ & new_n32636_;
  assign new_n32638_ = ~new_n32499_ & ~new_n32637_;
  assign new_n32639_ = ~new_n32635_ & new_n32638_;
  assign new_n32640_ = ~new_n32499_ & ~new_n32639_;
  assign new_n32641_ = \b[12]  & ~new_n32488_;
  assign new_n32642_ = ~new_n32482_ & new_n32641_;
  assign new_n32643_ = ~new_n32490_ & ~new_n32642_;
  assign new_n32644_ = ~new_n32640_ & new_n32643_;
  assign new_n32645_ = ~new_n32490_ & ~new_n32644_;
  assign new_n32646_ = \b[13]  & ~new_n32479_;
  assign new_n32647_ = ~new_n32473_ & new_n32646_;
  assign new_n32648_ = ~new_n32481_ & ~new_n32647_;
  assign new_n32649_ = ~new_n32645_ & new_n32648_;
  assign new_n32650_ = ~new_n32481_ & ~new_n32649_;
  assign new_n32651_ = \b[14]  & ~new_n32470_;
  assign new_n32652_ = ~new_n32464_ & new_n32651_;
  assign new_n32653_ = ~new_n32472_ & ~new_n32652_;
  assign new_n32654_ = ~new_n32650_ & new_n32653_;
  assign new_n32655_ = ~new_n32472_ & ~new_n32654_;
  assign new_n32656_ = \b[15]  & ~new_n32461_;
  assign new_n32657_ = ~new_n32455_ & new_n32656_;
  assign new_n32658_ = ~new_n32463_ & ~new_n32657_;
  assign new_n32659_ = ~new_n32655_ & new_n32658_;
  assign new_n32660_ = ~new_n32463_ & ~new_n32659_;
  assign new_n32661_ = \b[16]  & ~new_n32452_;
  assign new_n32662_ = ~new_n32446_ & new_n32661_;
  assign new_n32663_ = ~new_n32454_ & ~new_n32662_;
  assign new_n32664_ = ~new_n32660_ & new_n32663_;
  assign new_n32665_ = ~new_n32454_ & ~new_n32664_;
  assign new_n32666_ = \b[17]  & ~new_n32443_;
  assign new_n32667_ = ~new_n32437_ & new_n32666_;
  assign new_n32668_ = ~new_n32445_ & ~new_n32667_;
  assign new_n32669_ = ~new_n32665_ & new_n32668_;
  assign new_n32670_ = ~new_n32445_ & ~new_n32669_;
  assign new_n32671_ = \b[18]  & ~new_n32434_;
  assign new_n32672_ = ~new_n32428_ & new_n32671_;
  assign new_n32673_ = ~new_n32436_ & ~new_n32672_;
  assign new_n32674_ = ~new_n32670_ & new_n32673_;
  assign new_n32675_ = ~new_n32436_ & ~new_n32674_;
  assign new_n32676_ = \b[19]  & ~new_n32425_;
  assign new_n32677_ = ~new_n32419_ & new_n32676_;
  assign new_n32678_ = ~new_n32427_ & ~new_n32677_;
  assign new_n32679_ = ~new_n32675_ & new_n32678_;
  assign new_n32680_ = ~new_n32427_ & ~new_n32679_;
  assign new_n32681_ = \b[20]  & ~new_n32416_;
  assign new_n32682_ = ~new_n32410_ & new_n32681_;
  assign new_n32683_ = ~new_n32418_ & ~new_n32682_;
  assign new_n32684_ = ~new_n32680_ & new_n32683_;
  assign new_n32685_ = ~new_n32418_ & ~new_n32684_;
  assign new_n32686_ = \b[21]  & ~new_n32407_;
  assign new_n32687_ = ~new_n32401_ & new_n32686_;
  assign new_n32688_ = ~new_n32409_ & ~new_n32687_;
  assign new_n32689_ = ~new_n32685_ & new_n32688_;
  assign new_n32690_ = ~new_n32409_ & ~new_n32689_;
  assign new_n32691_ = \b[22]  & ~new_n32398_;
  assign new_n32692_ = ~new_n32392_ & new_n32691_;
  assign new_n32693_ = ~new_n32400_ & ~new_n32692_;
  assign new_n32694_ = ~new_n32690_ & new_n32693_;
  assign new_n32695_ = ~new_n32400_ & ~new_n32694_;
  assign new_n32696_ = ~new_n32102_ & ~new_n32391_;
  assign new_n32697_ = ~new_n32104_ & new_n32388_;
  assign new_n32698_ = ~new_n32384_ & new_n32697_;
  assign new_n32699_ = ~new_n32385_ & ~new_n32388_;
  assign new_n32700_ = ~new_n32698_ & ~new_n32699_;
  assign new_n32701_ = new_n32391_ & ~new_n32700_;
  assign new_n32702_ = ~new_n32696_ & ~new_n32701_;
  assign new_n32703_ = ~\b[23]  & ~new_n32702_;
  assign new_n32704_ = \b[23]  & ~new_n32696_;
  assign new_n32705_ = ~new_n32701_ & new_n32704_;
  assign new_n32706_ = new_n4471_ & ~new_n32705_;
  assign new_n32707_ = ~new_n32703_ & new_n32706_;
  assign new_n32708_ = ~new_n32695_ & new_n32707_;
  assign new_n32709_ = new_n4143_ & ~new_n32702_;
  assign new_n32710_ = ~new_n32708_ & ~new_n32709_;
  assign new_n32711_ = ~new_n32409_ & new_n32693_;
  assign new_n32712_ = ~new_n32689_ & new_n32711_;
  assign new_n32713_ = ~new_n32690_ & ~new_n32693_;
  assign new_n32714_ = ~new_n32712_ & ~new_n32713_;
  assign new_n32715_ = ~new_n32710_ & ~new_n32714_;
  assign new_n32716_ = ~new_n32399_ & ~new_n32709_;
  assign new_n32717_ = ~new_n32708_ & new_n32716_;
  assign new_n32718_ = ~new_n32715_ & ~new_n32717_;
  assign new_n32719_ = ~new_n32400_ & ~new_n32705_;
  assign new_n32720_ = ~new_n32703_ & new_n32719_;
  assign new_n32721_ = ~new_n32694_ & new_n32720_;
  assign new_n32722_ = ~new_n32703_ & ~new_n32705_;
  assign new_n32723_ = ~new_n32695_ & ~new_n32722_;
  assign new_n32724_ = ~new_n32721_ & ~new_n32723_;
  assign new_n32725_ = ~new_n32710_ & ~new_n32724_;
  assign new_n32726_ = ~new_n32702_ & ~new_n32709_;
  assign new_n32727_ = ~new_n32708_ & new_n32726_;
  assign new_n32728_ = ~new_n32725_ & ~new_n32727_;
  assign new_n32729_ = ~\b[24]  & ~new_n32728_;
  assign new_n32730_ = ~\b[23]  & ~new_n32718_;
  assign new_n32731_ = ~new_n32418_ & new_n32688_;
  assign new_n32732_ = ~new_n32684_ & new_n32731_;
  assign new_n32733_ = ~new_n32685_ & ~new_n32688_;
  assign new_n32734_ = ~new_n32732_ & ~new_n32733_;
  assign new_n32735_ = ~new_n32710_ & ~new_n32734_;
  assign new_n32736_ = ~new_n32408_ & ~new_n32709_;
  assign new_n32737_ = ~new_n32708_ & new_n32736_;
  assign new_n32738_ = ~new_n32735_ & ~new_n32737_;
  assign new_n32739_ = ~\b[22]  & ~new_n32738_;
  assign new_n32740_ = ~new_n32427_ & new_n32683_;
  assign new_n32741_ = ~new_n32679_ & new_n32740_;
  assign new_n32742_ = ~new_n32680_ & ~new_n32683_;
  assign new_n32743_ = ~new_n32741_ & ~new_n32742_;
  assign new_n32744_ = ~new_n32710_ & ~new_n32743_;
  assign new_n32745_ = ~new_n32417_ & ~new_n32709_;
  assign new_n32746_ = ~new_n32708_ & new_n32745_;
  assign new_n32747_ = ~new_n32744_ & ~new_n32746_;
  assign new_n32748_ = ~\b[21]  & ~new_n32747_;
  assign new_n32749_ = ~new_n32436_ & new_n32678_;
  assign new_n32750_ = ~new_n32674_ & new_n32749_;
  assign new_n32751_ = ~new_n32675_ & ~new_n32678_;
  assign new_n32752_ = ~new_n32750_ & ~new_n32751_;
  assign new_n32753_ = ~new_n32710_ & ~new_n32752_;
  assign new_n32754_ = ~new_n32426_ & ~new_n32709_;
  assign new_n32755_ = ~new_n32708_ & new_n32754_;
  assign new_n32756_ = ~new_n32753_ & ~new_n32755_;
  assign new_n32757_ = ~\b[20]  & ~new_n32756_;
  assign new_n32758_ = ~new_n32445_ & new_n32673_;
  assign new_n32759_ = ~new_n32669_ & new_n32758_;
  assign new_n32760_ = ~new_n32670_ & ~new_n32673_;
  assign new_n32761_ = ~new_n32759_ & ~new_n32760_;
  assign new_n32762_ = ~new_n32710_ & ~new_n32761_;
  assign new_n32763_ = ~new_n32435_ & ~new_n32709_;
  assign new_n32764_ = ~new_n32708_ & new_n32763_;
  assign new_n32765_ = ~new_n32762_ & ~new_n32764_;
  assign new_n32766_ = ~\b[19]  & ~new_n32765_;
  assign new_n32767_ = ~new_n32454_ & new_n32668_;
  assign new_n32768_ = ~new_n32664_ & new_n32767_;
  assign new_n32769_ = ~new_n32665_ & ~new_n32668_;
  assign new_n32770_ = ~new_n32768_ & ~new_n32769_;
  assign new_n32771_ = ~new_n32710_ & ~new_n32770_;
  assign new_n32772_ = ~new_n32444_ & ~new_n32709_;
  assign new_n32773_ = ~new_n32708_ & new_n32772_;
  assign new_n32774_ = ~new_n32771_ & ~new_n32773_;
  assign new_n32775_ = ~\b[18]  & ~new_n32774_;
  assign new_n32776_ = ~new_n32463_ & new_n32663_;
  assign new_n32777_ = ~new_n32659_ & new_n32776_;
  assign new_n32778_ = ~new_n32660_ & ~new_n32663_;
  assign new_n32779_ = ~new_n32777_ & ~new_n32778_;
  assign new_n32780_ = ~new_n32710_ & ~new_n32779_;
  assign new_n32781_ = ~new_n32453_ & ~new_n32709_;
  assign new_n32782_ = ~new_n32708_ & new_n32781_;
  assign new_n32783_ = ~new_n32780_ & ~new_n32782_;
  assign new_n32784_ = ~\b[17]  & ~new_n32783_;
  assign new_n32785_ = ~new_n32472_ & new_n32658_;
  assign new_n32786_ = ~new_n32654_ & new_n32785_;
  assign new_n32787_ = ~new_n32655_ & ~new_n32658_;
  assign new_n32788_ = ~new_n32786_ & ~new_n32787_;
  assign new_n32789_ = ~new_n32710_ & ~new_n32788_;
  assign new_n32790_ = ~new_n32462_ & ~new_n32709_;
  assign new_n32791_ = ~new_n32708_ & new_n32790_;
  assign new_n32792_ = ~new_n32789_ & ~new_n32791_;
  assign new_n32793_ = ~\b[16]  & ~new_n32792_;
  assign new_n32794_ = ~new_n32481_ & new_n32653_;
  assign new_n32795_ = ~new_n32649_ & new_n32794_;
  assign new_n32796_ = ~new_n32650_ & ~new_n32653_;
  assign new_n32797_ = ~new_n32795_ & ~new_n32796_;
  assign new_n32798_ = ~new_n32710_ & ~new_n32797_;
  assign new_n32799_ = ~new_n32471_ & ~new_n32709_;
  assign new_n32800_ = ~new_n32708_ & new_n32799_;
  assign new_n32801_ = ~new_n32798_ & ~new_n32800_;
  assign new_n32802_ = ~\b[15]  & ~new_n32801_;
  assign new_n32803_ = ~new_n32490_ & new_n32648_;
  assign new_n32804_ = ~new_n32644_ & new_n32803_;
  assign new_n32805_ = ~new_n32645_ & ~new_n32648_;
  assign new_n32806_ = ~new_n32804_ & ~new_n32805_;
  assign new_n32807_ = ~new_n32710_ & ~new_n32806_;
  assign new_n32808_ = ~new_n32480_ & ~new_n32709_;
  assign new_n32809_ = ~new_n32708_ & new_n32808_;
  assign new_n32810_ = ~new_n32807_ & ~new_n32809_;
  assign new_n32811_ = ~\b[14]  & ~new_n32810_;
  assign new_n32812_ = ~new_n32499_ & new_n32643_;
  assign new_n32813_ = ~new_n32639_ & new_n32812_;
  assign new_n32814_ = ~new_n32640_ & ~new_n32643_;
  assign new_n32815_ = ~new_n32813_ & ~new_n32814_;
  assign new_n32816_ = ~new_n32710_ & ~new_n32815_;
  assign new_n32817_ = ~new_n32489_ & ~new_n32709_;
  assign new_n32818_ = ~new_n32708_ & new_n32817_;
  assign new_n32819_ = ~new_n32816_ & ~new_n32818_;
  assign new_n32820_ = ~\b[13]  & ~new_n32819_;
  assign new_n32821_ = ~new_n32508_ & new_n32638_;
  assign new_n32822_ = ~new_n32634_ & new_n32821_;
  assign new_n32823_ = ~new_n32635_ & ~new_n32638_;
  assign new_n32824_ = ~new_n32822_ & ~new_n32823_;
  assign new_n32825_ = ~new_n32710_ & ~new_n32824_;
  assign new_n32826_ = ~new_n32498_ & ~new_n32709_;
  assign new_n32827_ = ~new_n32708_ & new_n32826_;
  assign new_n32828_ = ~new_n32825_ & ~new_n32827_;
  assign new_n32829_ = ~\b[12]  & ~new_n32828_;
  assign new_n32830_ = ~new_n32517_ & new_n32633_;
  assign new_n32831_ = ~new_n32629_ & new_n32830_;
  assign new_n32832_ = ~new_n32630_ & ~new_n32633_;
  assign new_n32833_ = ~new_n32831_ & ~new_n32832_;
  assign new_n32834_ = ~new_n32710_ & ~new_n32833_;
  assign new_n32835_ = ~new_n32507_ & ~new_n32709_;
  assign new_n32836_ = ~new_n32708_ & new_n32835_;
  assign new_n32837_ = ~new_n32834_ & ~new_n32836_;
  assign new_n32838_ = ~\b[11]  & ~new_n32837_;
  assign new_n32839_ = ~new_n32526_ & new_n32628_;
  assign new_n32840_ = ~new_n32624_ & new_n32839_;
  assign new_n32841_ = ~new_n32625_ & ~new_n32628_;
  assign new_n32842_ = ~new_n32840_ & ~new_n32841_;
  assign new_n32843_ = ~new_n32710_ & ~new_n32842_;
  assign new_n32844_ = ~new_n32516_ & ~new_n32709_;
  assign new_n32845_ = ~new_n32708_ & new_n32844_;
  assign new_n32846_ = ~new_n32843_ & ~new_n32845_;
  assign new_n32847_ = ~\b[10]  & ~new_n32846_;
  assign new_n32848_ = ~new_n32535_ & new_n32623_;
  assign new_n32849_ = ~new_n32619_ & new_n32848_;
  assign new_n32850_ = ~new_n32620_ & ~new_n32623_;
  assign new_n32851_ = ~new_n32849_ & ~new_n32850_;
  assign new_n32852_ = ~new_n32710_ & ~new_n32851_;
  assign new_n32853_ = ~new_n32525_ & ~new_n32709_;
  assign new_n32854_ = ~new_n32708_ & new_n32853_;
  assign new_n32855_ = ~new_n32852_ & ~new_n32854_;
  assign new_n32856_ = ~\b[9]  & ~new_n32855_;
  assign new_n32857_ = ~new_n32544_ & new_n32618_;
  assign new_n32858_ = ~new_n32614_ & new_n32857_;
  assign new_n32859_ = ~new_n32615_ & ~new_n32618_;
  assign new_n32860_ = ~new_n32858_ & ~new_n32859_;
  assign new_n32861_ = ~new_n32710_ & ~new_n32860_;
  assign new_n32862_ = ~new_n32534_ & ~new_n32709_;
  assign new_n32863_ = ~new_n32708_ & new_n32862_;
  assign new_n32864_ = ~new_n32861_ & ~new_n32863_;
  assign new_n32865_ = ~\b[8]  & ~new_n32864_;
  assign new_n32866_ = ~new_n32553_ & new_n32613_;
  assign new_n32867_ = ~new_n32609_ & new_n32866_;
  assign new_n32868_ = ~new_n32610_ & ~new_n32613_;
  assign new_n32869_ = ~new_n32867_ & ~new_n32868_;
  assign new_n32870_ = ~new_n32710_ & ~new_n32869_;
  assign new_n32871_ = ~new_n32543_ & ~new_n32709_;
  assign new_n32872_ = ~new_n32708_ & new_n32871_;
  assign new_n32873_ = ~new_n32870_ & ~new_n32872_;
  assign new_n32874_ = ~\b[7]  & ~new_n32873_;
  assign new_n32875_ = ~new_n32562_ & new_n32608_;
  assign new_n32876_ = ~new_n32604_ & new_n32875_;
  assign new_n32877_ = ~new_n32605_ & ~new_n32608_;
  assign new_n32878_ = ~new_n32876_ & ~new_n32877_;
  assign new_n32879_ = ~new_n32710_ & ~new_n32878_;
  assign new_n32880_ = ~new_n32552_ & ~new_n32709_;
  assign new_n32881_ = ~new_n32708_ & new_n32880_;
  assign new_n32882_ = ~new_n32879_ & ~new_n32881_;
  assign new_n32883_ = ~\b[6]  & ~new_n32882_;
  assign new_n32884_ = ~new_n32571_ & new_n32603_;
  assign new_n32885_ = ~new_n32599_ & new_n32884_;
  assign new_n32886_ = ~new_n32600_ & ~new_n32603_;
  assign new_n32887_ = ~new_n32885_ & ~new_n32886_;
  assign new_n32888_ = ~new_n32710_ & ~new_n32887_;
  assign new_n32889_ = ~new_n32561_ & ~new_n32709_;
  assign new_n32890_ = ~new_n32708_ & new_n32889_;
  assign new_n32891_ = ~new_n32888_ & ~new_n32890_;
  assign new_n32892_ = ~\b[5]  & ~new_n32891_;
  assign new_n32893_ = ~new_n32579_ & new_n32598_;
  assign new_n32894_ = ~new_n32594_ & new_n32893_;
  assign new_n32895_ = ~new_n32595_ & ~new_n32598_;
  assign new_n32896_ = ~new_n32894_ & ~new_n32895_;
  assign new_n32897_ = ~new_n32710_ & ~new_n32896_;
  assign new_n32898_ = ~new_n32570_ & ~new_n32709_;
  assign new_n32899_ = ~new_n32708_ & new_n32898_;
  assign new_n32900_ = ~new_n32897_ & ~new_n32899_;
  assign new_n32901_ = ~\b[4]  & ~new_n32900_;
  assign new_n32902_ = ~new_n32589_ & new_n32593_;
  assign new_n32903_ = ~new_n32588_ & new_n32902_;
  assign new_n32904_ = ~new_n32590_ & ~new_n32593_;
  assign new_n32905_ = ~new_n32903_ & ~new_n32904_;
  assign new_n32906_ = ~new_n32710_ & ~new_n32905_;
  assign new_n32907_ = ~new_n32578_ & ~new_n32709_;
  assign new_n32908_ = ~new_n32708_ & new_n32907_;
  assign new_n32909_ = ~new_n32906_ & ~new_n32908_;
  assign new_n32910_ = ~\b[3]  & ~new_n32909_;
  assign new_n32911_ = new_n4351_ & ~new_n32586_;
  assign new_n32912_ = ~new_n32584_ & new_n32911_;
  assign new_n32913_ = ~new_n32588_ & ~new_n32912_;
  assign new_n32914_ = ~new_n32710_ & new_n32913_;
  assign new_n32915_ = ~new_n32583_ & ~new_n32709_;
  assign new_n32916_ = ~new_n32708_ & new_n32915_;
  assign new_n32917_ = ~new_n32914_ & ~new_n32916_;
  assign new_n32918_ = ~\b[2]  & ~new_n32917_;
  assign new_n32919_ = \b[0]  & ~new_n32710_;
  assign new_n32920_ = \a[40]  & ~new_n32919_;
  assign new_n32921_ = new_n4351_ & ~new_n32710_;
  assign new_n32922_ = ~new_n32920_ & ~new_n32921_;
  assign new_n32923_ = \b[1]  & ~new_n32922_;
  assign new_n32924_ = ~\b[1]  & ~new_n32921_;
  assign new_n32925_ = ~new_n32920_ & new_n32924_;
  assign new_n32926_ = ~new_n32923_ & ~new_n32925_;
  assign new_n32927_ = ~new_n4693_ & ~new_n32926_;
  assign new_n32928_ = ~\b[1]  & ~new_n32922_;
  assign new_n32929_ = ~new_n32927_ & ~new_n32928_;
  assign new_n32930_ = \b[2]  & ~new_n32916_;
  assign new_n32931_ = ~new_n32914_ & new_n32930_;
  assign new_n32932_ = ~new_n32918_ & ~new_n32931_;
  assign new_n32933_ = ~new_n32929_ & new_n32932_;
  assign new_n32934_ = ~new_n32918_ & ~new_n32933_;
  assign new_n32935_ = \b[3]  & ~new_n32908_;
  assign new_n32936_ = ~new_n32906_ & new_n32935_;
  assign new_n32937_ = ~new_n32910_ & ~new_n32936_;
  assign new_n32938_ = ~new_n32934_ & new_n32937_;
  assign new_n32939_ = ~new_n32910_ & ~new_n32938_;
  assign new_n32940_ = \b[4]  & ~new_n32899_;
  assign new_n32941_ = ~new_n32897_ & new_n32940_;
  assign new_n32942_ = ~new_n32901_ & ~new_n32941_;
  assign new_n32943_ = ~new_n32939_ & new_n32942_;
  assign new_n32944_ = ~new_n32901_ & ~new_n32943_;
  assign new_n32945_ = \b[5]  & ~new_n32890_;
  assign new_n32946_ = ~new_n32888_ & new_n32945_;
  assign new_n32947_ = ~new_n32892_ & ~new_n32946_;
  assign new_n32948_ = ~new_n32944_ & new_n32947_;
  assign new_n32949_ = ~new_n32892_ & ~new_n32948_;
  assign new_n32950_ = \b[6]  & ~new_n32881_;
  assign new_n32951_ = ~new_n32879_ & new_n32950_;
  assign new_n32952_ = ~new_n32883_ & ~new_n32951_;
  assign new_n32953_ = ~new_n32949_ & new_n32952_;
  assign new_n32954_ = ~new_n32883_ & ~new_n32953_;
  assign new_n32955_ = \b[7]  & ~new_n32872_;
  assign new_n32956_ = ~new_n32870_ & new_n32955_;
  assign new_n32957_ = ~new_n32874_ & ~new_n32956_;
  assign new_n32958_ = ~new_n32954_ & new_n32957_;
  assign new_n32959_ = ~new_n32874_ & ~new_n32958_;
  assign new_n32960_ = \b[8]  & ~new_n32863_;
  assign new_n32961_ = ~new_n32861_ & new_n32960_;
  assign new_n32962_ = ~new_n32865_ & ~new_n32961_;
  assign new_n32963_ = ~new_n32959_ & new_n32962_;
  assign new_n32964_ = ~new_n32865_ & ~new_n32963_;
  assign new_n32965_ = \b[9]  & ~new_n32854_;
  assign new_n32966_ = ~new_n32852_ & new_n32965_;
  assign new_n32967_ = ~new_n32856_ & ~new_n32966_;
  assign new_n32968_ = ~new_n32964_ & new_n32967_;
  assign new_n32969_ = ~new_n32856_ & ~new_n32968_;
  assign new_n32970_ = \b[10]  & ~new_n32845_;
  assign new_n32971_ = ~new_n32843_ & new_n32970_;
  assign new_n32972_ = ~new_n32847_ & ~new_n32971_;
  assign new_n32973_ = ~new_n32969_ & new_n32972_;
  assign new_n32974_ = ~new_n32847_ & ~new_n32973_;
  assign new_n32975_ = \b[11]  & ~new_n32836_;
  assign new_n32976_ = ~new_n32834_ & new_n32975_;
  assign new_n32977_ = ~new_n32838_ & ~new_n32976_;
  assign new_n32978_ = ~new_n32974_ & new_n32977_;
  assign new_n32979_ = ~new_n32838_ & ~new_n32978_;
  assign new_n32980_ = \b[12]  & ~new_n32827_;
  assign new_n32981_ = ~new_n32825_ & new_n32980_;
  assign new_n32982_ = ~new_n32829_ & ~new_n32981_;
  assign new_n32983_ = ~new_n32979_ & new_n32982_;
  assign new_n32984_ = ~new_n32829_ & ~new_n32983_;
  assign new_n32985_ = \b[13]  & ~new_n32818_;
  assign new_n32986_ = ~new_n32816_ & new_n32985_;
  assign new_n32987_ = ~new_n32820_ & ~new_n32986_;
  assign new_n32988_ = ~new_n32984_ & new_n32987_;
  assign new_n32989_ = ~new_n32820_ & ~new_n32988_;
  assign new_n32990_ = \b[14]  & ~new_n32809_;
  assign new_n32991_ = ~new_n32807_ & new_n32990_;
  assign new_n32992_ = ~new_n32811_ & ~new_n32991_;
  assign new_n32993_ = ~new_n32989_ & new_n32992_;
  assign new_n32994_ = ~new_n32811_ & ~new_n32993_;
  assign new_n32995_ = \b[15]  & ~new_n32800_;
  assign new_n32996_ = ~new_n32798_ & new_n32995_;
  assign new_n32997_ = ~new_n32802_ & ~new_n32996_;
  assign new_n32998_ = ~new_n32994_ & new_n32997_;
  assign new_n32999_ = ~new_n32802_ & ~new_n32998_;
  assign new_n33000_ = \b[16]  & ~new_n32791_;
  assign new_n33001_ = ~new_n32789_ & new_n33000_;
  assign new_n33002_ = ~new_n32793_ & ~new_n33001_;
  assign new_n33003_ = ~new_n32999_ & new_n33002_;
  assign new_n33004_ = ~new_n32793_ & ~new_n33003_;
  assign new_n33005_ = \b[17]  & ~new_n32782_;
  assign new_n33006_ = ~new_n32780_ & new_n33005_;
  assign new_n33007_ = ~new_n32784_ & ~new_n33006_;
  assign new_n33008_ = ~new_n33004_ & new_n33007_;
  assign new_n33009_ = ~new_n32784_ & ~new_n33008_;
  assign new_n33010_ = \b[18]  & ~new_n32773_;
  assign new_n33011_ = ~new_n32771_ & new_n33010_;
  assign new_n33012_ = ~new_n32775_ & ~new_n33011_;
  assign new_n33013_ = ~new_n33009_ & new_n33012_;
  assign new_n33014_ = ~new_n32775_ & ~new_n33013_;
  assign new_n33015_ = \b[19]  & ~new_n32764_;
  assign new_n33016_ = ~new_n32762_ & new_n33015_;
  assign new_n33017_ = ~new_n32766_ & ~new_n33016_;
  assign new_n33018_ = ~new_n33014_ & new_n33017_;
  assign new_n33019_ = ~new_n32766_ & ~new_n33018_;
  assign new_n33020_ = \b[20]  & ~new_n32755_;
  assign new_n33021_ = ~new_n32753_ & new_n33020_;
  assign new_n33022_ = ~new_n32757_ & ~new_n33021_;
  assign new_n33023_ = ~new_n33019_ & new_n33022_;
  assign new_n33024_ = ~new_n32757_ & ~new_n33023_;
  assign new_n33025_ = \b[21]  & ~new_n32746_;
  assign new_n33026_ = ~new_n32744_ & new_n33025_;
  assign new_n33027_ = ~new_n32748_ & ~new_n33026_;
  assign new_n33028_ = ~new_n33024_ & new_n33027_;
  assign new_n33029_ = ~new_n32748_ & ~new_n33028_;
  assign new_n33030_ = \b[22]  & ~new_n32737_;
  assign new_n33031_ = ~new_n32735_ & new_n33030_;
  assign new_n33032_ = ~new_n32739_ & ~new_n33031_;
  assign new_n33033_ = ~new_n33029_ & new_n33032_;
  assign new_n33034_ = ~new_n32739_ & ~new_n33033_;
  assign new_n33035_ = \b[23]  & ~new_n32717_;
  assign new_n33036_ = ~new_n32715_ & new_n33035_;
  assign new_n33037_ = ~new_n32730_ & ~new_n33036_;
  assign new_n33038_ = ~new_n33034_ & new_n33037_;
  assign new_n33039_ = ~new_n32730_ & ~new_n33038_;
  assign new_n33040_ = \b[24]  & ~new_n32727_;
  assign new_n33041_ = ~new_n32725_ & new_n33040_;
  assign new_n33042_ = ~new_n32729_ & ~new_n33041_;
  assign new_n33043_ = ~new_n33039_ & new_n33042_;
  assign new_n33044_ = ~new_n32729_ & ~new_n33043_;
  assign new_n33045_ = new_n4813_ & ~new_n33044_;
  assign new_n33046_ = ~new_n32718_ & ~new_n33045_;
  assign new_n33047_ = ~new_n32739_ & new_n33037_;
  assign new_n33048_ = ~new_n33033_ & new_n33047_;
  assign new_n33049_ = ~new_n33034_ & ~new_n33037_;
  assign new_n33050_ = ~new_n33048_ & ~new_n33049_;
  assign new_n33051_ = new_n4813_ & ~new_n33050_;
  assign new_n33052_ = ~new_n33044_ & new_n33051_;
  assign new_n33053_ = ~new_n33046_ & ~new_n33052_;
  assign new_n33054_ = ~new_n32728_ & ~new_n33045_;
  assign new_n33055_ = ~new_n32730_ & new_n33042_;
  assign new_n33056_ = ~new_n33038_ & new_n33055_;
  assign new_n33057_ = ~new_n33039_ & ~new_n33042_;
  assign new_n33058_ = ~new_n33056_ & ~new_n33057_;
  assign new_n33059_ = new_n33045_ & ~new_n33058_;
  assign new_n33060_ = ~new_n33054_ & ~new_n33059_;
  assign new_n33061_ = ~\b[25]  & ~new_n33060_;
  assign new_n33062_ = ~\b[24]  & ~new_n33053_;
  assign new_n33063_ = ~new_n32738_ & ~new_n33045_;
  assign new_n33064_ = ~new_n32748_ & new_n33032_;
  assign new_n33065_ = ~new_n33028_ & new_n33064_;
  assign new_n33066_ = ~new_n33029_ & ~new_n33032_;
  assign new_n33067_ = ~new_n33065_ & ~new_n33066_;
  assign new_n33068_ = new_n4813_ & ~new_n33067_;
  assign new_n33069_ = ~new_n33044_ & new_n33068_;
  assign new_n33070_ = ~new_n33063_ & ~new_n33069_;
  assign new_n33071_ = ~\b[23]  & ~new_n33070_;
  assign new_n33072_ = ~new_n32747_ & ~new_n33045_;
  assign new_n33073_ = ~new_n32757_ & new_n33027_;
  assign new_n33074_ = ~new_n33023_ & new_n33073_;
  assign new_n33075_ = ~new_n33024_ & ~new_n33027_;
  assign new_n33076_ = ~new_n33074_ & ~new_n33075_;
  assign new_n33077_ = new_n4813_ & ~new_n33076_;
  assign new_n33078_ = ~new_n33044_ & new_n33077_;
  assign new_n33079_ = ~new_n33072_ & ~new_n33078_;
  assign new_n33080_ = ~\b[22]  & ~new_n33079_;
  assign new_n33081_ = ~new_n32756_ & ~new_n33045_;
  assign new_n33082_ = ~new_n32766_ & new_n33022_;
  assign new_n33083_ = ~new_n33018_ & new_n33082_;
  assign new_n33084_ = ~new_n33019_ & ~new_n33022_;
  assign new_n33085_ = ~new_n33083_ & ~new_n33084_;
  assign new_n33086_ = new_n4813_ & ~new_n33085_;
  assign new_n33087_ = ~new_n33044_ & new_n33086_;
  assign new_n33088_ = ~new_n33081_ & ~new_n33087_;
  assign new_n33089_ = ~\b[21]  & ~new_n33088_;
  assign new_n33090_ = ~new_n32765_ & ~new_n33045_;
  assign new_n33091_ = ~new_n32775_ & new_n33017_;
  assign new_n33092_ = ~new_n33013_ & new_n33091_;
  assign new_n33093_ = ~new_n33014_ & ~new_n33017_;
  assign new_n33094_ = ~new_n33092_ & ~new_n33093_;
  assign new_n33095_ = new_n4813_ & ~new_n33094_;
  assign new_n33096_ = ~new_n33044_ & new_n33095_;
  assign new_n33097_ = ~new_n33090_ & ~new_n33096_;
  assign new_n33098_ = ~\b[20]  & ~new_n33097_;
  assign new_n33099_ = ~new_n32774_ & ~new_n33045_;
  assign new_n33100_ = ~new_n32784_ & new_n33012_;
  assign new_n33101_ = ~new_n33008_ & new_n33100_;
  assign new_n33102_ = ~new_n33009_ & ~new_n33012_;
  assign new_n33103_ = ~new_n33101_ & ~new_n33102_;
  assign new_n33104_ = new_n4813_ & ~new_n33103_;
  assign new_n33105_ = ~new_n33044_ & new_n33104_;
  assign new_n33106_ = ~new_n33099_ & ~new_n33105_;
  assign new_n33107_ = ~\b[19]  & ~new_n33106_;
  assign new_n33108_ = ~new_n32783_ & ~new_n33045_;
  assign new_n33109_ = ~new_n32793_ & new_n33007_;
  assign new_n33110_ = ~new_n33003_ & new_n33109_;
  assign new_n33111_ = ~new_n33004_ & ~new_n33007_;
  assign new_n33112_ = ~new_n33110_ & ~new_n33111_;
  assign new_n33113_ = new_n4813_ & ~new_n33112_;
  assign new_n33114_ = ~new_n33044_ & new_n33113_;
  assign new_n33115_ = ~new_n33108_ & ~new_n33114_;
  assign new_n33116_ = ~\b[18]  & ~new_n33115_;
  assign new_n33117_ = ~new_n32792_ & ~new_n33045_;
  assign new_n33118_ = ~new_n32802_ & new_n33002_;
  assign new_n33119_ = ~new_n32998_ & new_n33118_;
  assign new_n33120_ = ~new_n32999_ & ~new_n33002_;
  assign new_n33121_ = ~new_n33119_ & ~new_n33120_;
  assign new_n33122_ = new_n4813_ & ~new_n33121_;
  assign new_n33123_ = ~new_n33044_ & new_n33122_;
  assign new_n33124_ = ~new_n33117_ & ~new_n33123_;
  assign new_n33125_ = ~\b[17]  & ~new_n33124_;
  assign new_n33126_ = ~new_n32801_ & ~new_n33045_;
  assign new_n33127_ = ~new_n32811_ & new_n32997_;
  assign new_n33128_ = ~new_n32993_ & new_n33127_;
  assign new_n33129_ = ~new_n32994_ & ~new_n32997_;
  assign new_n33130_ = ~new_n33128_ & ~new_n33129_;
  assign new_n33131_ = new_n4813_ & ~new_n33130_;
  assign new_n33132_ = ~new_n33044_ & new_n33131_;
  assign new_n33133_ = ~new_n33126_ & ~new_n33132_;
  assign new_n33134_ = ~\b[16]  & ~new_n33133_;
  assign new_n33135_ = ~new_n32810_ & ~new_n33045_;
  assign new_n33136_ = ~new_n32820_ & new_n32992_;
  assign new_n33137_ = ~new_n32988_ & new_n33136_;
  assign new_n33138_ = ~new_n32989_ & ~new_n32992_;
  assign new_n33139_ = ~new_n33137_ & ~new_n33138_;
  assign new_n33140_ = new_n4813_ & ~new_n33139_;
  assign new_n33141_ = ~new_n33044_ & new_n33140_;
  assign new_n33142_ = ~new_n33135_ & ~new_n33141_;
  assign new_n33143_ = ~\b[15]  & ~new_n33142_;
  assign new_n33144_ = ~new_n32819_ & ~new_n33045_;
  assign new_n33145_ = ~new_n32829_ & new_n32987_;
  assign new_n33146_ = ~new_n32983_ & new_n33145_;
  assign new_n33147_ = ~new_n32984_ & ~new_n32987_;
  assign new_n33148_ = ~new_n33146_ & ~new_n33147_;
  assign new_n33149_ = new_n4813_ & ~new_n33148_;
  assign new_n33150_ = ~new_n33044_ & new_n33149_;
  assign new_n33151_ = ~new_n33144_ & ~new_n33150_;
  assign new_n33152_ = ~\b[14]  & ~new_n33151_;
  assign new_n33153_ = ~new_n32828_ & ~new_n33045_;
  assign new_n33154_ = ~new_n32838_ & new_n32982_;
  assign new_n33155_ = ~new_n32978_ & new_n33154_;
  assign new_n33156_ = ~new_n32979_ & ~new_n32982_;
  assign new_n33157_ = ~new_n33155_ & ~new_n33156_;
  assign new_n33158_ = new_n4813_ & ~new_n33157_;
  assign new_n33159_ = ~new_n33044_ & new_n33158_;
  assign new_n33160_ = ~new_n33153_ & ~new_n33159_;
  assign new_n33161_ = ~\b[13]  & ~new_n33160_;
  assign new_n33162_ = ~new_n32837_ & ~new_n33045_;
  assign new_n33163_ = ~new_n32847_ & new_n32977_;
  assign new_n33164_ = ~new_n32973_ & new_n33163_;
  assign new_n33165_ = ~new_n32974_ & ~new_n32977_;
  assign new_n33166_ = ~new_n33164_ & ~new_n33165_;
  assign new_n33167_ = new_n4813_ & ~new_n33166_;
  assign new_n33168_ = ~new_n33044_ & new_n33167_;
  assign new_n33169_ = ~new_n33162_ & ~new_n33168_;
  assign new_n33170_ = ~\b[12]  & ~new_n33169_;
  assign new_n33171_ = ~new_n32846_ & ~new_n33045_;
  assign new_n33172_ = ~new_n32856_ & new_n32972_;
  assign new_n33173_ = ~new_n32968_ & new_n33172_;
  assign new_n33174_ = ~new_n32969_ & ~new_n32972_;
  assign new_n33175_ = ~new_n33173_ & ~new_n33174_;
  assign new_n33176_ = new_n4813_ & ~new_n33175_;
  assign new_n33177_ = ~new_n33044_ & new_n33176_;
  assign new_n33178_ = ~new_n33171_ & ~new_n33177_;
  assign new_n33179_ = ~\b[11]  & ~new_n33178_;
  assign new_n33180_ = ~new_n32855_ & ~new_n33045_;
  assign new_n33181_ = ~new_n32865_ & new_n32967_;
  assign new_n33182_ = ~new_n32963_ & new_n33181_;
  assign new_n33183_ = ~new_n32964_ & ~new_n32967_;
  assign new_n33184_ = ~new_n33182_ & ~new_n33183_;
  assign new_n33185_ = new_n4813_ & ~new_n33184_;
  assign new_n33186_ = ~new_n33044_ & new_n33185_;
  assign new_n33187_ = ~new_n33180_ & ~new_n33186_;
  assign new_n33188_ = ~\b[10]  & ~new_n33187_;
  assign new_n33189_ = ~new_n32864_ & ~new_n33045_;
  assign new_n33190_ = ~new_n32874_ & new_n32962_;
  assign new_n33191_ = ~new_n32958_ & new_n33190_;
  assign new_n33192_ = ~new_n32959_ & ~new_n32962_;
  assign new_n33193_ = ~new_n33191_ & ~new_n33192_;
  assign new_n33194_ = new_n4813_ & ~new_n33193_;
  assign new_n33195_ = ~new_n33044_ & new_n33194_;
  assign new_n33196_ = ~new_n33189_ & ~new_n33195_;
  assign new_n33197_ = ~\b[9]  & ~new_n33196_;
  assign new_n33198_ = ~new_n32873_ & ~new_n33045_;
  assign new_n33199_ = ~new_n32883_ & new_n32957_;
  assign new_n33200_ = ~new_n32953_ & new_n33199_;
  assign new_n33201_ = ~new_n32954_ & ~new_n32957_;
  assign new_n33202_ = ~new_n33200_ & ~new_n33201_;
  assign new_n33203_ = new_n4813_ & ~new_n33202_;
  assign new_n33204_ = ~new_n33044_ & new_n33203_;
  assign new_n33205_ = ~new_n33198_ & ~new_n33204_;
  assign new_n33206_ = ~\b[8]  & ~new_n33205_;
  assign new_n33207_ = ~new_n32882_ & ~new_n33045_;
  assign new_n33208_ = ~new_n32892_ & new_n32952_;
  assign new_n33209_ = ~new_n32948_ & new_n33208_;
  assign new_n33210_ = ~new_n32949_ & ~new_n32952_;
  assign new_n33211_ = ~new_n33209_ & ~new_n33210_;
  assign new_n33212_ = new_n4813_ & ~new_n33211_;
  assign new_n33213_ = ~new_n33044_ & new_n33212_;
  assign new_n33214_ = ~new_n33207_ & ~new_n33213_;
  assign new_n33215_ = ~\b[7]  & ~new_n33214_;
  assign new_n33216_ = ~new_n32891_ & ~new_n33045_;
  assign new_n33217_ = ~new_n32901_ & new_n32947_;
  assign new_n33218_ = ~new_n32943_ & new_n33217_;
  assign new_n33219_ = ~new_n32944_ & ~new_n32947_;
  assign new_n33220_ = ~new_n33218_ & ~new_n33219_;
  assign new_n33221_ = new_n4813_ & ~new_n33220_;
  assign new_n33222_ = ~new_n33044_ & new_n33221_;
  assign new_n33223_ = ~new_n33216_ & ~new_n33222_;
  assign new_n33224_ = ~\b[6]  & ~new_n33223_;
  assign new_n33225_ = ~new_n32900_ & ~new_n33045_;
  assign new_n33226_ = ~new_n32910_ & new_n32942_;
  assign new_n33227_ = ~new_n32938_ & new_n33226_;
  assign new_n33228_ = ~new_n32939_ & ~new_n32942_;
  assign new_n33229_ = ~new_n33227_ & ~new_n33228_;
  assign new_n33230_ = new_n4813_ & ~new_n33229_;
  assign new_n33231_ = ~new_n33044_ & new_n33230_;
  assign new_n33232_ = ~new_n33225_ & ~new_n33231_;
  assign new_n33233_ = ~\b[5]  & ~new_n33232_;
  assign new_n33234_ = ~new_n32909_ & ~new_n33045_;
  assign new_n33235_ = ~new_n32918_ & new_n32937_;
  assign new_n33236_ = ~new_n32933_ & new_n33235_;
  assign new_n33237_ = ~new_n32934_ & ~new_n32937_;
  assign new_n33238_ = ~new_n33236_ & ~new_n33237_;
  assign new_n33239_ = new_n4813_ & ~new_n33238_;
  assign new_n33240_ = ~new_n33044_ & new_n33239_;
  assign new_n33241_ = ~new_n33234_ & ~new_n33240_;
  assign new_n33242_ = ~\b[4]  & ~new_n33241_;
  assign new_n33243_ = ~new_n32917_ & ~new_n33045_;
  assign new_n33244_ = ~new_n32928_ & new_n32932_;
  assign new_n33245_ = ~new_n32927_ & new_n33244_;
  assign new_n33246_ = ~new_n32929_ & ~new_n32932_;
  assign new_n33247_ = ~new_n33245_ & ~new_n33246_;
  assign new_n33248_ = new_n4813_ & ~new_n33247_;
  assign new_n33249_ = ~new_n33044_ & new_n33248_;
  assign new_n33250_ = ~new_n33243_ & ~new_n33249_;
  assign new_n33251_ = ~\b[3]  & ~new_n33250_;
  assign new_n33252_ = ~new_n32922_ & ~new_n33045_;
  assign new_n33253_ = new_n4693_ & ~new_n32925_;
  assign new_n33254_ = ~new_n32923_ & new_n33253_;
  assign new_n33255_ = new_n4813_ & ~new_n33254_;
  assign new_n33256_ = ~new_n32927_ & new_n33255_;
  assign new_n33257_ = ~new_n33044_ & new_n33256_;
  assign new_n33258_ = ~new_n33252_ & ~new_n33257_;
  assign new_n33259_ = ~\b[2]  & ~new_n33258_;
  assign new_n33260_ = new_n5033_ & ~new_n33044_;
  assign new_n33261_ = \a[39]  & ~new_n33260_;
  assign new_n33262_ = new_n5039_ & ~new_n33044_;
  assign new_n33263_ = ~new_n33261_ & ~new_n33262_;
  assign new_n33264_ = \b[1]  & ~new_n33263_;
  assign new_n33265_ = ~\b[1]  & ~new_n33262_;
  assign new_n33266_ = ~new_n33261_ & new_n33265_;
  assign new_n33267_ = ~new_n33264_ & ~new_n33266_;
  assign new_n33268_ = ~new_n5046_ & ~new_n33267_;
  assign new_n33269_ = ~\b[1]  & ~new_n33263_;
  assign new_n33270_ = ~new_n33268_ & ~new_n33269_;
  assign new_n33271_ = \b[2]  & ~new_n33257_;
  assign new_n33272_ = ~new_n33252_ & new_n33271_;
  assign new_n33273_ = ~new_n33259_ & ~new_n33272_;
  assign new_n33274_ = ~new_n33270_ & new_n33273_;
  assign new_n33275_ = ~new_n33259_ & ~new_n33274_;
  assign new_n33276_ = \b[3]  & ~new_n33249_;
  assign new_n33277_ = ~new_n33243_ & new_n33276_;
  assign new_n33278_ = ~new_n33251_ & ~new_n33277_;
  assign new_n33279_ = ~new_n33275_ & new_n33278_;
  assign new_n33280_ = ~new_n33251_ & ~new_n33279_;
  assign new_n33281_ = \b[4]  & ~new_n33240_;
  assign new_n33282_ = ~new_n33234_ & new_n33281_;
  assign new_n33283_ = ~new_n33242_ & ~new_n33282_;
  assign new_n33284_ = ~new_n33280_ & new_n33283_;
  assign new_n33285_ = ~new_n33242_ & ~new_n33284_;
  assign new_n33286_ = \b[5]  & ~new_n33231_;
  assign new_n33287_ = ~new_n33225_ & new_n33286_;
  assign new_n33288_ = ~new_n33233_ & ~new_n33287_;
  assign new_n33289_ = ~new_n33285_ & new_n33288_;
  assign new_n33290_ = ~new_n33233_ & ~new_n33289_;
  assign new_n33291_ = \b[6]  & ~new_n33222_;
  assign new_n33292_ = ~new_n33216_ & new_n33291_;
  assign new_n33293_ = ~new_n33224_ & ~new_n33292_;
  assign new_n33294_ = ~new_n33290_ & new_n33293_;
  assign new_n33295_ = ~new_n33224_ & ~new_n33294_;
  assign new_n33296_ = \b[7]  & ~new_n33213_;
  assign new_n33297_ = ~new_n33207_ & new_n33296_;
  assign new_n33298_ = ~new_n33215_ & ~new_n33297_;
  assign new_n33299_ = ~new_n33295_ & new_n33298_;
  assign new_n33300_ = ~new_n33215_ & ~new_n33299_;
  assign new_n33301_ = \b[8]  & ~new_n33204_;
  assign new_n33302_ = ~new_n33198_ & new_n33301_;
  assign new_n33303_ = ~new_n33206_ & ~new_n33302_;
  assign new_n33304_ = ~new_n33300_ & new_n33303_;
  assign new_n33305_ = ~new_n33206_ & ~new_n33304_;
  assign new_n33306_ = \b[9]  & ~new_n33195_;
  assign new_n33307_ = ~new_n33189_ & new_n33306_;
  assign new_n33308_ = ~new_n33197_ & ~new_n33307_;
  assign new_n33309_ = ~new_n33305_ & new_n33308_;
  assign new_n33310_ = ~new_n33197_ & ~new_n33309_;
  assign new_n33311_ = \b[10]  & ~new_n33186_;
  assign new_n33312_ = ~new_n33180_ & new_n33311_;
  assign new_n33313_ = ~new_n33188_ & ~new_n33312_;
  assign new_n33314_ = ~new_n33310_ & new_n33313_;
  assign new_n33315_ = ~new_n33188_ & ~new_n33314_;
  assign new_n33316_ = \b[11]  & ~new_n33177_;
  assign new_n33317_ = ~new_n33171_ & new_n33316_;
  assign new_n33318_ = ~new_n33179_ & ~new_n33317_;
  assign new_n33319_ = ~new_n33315_ & new_n33318_;
  assign new_n33320_ = ~new_n33179_ & ~new_n33319_;
  assign new_n33321_ = \b[12]  & ~new_n33168_;
  assign new_n33322_ = ~new_n33162_ & new_n33321_;
  assign new_n33323_ = ~new_n33170_ & ~new_n33322_;
  assign new_n33324_ = ~new_n33320_ & new_n33323_;
  assign new_n33325_ = ~new_n33170_ & ~new_n33324_;
  assign new_n33326_ = \b[13]  & ~new_n33159_;
  assign new_n33327_ = ~new_n33153_ & new_n33326_;
  assign new_n33328_ = ~new_n33161_ & ~new_n33327_;
  assign new_n33329_ = ~new_n33325_ & new_n33328_;
  assign new_n33330_ = ~new_n33161_ & ~new_n33329_;
  assign new_n33331_ = \b[14]  & ~new_n33150_;
  assign new_n33332_ = ~new_n33144_ & new_n33331_;
  assign new_n33333_ = ~new_n33152_ & ~new_n33332_;
  assign new_n33334_ = ~new_n33330_ & new_n33333_;
  assign new_n33335_ = ~new_n33152_ & ~new_n33334_;
  assign new_n33336_ = \b[15]  & ~new_n33141_;
  assign new_n33337_ = ~new_n33135_ & new_n33336_;
  assign new_n33338_ = ~new_n33143_ & ~new_n33337_;
  assign new_n33339_ = ~new_n33335_ & new_n33338_;
  assign new_n33340_ = ~new_n33143_ & ~new_n33339_;
  assign new_n33341_ = \b[16]  & ~new_n33132_;
  assign new_n33342_ = ~new_n33126_ & new_n33341_;
  assign new_n33343_ = ~new_n33134_ & ~new_n33342_;
  assign new_n33344_ = ~new_n33340_ & new_n33343_;
  assign new_n33345_ = ~new_n33134_ & ~new_n33344_;
  assign new_n33346_ = \b[17]  & ~new_n33123_;
  assign new_n33347_ = ~new_n33117_ & new_n33346_;
  assign new_n33348_ = ~new_n33125_ & ~new_n33347_;
  assign new_n33349_ = ~new_n33345_ & new_n33348_;
  assign new_n33350_ = ~new_n33125_ & ~new_n33349_;
  assign new_n33351_ = \b[18]  & ~new_n33114_;
  assign new_n33352_ = ~new_n33108_ & new_n33351_;
  assign new_n33353_ = ~new_n33116_ & ~new_n33352_;
  assign new_n33354_ = ~new_n33350_ & new_n33353_;
  assign new_n33355_ = ~new_n33116_ & ~new_n33354_;
  assign new_n33356_ = \b[19]  & ~new_n33105_;
  assign new_n33357_ = ~new_n33099_ & new_n33356_;
  assign new_n33358_ = ~new_n33107_ & ~new_n33357_;
  assign new_n33359_ = ~new_n33355_ & new_n33358_;
  assign new_n33360_ = ~new_n33107_ & ~new_n33359_;
  assign new_n33361_ = \b[20]  & ~new_n33096_;
  assign new_n33362_ = ~new_n33090_ & new_n33361_;
  assign new_n33363_ = ~new_n33098_ & ~new_n33362_;
  assign new_n33364_ = ~new_n33360_ & new_n33363_;
  assign new_n33365_ = ~new_n33098_ & ~new_n33364_;
  assign new_n33366_ = \b[21]  & ~new_n33087_;
  assign new_n33367_ = ~new_n33081_ & new_n33366_;
  assign new_n33368_ = ~new_n33089_ & ~new_n33367_;
  assign new_n33369_ = ~new_n33365_ & new_n33368_;
  assign new_n33370_ = ~new_n33089_ & ~new_n33369_;
  assign new_n33371_ = \b[22]  & ~new_n33078_;
  assign new_n33372_ = ~new_n33072_ & new_n33371_;
  assign new_n33373_ = ~new_n33080_ & ~new_n33372_;
  assign new_n33374_ = ~new_n33370_ & new_n33373_;
  assign new_n33375_ = ~new_n33080_ & ~new_n33374_;
  assign new_n33376_ = \b[23]  & ~new_n33069_;
  assign new_n33377_ = ~new_n33063_ & new_n33376_;
  assign new_n33378_ = ~new_n33071_ & ~new_n33377_;
  assign new_n33379_ = ~new_n33375_ & new_n33378_;
  assign new_n33380_ = ~new_n33071_ & ~new_n33379_;
  assign new_n33381_ = \b[24]  & ~new_n33052_;
  assign new_n33382_ = ~new_n33046_ & new_n33381_;
  assign new_n33383_ = ~new_n33062_ & ~new_n33382_;
  assign new_n33384_ = ~new_n33380_ & new_n33383_;
  assign new_n33385_ = ~new_n33062_ & ~new_n33384_;
  assign new_n33386_ = \b[25]  & ~new_n33054_;
  assign new_n33387_ = ~new_n33059_ & new_n33386_;
  assign new_n33388_ = ~new_n33061_ & ~new_n33387_;
  assign new_n33389_ = ~new_n33385_ & new_n33388_;
  assign new_n33390_ = ~new_n33061_ & ~new_n33389_;
  assign new_n33391_ = new_n5172_ & ~new_n33390_;
  assign new_n33392_ = ~new_n33053_ & ~new_n33391_;
  assign new_n33393_ = ~new_n33071_ & new_n33383_;
  assign new_n33394_ = ~new_n33379_ & new_n33393_;
  assign new_n33395_ = ~new_n33380_ & ~new_n33383_;
  assign new_n33396_ = ~new_n33394_ & ~new_n33395_;
  assign new_n33397_ = new_n5172_ & ~new_n33396_;
  assign new_n33398_ = ~new_n33390_ & new_n33397_;
  assign new_n33399_ = ~new_n33392_ & ~new_n33398_;
  assign new_n33400_ = ~\b[25]  & ~new_n33399_;
  assign new_n33401_ = ~new_n33070_ & ~new_n33391_;
  assign new_n33402_ = ~new_n33080_ & new_n33378_;
  assign new_n33403_ = ~new_n33374_ & new_n33402_;
  assign new_n33404_ = ~new_n33375_ & ~new_n33378_;
  assign new_n33405_ = ~new_n33403_ & ~new_n33404_;
  assign new_n33406_ = new_n5172_ & ~new_n33405_;
  assign new_n33407_ = ~new_n33390_ & new_n33406_;
  assign new_n33408_ = ~new_n33401_ & ~new_n33407_;
  assign new_n33409_ = ~\b[24]  & ~new_n33408_;
  assign new_n33410_ = ~new_n33079_ & ~new_n33391_;
  assign new_n33411_ = ~new_n33089_ & new_n33373_;
  assign new_n33412_ = ~new_n33369_ & new_n33411_;
  assign new_n33413_ = ~new_n33370_ & ~new_n33373_;
  assign new_n33414_ = ~new_n33412_ & ~new_n33413_;
  assign new_n33415_ = new_n5172_ & ~new_n33414_;
  assign new_n33416_ = ~new_n33390_ & new_n33415_;
  assign new_n33417_ = ~new_n33410_ & ~new_n33416_;
  assign new_n33418_ = ~\b[23]  & ~new_n33417_;
  assign new_n33419_ = ~new_n33088_ & ~new_n33391_;
  assign new_n33420_ = ~new_n33098_ & new_n33368_;
  assign new_n33421_ = ~new_n33364_ & new_n33420_;
  assign new_n33422_ = ~new_n33365_ & ~new_n33368_;
  assign new_n33423_ = ~new_n33421_ & ~new_n33422_;
  assign new_n33424_ = new_n5172_ & ~new_n33423_;
  assign new_n33425_ = ~new_n33390_ & new_n33424_;
  assign new_n33426_ = ~new_n33419_ & ~new_n33425_;
  assign new_n33427_ = ~\b[22]  & ~new_n33426_;
  assign new_n33428_ = ~new_n33097_ & ~new_n33391_;
  assign new_n33429_ = ~new_n33107_ & new_n33363_;
  assign new_n33430_ = ~new_n33359_ & new_n33429_;
  assign new_n33431_ = ~new_n33360_ & ~new_n33363_;
  assign new_n33432_ = ~new_n33430_ & ~new_n33431_;
  assign new_n33433_ = new_n5172_ & ~new_n33432_;
  assign new_n33434_ = ~new_n33390_ & new_n33433_;
  assign new_n33435_ = ~new_n33428_ & ~new_n33434_;
  assign new_n33436_ = ~\b[21]  & ~new_n33435_;
  assign new_n33437_ = ~new_n33106_ & ~new_n33391_;
  assign new_n33438_ = ~new_n33116_ & new_n33358_;
  assign new_n33439_ = ~new_n33354_ & new_n33438_;
  assign new_n33440_ = ~new_n33355_ & ~new_n33358_;
  assign new_n33441_ = ~new_n33439_ & ~new_n33440_;
  assign new_n33442_ = new_n5172_ & ~new_n33441_;
  assign new_n33443_ = ~new_n33390_ & new_n33442_;
  assign new_n33444_ = ~new_n33437_ & ~new_n33443_;
  assign new_n33445_ = ~\b[20]  & ~new_n33444_;
  assign new_n33446_ = ~new_n33115_ & ~new_n33391_;
  assign new_n33447_ = ~new_n33125_ & new_n33353_;
  assign new_n33448_ = ~new_n33349_ & new_n33447_;
  assign new_n33449_ = ~new_n33350_ & ~new_n33353_;
  assign new_n33450_ = ~new_n33448_ & ~new_n33449_;
  assign new_n33451_ = new_n5172_ & ~new_n33450_;
  assign new_n33452_ = ~new_n33390_ & new_n33451_;
  assign new_n33453_ = ~new_n33446_ & ~new_n33452_;
  assign new_n33454_ = ~\b[19]  & ~new_n33453_;
  assign new_n33455_ = ~new_n33124_ & ~new_n33391_;
  assign new_n33456_ = ~new_n33134_ & new_n33348_;
  assign new_n33457_ = ~new_n33344_ & new_n33456_;
  assign new_n33458_ = ~new_n33345_ & ~new_n33348_;
  assign new_n33459_ = ~new_n33457_ & ~new_n33458_;
  assign new_n33460_ = new_n5172_ & ~new_n33459_;
  assign new_n33461_ = ~new_n33390_ & new_n33460_;
  assign new_n33462_ = ~new_n33455_ & ~new_n33461_;
  assign new_n33463_ = ~\b[18]  & ~new_n33462_;
  assign new_n33464_ = ~new_n33133_ & ~new_n33391_;
  assign new_n33465_ = ~new_n33143_ & new_n33343_;
  assign new_n33466_ = ~new_n33339_ & new_n33465_;
  assign new_n33467_ = ~new_n33340_ & ~new_n33343_;
  assign new_n33468_ = ~new_n33466_ & ~new_n33467_;
  assign new_n33469_ = new_n5172_ & ~new_n33468_;
  assign new_n33470_ = ~new_n33390_ & new_n33469_;
  assign new_n33471_ = ~new_n33464_ & ~new_n33470_;
  assign new_n33472_ = ~\b[17]  & ~new_n33471_;
  assign new_n33473_ = ~new_n33142_ & ~new_n33391_;
  assign new_n33474_ = ~new_n33152_ & new_n33338_;
  assign new_n33475_ = ~new_n33334_ & new_n33474_;
  assign new_n33476_ = ~new_n33335_ & ~new_n33338_;
  assign new_n33477_ = ~new_n33475_ & ~new_n33476_;
  assign new_n33478_ = new_n5172_ & ~new_n33477_;
  assign new_n33479_ = ~new_n33390_ & new_n33478_;
  assign new_n33480_ = ~new_n33473_ & ~new_n33479_;
  assign new_n33481_ = ~\b[16]  & ~new_n33480_;
  assign new_n33482_ = ~new_n33151_ & ~new_n33391_;
  assign new_n33483_ = ~new_n33161_ & new_n33333_;
  assign new_n33484_ = ~new_n33329_ & new_n33483_;
  assign new_n33485_ = ~new_n33330_ & ~new_n33333_;
  assign new_n33486_ = ~new_n33484_ & ~new_n33485_;
  assign new_n33487_ = new_n5172_ & ~new_n33486_;
  assign new_n33488_ = ~new_n33390_ & new_n33487_;
  assign new_n33489_ = ~new_n33482_ & ~new_n33488_;
  assign new_n33490_ = ~\b[15]  & ~new_n33489_;
  assign new_n33491_ = ~new_n33160_ & ~new_n33391_;
  assign new_n33492_ = ~new_n33170_ & new_n33328_;
  assign new_n33493_ = ~new_n33324_ & new_n33492_;
  assign new_n33494_ = ~new_n33325_ & ~new_n33328_;
  assign new_n33495_ = ~new_n33493_ & ~new_n33494_;
  assign new_n33496_ = new_n5172_ & ~new_n33495_;
  assign new_n33497_ = ~new_n33390_ & new_n33496_;
  assign new_n33498_ = ~new_n33491_ & ~new_n33497_;
  assign new_n33499_ = ~\b[14]  & ~new_n33498_;
  assign new_n33500_ = ~new_n33169_ & ~new_n33391_;
  assign new_n33501_ = ~new_n33179_ & new_n33323_;
  assign new_n33502_ = ~new_n33319_ & new_n33501_;
  assign new_n33503_ = ~new_n33320_ & ~new_n33323_;
  assign new_n33504_ = ~new_n33502_ & ~new_n33503_;
  assign new_n33505_ = new_n5172_ & ~new_n33504_;
  assign new_n33506_ = ~new_n33390_ & new_n33505_;
  assign new_n33507_ = ~new_n33500_ & ~new_n33506_;
  assign new_n33508_ = ~\b[13]  & ~new_n33507_;
  assign new_n33509_ = ~new_n33178_ & ~new_n33391_;
  assign new_n33510_ = ~new_n33188_ & new_n33318_;
  assign new_n33511_ = ~new_n33314_ & new_n33510_;
  assign new_n33512_ = ~new_n33315_ & ~new_n33318_;
  assign new_n33513_ = ~new_n33511_ & ~new_n33512_;
  assign new_n33514_ = new_n5172_ & ~new_n33513_;
  assign new_n33515_ = ~new_n33390_ & new_n33514_;
  assign new_n33516_ = ~new_n33509_ & ~new_n33515_;
  assign new_n33517_ = ~\b[12]  & ~new_n33516_;
  assign new_n33518_ = ~new_n33187_ & ~new_n33391_;
  assign new_n33519_ = ~new_n33197_ & new_n33313_;
  assign new_n33520_ = ~new_n33309_ & new_n33519_;
  assign new_n33521_ = ~new_n33310_ & ~new_n33313_;
  assign new_n33522_ = ~new_n33520_ & ~new_n33521_;
  assign new_n33523_ = new_n5172_ & ~new_n33522_;
  assign new_n33524_ = ~new_n33390_ & new_n33523_;
  assign new_n33525_ = ~new_n33518_ & ~new_n33524_;
  assign new_n33526_ = ~\b[11]  & ~new_n33525_;
  assign new_n33527_ = ~new_n33196_ & ~new_n33391_;
  assign new_n33528_ = ~new_n33206_ & new_n33308_;
  assign new_n33529_ = ~new_n33304_ & new_n33528_;
  assign new_n33530_ = ~new_n33305_ & ~new_n33308_;
  assign new_n33531_ = ~new_n33529_ & ~new_n33530_;
  assign new_n33532_ = new_n5172_ & ~new_n33531_;
  assign new_n33533_ = ~new_n33390_ & new_n33532_;
  assign new_n33534_ = ~new_n33527_ & ~new_n33533_;
  assign new_n33535_ = ~\b[10]  & ~new_n33534_;
  assign new_n33536_ = ~new_n33205_ & ~new_n33391_;
  assign new_n33537_ = ~new_n33215_ & new_n33303_;
  assign new_n33538_ = ~new_n33299_ & new_n33537_;
  assign new_n33539_ = ~new_n33300_ & ~new_n33303_;
  assign new_n33540_ = ~new_n33538_ & ~new_n33539_;
  assign new_n33541_ = new_n5172_ & ~new_n33540_;
  assign new_n33542_ = ~new_n33390_ & new_n33541_;
  assign new_n33543_ = ~new_n33536_ & ~new_n33542_;
  assign new_n33544_ = ~\b[9]  & ~new_n33543_;
  assign new_n33545_ = ~new_n33214_ & ~new_n33391_;
  assign new_n33546_ = ~new_n33224_ & new_n33298_;
  assign new_n33547_ = ~new_n33294_ & new_n33546_;
  assign new_n33548_ = ~new_n33295_ & ~new_n33298_;
  assign new_n33549_ = ~new_n33547_ & ~new_n33548_;
  assign new_n33550_ = new_n5172_ & ~new_n33549_;
  assign new_n33551_ = ~new_n33390_ & new_n33550_;
  assign new_n33552_ = ~new_n33545_ & ~new_n33551_;
  assign new_n33553_ = ~\b[8]  & ~new_n33552_;
  assign new_n33554_ = ~new_n33223_ & ~new_n33391_;
  assign new_n33555_ = ~new_n33233_ & new_n33293_;
  assign new_n33556_ = ~new_n33289_ & new_n33555_;
  assign new_n33557_ = ~new_n33290_ & ~new_n33293_;
  assign new_n33558_ = ~new_n33556_ & ~new_n33557_;
  assign new_n33559_ = new_n5172_ & ~new_n33558_;
  assign new_n33560_ = ~new_n33390_ & new_n33559_;
  assign new_n33561_ = ~new_n33554_ & ~new_n33560_;
  assign new_n33562_ = ~\b[7]  & ~new_n33561_;
  assign new_n33563_ = ~new_n33232_ & ~new_n33391_;
  assign new_n33564_ = ~new_n33242_ & new_n33288_;
  assign new_n33565_ = ~new_n33284_ & new_n33564_;
  assign new_n33566_ = ~new_n33285_ & ~new_n33288_;
  assign new_n33567_ = ~new_n33565_ & ~new_n33566_;
  assign new_n33568_ = new_n5172_ & ~new_n33567_;
  assign new_n33569_ = ~new_n33390_ & new_n33568_;
  assign new_n33570_ = ~new_n33563_ & ~new_n33569_;
  assign new_n33571_ = ~\b[6]  & ~new_n33570_;
  assign new_n33572_ = ~new_n33241_ & ~new_n33391_;
  assign new_n33573_ = ~new_n33251_ & new_n33283_;
  assign new_n33574_ = ~new_n33279_ & new_n33573_;
  assign new_n33575_ = ~new_n33280_ & ~new_n33283_;
  assign new_n33576_ = ~new_n33574_ & ~new_n33575_;
  assign new_n33577_ = new_n5172_ & ~new_n33576_;
  assign new_n33578_ = ~new_n33390_ & new_n33577_;
  assign new_n33579_ = ~new_n33572_ & ~new_n33578_;
  assign new_n33580_ = ~\b[5]  & ~new_n33579_;
  assign new_n33581_ = ~new_n33250_ & ~new_n33391_;
  assign new_n33582_ = ~new_n33259_ & new_n33278_;
  assign new_n33583_ = ~new_n33274_ & new_n33582_;
  assign new_n33584_ = ~new_n33275_ & ~new_n33278_;
  assign new_n33585_ = ~new_n33583_ & ~new_n33584_;
  assign new_n33586_ = new_n5172_ & ~new_n33585_;
  assign new_n33587_ = ~new_n33390_ & new_n33586_;
  assign new_n33588_ = ~new_n33581_ & ~new_n33587_;
  assign new_n33589_ = ~\b[4]  & ~new_n33588_;
  assign new_n33590_ = ~new_n33258_ & ~new_n33391_;
  assign new_n33591_ = ~new_n33269_ & new_n33273_;
  assign new_n33592_ = ~new_n33268_ & new_n33591_;
  assign new_n33593_ = ~new_n33270_ & ~new_n33273_;
  assign new_n33594_ = ~new_n33592_ & ~new_n33593_;
  assign new_n33595_ = new_n5172_ & ~new_n33594_;
  assign new_n33596_ = ~new_n33390_ & new_n33595_;
  assign new_n33597_ = ~new_n33590_ & ~new_n33596_;
  assign new_n33598_ = ~\b[3]  & ~new_n33597_;
  assign new_n33599_ = ~new_n33263_ & ~new_n33391_;
  assign new_n33600_ = new_n5046_ & ~new_n33266_;
  assign new_n33601_ = ~new_n33264_ & new_n33600_;
  assign new_n33602_ = new_n5172_ & ~new_n33601_;
  assign new_n33603_ = ~new_n33268_ & new_n33602_;
  assign new_n33604_ = ~new_n33390_ & new_n33603_;
  assign new_n33605_ = ~new_n33599_ & ~new_n33604_;
  assign new_n33606_ = ~\b[2]  & ~new_n33605_;
  assign new_n33607_ = new_n5393_ & ~new_n33390_;
  assign new_n33608_ = \a[38]  & ~new_n33607_;
  assign new_n33609_ = new_n5399_ & ~new_n33390_;
  assign new_n33610_ = ~new_n33608_ & ~new_n33609_;
  assign new_n33611_ = \b[1]  & ~new_n33610_;
  assign new_n33612_ = ~\b[1]  & ~new_n33609_;
  assign new_n33613_ = ~new_n33608_ & new_n33612_;
  assign new_n33614_ = ~new_n33611_ & ~new_n33613_;
  assign new_n33615_ = ~new_n5406_ & ~new_n33614_;
  assign new_n33616_ = ~\b[1]  & ~new_n33610_;
  assign new_n33617_ = ~new_n33615_ & ~new_n33616_;
  assign new_n33618_ = \b[2]  & ~new_n33604_;
  assign new_n33619_ = ~new_n33599_ & new_n33618_;
  assign new_n33620_ = ~new_n33606_ & ~new_n33619_;
  assign new_n33621_ = ~new_n33617_ & new_n33620_;
  assign new_n33622_ = ~new_n33606_ & ~new_n33621_;
  assign new_n33623_ = \b[3]  & ~new_n33596_;
  assign new_n33624_ = ~new_n33590_ & new_n33623_;
  assign new_n33625_ = ~new_n33598_ & ~new_n33624_;
  assign new_n33626_ = ~new_n33622_ & new_n33625_;
  assign new_n33627_ = ~new_n33598_ & ~new_n33626_;
  assign new_n33628_ = \b[4]  & ~new_n33587_;
  assign new_n33629_ = ~new_n33581_ & new_n33628_;
  assign new_n33630_ = ~new_n33589_ & ~new_n33629_;
  assign new_n33631_ = ~new_n33627_ & new_n33630_;
  assign new_n33632_ = ~new_n33589_ & ~new_n33631_;
  assign new_n33633_ = \b[5]  & ~new_n33578_;
  assign new_n33634_ = ~new_n33572_ & new_n33633_;
  assign new_n33635_ = ~new_n33580_ & ~new_n33634_;
  assign new_n33636_ = ~new_n33632_ & new_n33635_;
  assign new_n33637_ = ~new_n33580_ & ~new_n33636_;
  assign new_n33638_ = \b[6]  & ~new_n33569_;
  assign new_n33639_ = ~new_n33563_ & new_n33638_;
  assign new_n33640_ = ~new_n33571_ & ~new_n33639_;
  assign new_n33641_ = ~new_n33637_ & new_n33640_;
  assign new_n33642_ = ~new_n33571_ & ~new_n33641_;
  assign new_n33643_ = \b[7]  & ~new_n33560_;
  assign new_n33644_ = ~new_n33554_ & new_n33643_;
  assign new_n33645_ = ~new_n33562_ & ~new_n33644_;
  assign new_n33646_ = ~new_n33642_ & new_n33645_;
  assign new_n33647_ = ~new_n33562_ & ~new_n33646_;
  assign new_n33648_ = \b[8]  & ~new_n33551_;
  assign new_n33649_ = ~new_n33545_ & new_n33648_;
  assign new_n33650_ = ~new_n33553_ & ~new_n33649_;
  assign new_n33651_ = ~new_n33647_ & new_n33650_;
  assign new_n33652_ = ~new_n33553_ & ~new_n33651_;
  assign new_n33653_ = \b[9]  & ~new_n33542_;
  assign new_n33654_ = ~new_n33536_ & new_n33653_;
  assign new_n33655_ = ~new_n33544_ & ~new_n33654_;
  assign new_n33656_ = ~new_n33652_ & new_n33655_;
  assign new_n33657_ = ~new_n33544_ & ~new_n33656_;
  assign new_n33658_ = \b[10]  & ~new_n33533_;
  assign new_n33659_ = ~new_n33527_ & new_n33658_;
  assign new_n33660_ = ~new_n33535_ & ~new_n33659_;
  assign new_n33661_ = ~new_n33657_ & new_n33660_;
  assign new_n33662_ = ~new_n33535_ & ~new_n33661_;
  assign new_n33663_ = \b[11]  & ~new_n33524_;
  assign new_n33664_ = ~new_n33518_ & new_n33663_;
  assign new_n33665_ = ~new_n33526_ & ~new_n33664_;
  assign new_n33666_ = ~new_n33662_ & new_n33665_;
  assign new_n33667_ = ~new_n33526_ & ~new_n33666_;
  assign new_n33668_ = \b[12]  & ~new_n33515_;
  assign new_n33669_ = ~new_n33509_ & new_n33668_;
  assign new_n33670_ = ~new_n33517_ & ~new_n33669_;
  assign new_n33671_ = ~new_n33667_ & new_n33670_;
  assign new_n33672_ = ~new_n33517_ & ~new_n33671_;
  assign new_n33673_ = \b[13]  & ~new_n33506_;
  assign new_n33674_ = ~new_n33500_ & new_n33673_;
  assign new_n33675_ = ~new_n33508_ & ~new_n33674_;
  assign new_n33676_ = ~new_n33672_ & new_n33675_;
  assign new_n33677_ = ~new_n33508_ & ~new_n33676_;
  assign new_n33678_ = \b[14]  & ~new_n33497_;
  assign new_n33679_ = ~new_n33491_ & new_n33678_;
  assign new_n33680_ = ~new_n33499_ & ~new_n33679_;
  assign new_n33681_ = ~new_n33677_ & new_n33680_;
  assign new_n33682_ = ~new_n33499_ & ~new_n33681_;
  assign new_n33683_ = \b[15]  & ~new_n33488_;
  assign new_n33684_ = ~new_n33482_ & new_n33683_;
  assign new_n33685_ = ~new_n33490_ & ~new_n33684_;
  assign new_n33686_ = ~new_n33682_ & new_n33685_;
  assign new_n33687_ = ~new_n33490_ & ~new_n33686_;
  assign new_n33688_ = \b[16]  & ~new_n33479_;
  assign new_n33689_ = ~new_n33473_ & new_n33688_;
  assign new_n33690_ = ~new_n33481_ & ~new_n33689_;
  assign new_n33691_ = ~new_n33687_ & new_n33690_;
  assign new_n33692_ = ~new_n33481_ & ~new_n33691_;
  assign new_n33693_ = \b[17]  & ~new_n33470_;
  assign new_n33694_ = ~new_n33464_ & new_n33693_;
  assign new_n33695_ = ~new_n33472_ & ~new_n33694_;
  assign new_n33696_ = ~new_n33692_ & new_n33695_;
  assign new_n33697_ = ~new_n33472_ & ~new_n33696_;
  assign new_n33698_ = \b[18]  & ~new_n33461_;
  assign new_n33699_ = ~new_n33455_ & new_n33698_;
  assign new_n33700_ = ~new_n33463_ & ~new_n33699_;
  assign new_n33701_ = ~new_n33697_ & new_n33700_;
  assign new_n33702_ = ~new_n33463_ & ~new_n33701_;
  assign new_n33703_ = \b[19]  & ~new_n33452_;
  assign new_n33704_ = ~new_n33446_ & new_n33703_;
  assign new_n33705_ = ~new_n33454_ & ~new_n33704_;
  assign new_n33706_ = ~new_n33702_ & new_n33705_;
  assign new_n33707_ = ~new_n33454_ & ~new_n33706_;
  assign new_n33708_ = \b[20]  & ~new_n33443_;
  assign new_n33709_ = ~new_n33437_ & new_n33708_;
  assign new_n33710_ = ~new_n33445_ & ~new_n33709_;
  assign new_n33711_ = ~new_n33707_ & new_n33710_;
  assign new_n33712_ = ~new_n33445_ & ~new_n33711_;
  assign new_n33713_ = \b[21]  & ~new_n33434_;
  assign new_n33714_ = ~new_n33428_ & new_n33713_;
  assign new_n33715_ = ~new_n33436_ & ~new_n33714_;
  assign new_n33716_ = ~new_n33712_ & new_n33715_;
  assign new_n33717_ = ~new_n33436_ & ~new_n33716_;
  assign new_n33718_ = \b[22]  & ~new_n33425_;
  assign new_n33719_ = ~new_n33419_ & new_n33718_;
  assign new_n33720_ = ~new_n33427_ & ~new_n33719_;
  assign new_n33721_ = ~new_n33717_ & new_n33720_;
  assign new_n33722_ = ~new_n33427_ & ~new_n33721_;
  assign new_n33723_ = \b[23]  & ~new_n33416_;
  assign new_n33724_ = ~new_n33410_ & new_n33723_;
  assign new_n33725_ = ~new_n33418_ & ~new_n33724_;
  assign new_n33726_ = ~new_n33722_ & new_n33725_;
  assign new_n33727_ = ~new_n33418_ & ~new_n33726_;
  assign new_n33728_ = \b[24]  & ~new_n33407_;
  assign new_n33729_ = ~new_n33401_ & new_n33728_;
  assign new_n33730_ = ~new_n33409_ & ~new_n33729_;
  assign new_n33731_ = ~new_n33727_ & new_n33730_;
  assign new_n33732_ = ~new_n33409_ & ~new_n33731_;
  assign new_n33733_ = \b[25]  & ~new_n33398_;
  assign new_n33734_ = ~new_n33392_ & new_n33733_;
  assign new_n33735_ = ~new_n33400_ & ~new_n33734_;
  assign new_n33736_ = ~new_n33732_ & new_n33735_;
  assign new_n33737_ = ~new_n33400_ & ~new_n33736_;
  assign new_n33738_ = ~new_n33060_ & ~new_n33391_;
  assign new_n33739_ = ~new_n33062_ & new_n33388_;
  assign new_n33740_ = ~new_n33384_ & new_n33739_;
  assign new_n33741_ = ~new_n33385_ & ~new_n33388_;
  assign new_n33742_ = ~new_n33740_ & ~new_n33741_;
  assign new_n33743_ = new_n33391_ & ~new_n33742_;
  assign new_n33744_ = ~new_n33738_ & ~new_n33743_;
  assign new_n33745_ = ~\b[26]  & ~new_n33744_;
  assign new_n33746_ = \b[26]  & ~new_n33738_;
  assign new_n33747_ = ~new_n33743_ & new_n33746_;
  assign new_n33748_ = new_n5542_ & ~new_n33747_;
  assign new_n33749_ = ~new_n33745_ & new_n33748_;
  assign new_n33750_ = ~new_n33737_ & new_n33749_;
  assign new_n33751_ = new_n5172_ & ~new_n33744_;
  assign new_n33752_ = ~new_n33750_ & ~new_n33751_;
  assign new_n33753_ = ~new_n33409_ & new_n33735_;
  assign new_n33754_ = ~new_n33731_ & new_n33753_;
  assign new_n33755_ = ~new_n33732_ & ~new_n33735_;
  assign new_n33756_ = ~new_n33754_ & ~new_n33755_;
  assign new_n33757_ = ~new_n33752_ & ~new_n33756_;
  assign new_n33758_ = ~new_n33399_ & ~new_n33751_;
  assign new_n33759_ = ~new_n33750_ & new_n33758_;
  assign new_n33760_ = ~new_n33757_ & ~new_n33759_;
  assign new_n33761_ = ~new_n33400_ & ~new_n33747_;
  assign new_n33762_ = ~new_n33745_ & new_n33761_;
  assign new_n33763_ = ~new_n33736_ & new_n33762_;
  assign new_n33764_ = ~new_n33745_ & ~new_n33747_;
  assign new_n33765_ = ~new_n33737_ & ~new_n33764_;
  assign new_n33766_ = ~new_n33763_ & ~new_n33765_;
  assign new_n33767_ = ~new_n33752_ & ~new_n33766_;
  assign new_n33768_ = ~new_n33744_ & ~new_n33751_;
  assign new_n33769_ = ~new_n33750_ & new_n33768_;
  assign new_n33770_ = ~new_n33767_ & ~new_n33769_;
  assign new_n33771_ = ~\b[27]  & ~new_n33770_;
  assign new_n33772_ = ~\b[26]  & ~new_n33760_;
  assign new_n33773_ = ~new_n33418_ & new_n33730_;
  assign new_n33774_ = ~new_n33726_ & new_n33773_;
  assign new_n33775_ = ~new_n33727_ & ~new_n33730_;
  assign new_n33776_ = ~new_n33774_ & ~new_n33775_;
  assign new_n33777_ = ~new_n33752_ & ~new_n33776_;
  assign new_n33778_ = ~new_n33408_ & ~new_n33751_;
  assign new_n33779_ = ~new_n33750_ & new_n33778_;
  assign new_n33780_ = ~new_n33777_ & ~new_n33779_;
  assign new_n33781_ = ~\b[25]  & ~new_n33780_;
  assign new_n33782_ = ~new_n33427_ & new_n33725_;
  assign new_n33783_ = ~new_n33721_ & new_n33782_;
  assign new_n33784_ = ~new_n33722_ & ~new_n33725_;
  assign new_n33785_ = ~new_n33783_ & ~new_n33784_;
  assign new_n33786_ = ~new_n33752_ & ~new_n33785_;
  assign new_n33787_ = ~new_n33417_ & ~new_n33751_;
  assign new_n33788_ = ~new_n33750_ & new_n33787_;
  assign new_n33789_ = ~new_n33786_ & ~new_n33788_;
  assign new_n33790_ = ~\b[24]  & ~new_n33789_;
  assign new_n33791_ = ~new_n33436_ & new_n33720_;
  assign new_n33792_ = ~new_n33716_ & new_n33791_;
  assign new_n33793_ = ~new_n33717_ & ~new_n33720_;
  assign new_n33794_ = ~new_n33792_ & ~new_n33793_;
  assign new_n33795_ = ~new_n33752_ & ~new_n33794_;
  assign new_n33796_ = ~new_n33426_ & ~new_n33751_;
  assign new_n33797_ = ~new_n33750_ & new_n33796_;
  assign new_n33798_ = ~new_n33795_ & ~new_n33797_;
  assign new_n33799_ = ~\b[23]  & ~new_n33798_;
  assign new_n33800_ = ~new_n33445_ & new_n33715_;
  assign new_n33801_ = ~new_n33711_ & new_n33800_;
  assign new_n33802_ = ~new_n33712_ & ~new_n33715_;
  assign new_n33803_ = ~new_n33801_ & ~new_n33802_;
  assign new_n33804_ = ~new_n33752_ & ~new_n33803_;
  assign new_n33805_ = ~new_n33435_ & ~new_n33751_;
  assign new_n33806_ = ~new_n33750_ & new_n33805_;
  assign new_n33807_ = ~new_n33804_ & ~new_n33806_;
  assign new_n33808_ = ~\b[22]  & ~new_n33807_;
  assign new_n33809_ = ~new_n33454_ & new_n33710_;
  assign new_n33810_ = ~new_n33706_ & new_n33809_;
  assign new_n33811_ = ~new_n33707_ & ~new_n33710_;
  assign new_n33812_ = ~new_n33810_ & ~new_n33811_;
  assign new_n33813_ = ~new_n33752_ & ~new_n33812_;
  assign new_n33814_ = ~new_n33444_ & ~new_n33751_;
  assign new_n33815_ = ~new_n33750_ & new_n33814_;
  assign new_n33816_ = ~new_n33813_ & ~new_n33815_;
  assign new_n33817_ = ~\b[21]  & ~new_n33816_;
  assign new_n33818_ = ~new_n33463_ & new_n33705_;
  assign new_n33819_ = ~new_n33701_ & new_n33818_;
  assign new_n33820_ = ~new_n33702_ & ~new_n33705_;
  assign new_n33821_ = ~new_n33819_ & ~new_n33820_;
  assign new_n33822_ = ~new_n33752_ & ~new_n33821_;
  assign new_n33823_ = ~new_n33453_ & ~new_n33751_;
  assign new_n33824_ = ~new_n33750_ & new_n33823_;
  assign new_n33825_ = ~new_n33822_ & ~new_n33824_;
  assign new_n33826_ = ~\b[20]  & ~new_n33825_;
  assign new_n33827_ = ~new_n33472_ & new_n33700_;
  assign new_n33828_ = ~new_n33696_ & new_n33827_;
  assign new_n33829_ = ~new_n33697_ & ~new_n33700_;
  assign new_n33830_ = ~new_n33828_ & ~new_n33829_;
  assign new_n33831_ = ~new_n33752_ & ~new_n33830_;
  assign new_n33832_ = ~new_n33462_ & ~new_n33751_;
  assign new_n33833_ = ~new_n33750_ & new_n33832_;
  assign new_n33834_ = ~new_n33831_ & ~new_n33833_;
  assign new_n33835_ = ~\b[19]  & ~new_n33834_;
  assign new_n33836_ = ~new_n33481_ & new_n33695_;
  assign new_n33837_ = ~new_n33691_ & new_n33836_;
  assign new_n33838_ = ~new_n33692_ & ~new_n33695_;
  assign new_n33839_ = ~new_n33837_ & ~new_n33838_;
  assign new_n33840_ = ~new_n33752_ & ~new_n33839_;
  assign new_n33841_ = ~new_n33471_ & ~new_n33751_;
  assign new_n33842_ = ~new_n33750_ & new_n33841_;
  assign new_n33843_ = ~new_n33840_ & ~new_n33842_;
  assign new_n33844_ = ~\b[18]  & ~new_n33843_;
  assign new_n33845_ = ~new_n33490_ & new_n33690_;
  assign new_n33846_ = ~new_n33686_ & new_n33845_;
  assign new_n33847_ = ~new_n33687_ & ~new_n33690_;
  assign new_n33848_ = ~new_n33846_ & ~new_n33847_;
  assign new_n33849_ = ~new_n33752_ & ~new_n33848_;
  assign new_n33850_ = ~new_n33480_ & ~new_n33751_;
  assign new_n33851_ = ~new_n33750_ & new_n33850_;
  assign new_n33852_ = ~new_n33849_ & ~new_n33851_;
  assign new_n33853_ = ~\b[17]  & ~new_n33852_;
  assign new_n33854_ = ~new_n33499_ & new_n33685_;
  assign new_n33855_ = ~new_n33681_ & new_n33854_;
  assign new_n33856_ = ~new_n33682_ & ~new_n33685_;
  assign new_n33857_ = ~new_n33855_ & ~new_n33856_;
  assign new_n33858_ = ~new_n33752_ & ~new_n33857_;
  assign new_n33859_ = ~new_n33489_ & ~new_n33751_;
  assign new_n33860_ = ~new_n33750_ & new_n33859_;
  assign new_n33861_ = ~new_n33858_ & ~new_n33860_;
  assign new_n33862_ = ~\b[16]  & ~new_n33861_;
  assign new_n33863_ = ~new_n33508_ & new_n33680_;
  assign new_n33864_ = ~new_n33676_ & new_n33863_;
  assign new_n33865_ = ~new_n33677_ & ~new_n33680_;
  assign new_n33866_ = ~new_n33864_ & ~new_n33865_;
  assign new_n33867_ = ~new_n33752_ & ~new_n33866_;
  assign new_n33868_ = ~new_n33498_ & ~new_n33751_;
  assign new_n33869_ = ~new_n33750_ & new_n33868_;
  assign new_n33870_ = ~new_n33867_ & ~new_n33869_;
  assign new_n33871_ = ~\b[15]  & ~new_n33870_;
  assign new_n33872_ = ~new_n33517_ & new_n33675_;
  assign new_n33873_ = ~new_n33671_ & new_n33872_;
  assign new_n33874_ = ~new_n33672_ & ~new_n33675_;
  assign new_n33875_ = ~new_n33873_ & ~new_n33874_;
  assign new_n33876_ = ~new_n33752_ & ~new_n33875_;
  assign new_n33877_ = ~new_n33507_ & ~new_n33751_;
  assign new_n33878_ = ~new_n33750_ & new_n33877_;
  assign new_n33879_ = ~new_n33876_ & ~new_n33878_;
  assign new_n33880_ = ~\b[14]  & ~new_n33879_;
  assign new_n33881_ = ~new_n33526_ & new_n33670_;
  assign new_n33882_ = ~new_n33666_ & new_n33881_;
  assign new_n33883_ = ~new_n33667_ & ~new_n33670_;
  assign new_n33884_ = ~new_n33882_ & ~new_n33883_;
  assign new_n33885_ = ~new_n33752_ & ~new_n33884_;
  assign new_n33886_ = ~new_n33516_ & ~new_n33751_;
  assign new_n33887_ = ~new_n33750_ & new_n33886_;
  assign new_n33888_ = ~new_n33885_ & ~new_n33887_;
  assign new_n33889_ = ~\b[13]  & ~new_n33888_;
  assign new_n33890_ = ~new_n33535_ & new_n33665_;
  assign new_n33891_ = ~new_n33661_ & new_n33890_;
  assign new_n33892_ = ~new_n33662_ & ~new_n33665_;
  assign new_n33893_ = ~new_n33891_ & ~new_n33892_;
  assign new_n33894_ = ~new_n33752_ & ~new_n33893_;
  assign new_n33895_ = ~new_n33525_ & ~new_n33751_;
  assign new_n33896_ = ~new_n33750_ & new_n33895_;
  assign new_n33897_ = ~new_n33894_ & ~new_n33896_;
  assign new_n33898_ = ~\b[12]  & ~new_n33897_;
  assign new_n33899_ = ~new_n33544_ & new_n33660_;
  assign new_n33900_ = ~new_n33656_ & new_n33899_;
  assign new_n33901_ = ~new_n33657_ & ~new_n33660_;
  assign new_n33902_ = ~new_n33900_ & ~new_n33901_;
  assign new_n33903_ = ~new_n33752_ & ~new_n33902_;
  assign new_n33904_ = ~new_n33534_ & ~new_n33751_;
  assign new_n33905_ = ~new_n33750_ & new_n33904_;
  assign new_n33906_ = ~new_n33903_ & ~new_n33905_;
  assign new_n33907_ = ~\b[11]  & ~new_n33906_;
  assign new_n33908_ = ~new_n33553_ & new_n33655_;
  assign new_n33909_ = ~new_n33651_ & new_n33908_;
  assign new_n33910_ = ~new_n33652_ & ~new_n33655_;
  assign new_n33911_ = ~new_n33909_ & ~new_n33910_;
  assign new_n33912_ = ~new_n33752_ & ~new_n33911_;
  assign new_n33913_ = ~new_n33543_ & ~new_n33751_;
  assign new_n33914_ = ~new_n33750_ & new_n33913_;
  assign new_n33915_ = ~new_n33912_ & ~new_n33914_;
  assign new_n33916_ = ~\b[10]  & ~new_n33915_;
  assign new_n33917_ = ~new_n33562_ & new_n33650_;
  assign new_n33918_ = ~new_n33646_ & new_n33917_;
  assign new_n33919_ = ~new_n33647_ & ~new_n33650_;
  assign new_n33920_ = ~new_n33918_ & ~new_n33919_;
  assign new_n33921_ = ~new_n33752_ & ~new_n33920_;
  assign new_n33922_ = ~new_n33552_ & ~new_n33751_;
  assign new_n33923_ = ~new_n33750_ & new_n33922_;
  assign new_n33924_ = ~new_n33921_ & ~new_n33923_;
  assign new_n33925_ = ~\b[9]  & ~new_n33924_;
  assign new_n33926_ = ~new_n33571_ & new_n33645_;
  assign new_n33927_ = ~new_n33641_ & new_n33926_;
  assign new_n33928_ = ~new_n33642_ & ~new_n33645_;
  assign new_n33929_ = ~new_n33927_ & ~new_n33928_;
  assign new_n33930_ = ~new_n33752_ & ~new_n33929_;
  assign new_n33931_ = ~new_n33561_ & ~new_n33751_;
  assign new_n33932_ = ~new_n33750_ & new_n33931_;
  assign new_n33933_ = ~new_n33930_ & ~new_n33932_;
  assign new_n33934_ = ~\b[8]  & ~new_n33933_;
  assign new_n33935_ = ~new_n33580_ & new_n33640_;
  assign new_n33936_ = ~new_n33636_ & new_n33935_;
  assign new_n33937_ = ~new_n33637_ & ~new_n33640_;
  assign new_n33938_ = ~new_n33936_ & ~new_n33937_;
  assign new_n33939_ = ~new_n33752_ & ~new_n33938_;
  assign new_n33940_ = ~new_n33570_ & ~new_n33751_;
  assign new_n33941_ = ~new_n33750_ & new_n33940_;
  assign new_n33942_ = ~new_n33939_ & ~new_n33941_;
  assign new_n33943_ = ~\b[7]  & ~new_n33942_;
  assign new_n33944_ = ~new_n33589_ & new_n33635_;
  assign new_n33945_ = ~new_n33631_ & new_n33944_;
  assign new_n33946_ = ~new_n33632_ & ~new_n33635_;
  assign new_n33947_ = ~new_n33945_ & ~new_n33946_;
  assign new_n33948_ = ~new_n33752_ & ~new_n33947_;
  assign new_n33949_ = ~new_n33579_ & ~new_n33751_;
  assign new_n33950_ = ~new_n33750_ & new_n33949_;
  assign new_n33951_ = ~new_n33948_ & ~new_n33950_;
  assign new_n33952_ = ~\b[6]  & ~new_n33951_;
  assign new_n33953_ = ~new_n33598_ & new_n33630_;
  assign new_n33954_ = ~new_n33626_ & new_n33953_;
  assign new_n33955_ = ~new_n33627_ & ~new_n33630_;
  assign new_n33956_ = ~new_n33954_ & ~new_n33955_;
  assign new_n33957_ = ~new_n33752_ & ~new_n33956_;
  assign new_n33958_ = ~new_n33588_ & ~new_n33751_;
  assign new_n33959_ = ~new_n33750_ & new_n33958_;
  assign new_n33960_ = ~new_n33957_ & ~new_n33959_;
  assign new_n33961_ = ~\b[5]  & ~new_n33960_;
  assign new_n33962_ = ~new_n33606_ & new_n33625_;
  assign new_n33963_ = ~new_n33621_ & new_n33962_;
  assign new_n33964_ = ~new_n33622_ & ~new_n33625_;
  assign new_n33965_ = ~new_n33963_ & ~new_n33964_;
  assign new_n33966_ = ~new_n33752_ & ~new_n33965_;
  assign new_n33967_ = ~new_n33597_ & ~new_n33751_;
  assign new_n33968_ = ~new_n33750_ & new_n33967_;
  assign new_n33969_ = ~new_n33966_ & ~new_n33968_;
  assign new_n33970_ = ~\b[4]  & ~new_n33969_;
  assign new_n33971_ = ~new_n33616_ & new_n33620_;
  assign new_n33972_ = ~new_n33615_ & new_n33971_;
  assign new_n33973_ = ~new_n33617_ & ~new_n33620_;
  assign new_n33974_ = ~new_n33972_ & ~new_n33973_;
  assign new_n33975_ = ~new_n33752_ & ~new_n33974_;
  assign new_n33976_ = ~new_n33605_ & ~new_n33751_;
  assign new_n33977_ = ~new_n33750_ & new_n33976_;
  assign new_n33978_ = ~new_n33975_ & ~new_n33977_;
  assign new_n33979_ = ~\b[3]  & ~new_n33978_;
  assign new_n33980_ = new_n5406_ & ~new_n33613_;
  assign new_n33981_ = ~new_n33611_ & new_n33980_;
  assign new_n33982_ = ~new_n33615_ & ~new_n33981_;
  assign new_n33983_ = ~new_n33752_ & new_n33982_;
  assign new_n33984_ = ~new_n33610_ & ~new_n33751_;
  assign new_n33985_ = ~new_n33750_ & new_n33984_;
  assign new_n33986_ = ~new_n33983_ & ~new_n33985_;
  assign new_n33987_ = ~\b[2]  & ~new_n33986_;
  assign new_n33988_ = \b[0]  & ~new_n33752_;
  assign new_n33989_ = \a[37]  & ~new_n33988_;
  assign new_n33990_ = new_n5406_ & ~new_n33752_;
  assign new_n33991_ = ~new_n33989_ & ~new_n33990_;
  assign new_n33992_ = \b[1]  & ~new_n33991_;
  assign new_n33993_ = ~\b[1]  & ~new_n33990_;
  assign new_n33994_ = ~new_n33989_ & new_n33993_;
  assign new_n33995_ = ~new_n33992_ & ~new_n33994_;
  assign new_n33996_ = ~new_n5791_ & ~new_n33995_;
  assign new_n33997_ = ~\b[1]  & ~new_n33991_;
  assign new_n33998_ = ~new_n33996_ & ~new_n33997_;
  assign new_n33999_ = \b[2]  & ~new_n33985_;
  assign new_n34000_ = ~new_n33983_ & new_n33999_;
  assign new_n34001_ = ~new_n33987_ & ~new_n34000_;
  assign new_n34002_ = ~new_n33998_ & new_n34001_;
  assign new_n34003_ = ~new_n33987_ & ~new_n34002_;
  assign new_n34004_ = \b[3]  & ~new_n33977_;
  assign new_n34005_ = ~new_n33975_ & new_n34004_;
  assign new_n34006_ = ~new_n33979_ & ~new_n34005_;
  assign new_n34007_ = ~new_n34003_ & new_n34006_;
  assign new_n34008_ = ~new_n33979_ & ~new_n34007_;
  assign new_n34009_ = \b[4]  & ~new_n33968_;
  assign new_n34010_ = ~new_n33966_ & new_n34009_;
  assign new_n34011_ = ~new_n33970_ & ~new_n34010_;
  assign new_n34012_ = ~new_n34008_ & new_n34011_;
  assign new_n34013_ = ~new_n33970_ & ~new_n34012_;
  assign new_n34014_ = \b[5]  & ~new_n33959_;
  assign new_n34015_ = ~new_n33957_ & new_n34014_;
  assign new_n34016_ = ~new_n33961_ & ~new_n34015_;
  assign new_n34017_ = ~new_n34013_ & new_n34016_;
  assign new_n34018_ = ~new_n33961_ & ~new_n34017_;
  assign new_n34019_ = \b[6]  & ~new_n33950_;
  assign new_n34020_ = ~new_n33948_ & new_n34019_;
  assign new_n34021_ = ~new_n33952_ & ~new_n34020_;
  assign new_n34022_ = ~new_n34018_ & new_n34021_;
  assign new_n34023_ = ~new_n33952_ & ~new_n34022_;
  assign new_n34024_ = \b[7]  & ~new_n33941_;
  assign new_n34025_ = ~new_n33939_ & new_n34024_;
  assign new_n34026_ = ~new_n33943_ & ~new_n34025_;
  assign new_n34027_ = ~new_n34023_ & new_n34026_;
  assign new_n34028_ = ~new_n33943_ & ~new_n34027_;
  assign new_n34029_ = \b[8]  & ~new_n33932_;
  assign new_n34030_ = ~new_n33930_ & new_n34029_;
  assign new_n34031_ = ~new_n33934_ & ~new_n34030_;
  assign new_n34032_ = ~new_n34028_ & new_n34031_;
  assign new_n34033_ = ~new_n33934_ & ~new_n34032_;
  assign new_n34034_ = \b[9]  & ~new_n33923_;
  assign new_n34035_ = ~new_n33921_ & new_n34034_;
  assign new_n34036_ = ~new_n33925_ & ~new_n34035_;
  assign new_n34037_ = ~new_n34033_ & new_n34036_;
  assign new_n34038_ = ~new_n33925_ & ~new_n34037_;
  assign new_n34039_ = \b[10]  & ~new_n33914_;
  assign new_n34040_ = ~new_n33912_ & new_n34039_;
  assign new_n34041_ = ~new_n33916_ & ~new_n34040_;
  assign new_n34042_ = ~new_n34038_ & new_n34041_;
  assign new_n34043_ = ~new_n33916_ & ~new_n34042_;
  assign new_n34044_ = \b[11]  & ~new_n33905_;
  assign new_n34045_ = ~new_n33903_ & new_n34044_;
  assign new_n34046_ = ~new_n33907_ & ~new_n34045_;
  assign new_n34047_ = ~new_n34043_ & new_n34046_;
  assign new_n34048_ = ~new_n33907_ & ~new_n34047_;
  assign new_n34049_ = \b[12]  & ~new_n33896_;
  assign new_n34050_ = ~new_n33894_ & new_n34049_;
  assign new_n34051_ = ~new_n33898_ & ~new_n34050_;
  assign new_n34052_ = ~new_n34048_ & new_n34051_;
  assign new_n34053_ = ~new_n33898_ & ~new_n34052_;
  assign new_n34054_ = \b[13]  & ~new_n33887_;
  assign new_n34055_ = ~new_n33885_ & new_n34054_;
  assign new_n34056_ = ~new_n33889_ & ~new_n34055_;
  assign new_n34057_ = ~new_n34053_ & new_n34056_;
  assign new_n34058_ = ~new_n33889_ & ~new_n34057_;
  assign new_n34059_ = \b[14]  & ~new_n33878_;
  assign new_n34060_ = ~new_n33876_ & new_n34059_;
  assign new_n34061_ = ~new_n33880_ & ~new_n34060_;
  assign new_n34062_ = ~new_n34058_ & new_n34061_;
  assign new_n34063_ = ~new_n33880_ & ~new_n34062_;
  assign new_n34064_ = \b[15]  & ~new_n33869_;
  assign new_n34065_ = ~new_n33867_ & new_n34064_;
  assign new_n34066_ = ~new_n33871_ & ~new_n34065_;
  assign new_n34067_ = ~new_n34063_ & new_n34066_;
  assign new_n34068_ = ~new_n33871_ & ~new_n34067_;
  assign new_n34069_ = \b[16]  & ~new_n33860_;
  assign new_n34070_ = ~new_n33858_ & new_n34069_;
  assign new_n34071_ = ~new_n33862_ & ~new_n34070_;
  assign new_n34072_ = ~new_n34068_ & new_n34071_;
  assign new_n34073_ = ~new_n33862_ & ~new_n34072_;
  assign new_n34074_ = \b[17]  & ~new_n33851_;
  assign new_n34075_ = ~new_n33849_ & new_n34074_;
  assign new_n34076_ = ~new_n33853_ & ~new_n34075_;
  assign new_n34077_ = ~new_n34073_ & new_n34076_;
  assign new_n34078_ = ~new_n33853_ & ~new_n34077_;
  assign new_n34079_ = \b[18]  & ~new_n33842_;
  assign new_n34080_ = ~new_n33840_ & new_n34079_;
  assign new_n34081_ = ~new_n33844_ & ~new_n34080_;
  assign new_n34082_ = ~new_n34078_ & new_n34081_;
  assign new_n34083_ = ~new_n33844_ & ~new_n34082_;
  assign new_n34084_ = \b[19]  & ~new_n33833_;
  assign new_n34085_ = ~new_n33831_ & new_n34084_;
  assign new_n34086_ = ~new_n33835_ & ~new_n34085_;
  assign new_n34087_ = ~new_n34083_ & new_n34086_;
  assign new_n34088_ = ~new_n33835_ & ~new_n34087_;
  assign new_n34089_ = \b[20]  & ~new_n33824_;
  assign new_n34090_ = ~new_n33822_ & new_n34089_;
  assign new_n34091_ = ~new_n33826_ & ~new_n34090_;
  assign new_n34092_ = ~new_n34088_ & new_n34091_;
  assign new_n34093_ = ~new_n33826_ & ~new_n34092_;
  assign new_n34094_ = \b[21]  & ~new_n33815_;
  assign new_n34095_ = ~new_n33813_ & new_n34094_;
  assign new_n34096_ = ~new_n33817_ & ~new_n34095_;
  assign new_n34097_ = ~new_n34093_ & new_n34096_;
  assign new_n34098_ = ~new_n33817_ & ~new_n34097_;
  assign new_n34099_ = \b[22]  & ~new_n33806_;
  assign new_n34100_ = ~new_n33804_ & new_n34099_;
  assign new_n34101_ = ~new_n33808_ & ~new_n34100_;
  assign new_n34102_ = ~new_n34098_ & new_n34101_;
  assign new_n34103_ = ~new_n33808_ & ~new_n34102_;
  assign new_n34104_ = \b[23]  & ~new_n33797_;
  assign new_n34105_ = ~new_n33795_ & new_n34104_;
  assign new_n34106_ = ~new_n33799_ & ~new_n34105_;
  assign new_n34107_ = ~new_n34103_ & new_n34106_;
  assign new_n34108_ = ~new_n33799_ & ~new_n34107_;
  assign new_n34109_ = \b[24]  & ~new_n33788_;
  assign new_n34110_ = ~new_n33786_ & new_n34109_;
  assign new_n34111_ = ~new_n33790_ & ~new_n34110_;
  assign new_n34112_ = ~new_n34108_ & new_n34111_;
  assign new_n34113_ = ~new_n33790_ & ~new_n34112_;
  assign new_n34114_ = \b[25]  & ~new_n33779_;
  assign new_n34115_ = ~new_n33777_ & new_n34114_;
  assign new_n34116_ = ~new_n33781_ & ~new_n34115_;
  assign new_n34117_ = ~new_n34113_ & new_n34116_;
  assign new_n34118_ = ~new_n33781_ & ~new_n34117_;
  assign new_n34119_ = \b[26]  & ~new_n33759_;
  assign new_n34120_ = ~new_n33757_ & new_n34119_;
  assign new_n34121_ = ~new_n33772_ & ~new_n34120_;
  assign new_n34122_ = ~new_n34118_ & new_n34121_;
  assign new_n34123_ = ~new_n33772_ & ~new_n34122_;
  assign new_n34124_ = \b[27]  & ~new_n33769_;
  assign new_n34125_ = ~new_n33767_ & new_n34124_;
  assign new_n34126_ = ~new_n33771_ & ~new_n34125_;
  assign new_n34127_ = ~new_n34123_ & new_n34126_;
  assign new_n34128_ = ~new_n33771_ & ~new_n34127_;
  assign new_n34129_ = new_n5926_ & ~new_n34128_;
  assign new_n34130_ = ~new_n33760_ & ~new_n34129_;
  assign new_n34131_ = ~new_n33781_ & new_n34121_;
  assign new_n34132_ = ~new_n34117_ & new_n34131_;
  assign new_n34133_ = ~new_n34118_ & ~new_n34121_;
  assign new_n34134_ = ~new_n34132_ & ~new_n34133_;
  assign new_n34135_ = new_n5926_ & ~new_n34134_;
  assign new_n34136_ = ~new_n34128_ & new_n34135_;
  assign new_n34137_ = ~new_n34130_ & ~new_n34136_;
  assign new_n34138_ = ~new_n33770_ & ~new_n34129_;
  assign new_n34139_ = ~new_n33772_ & new_n34126_;
  assign new_n34140_ = ~new_n34122_ & new_n34139_;
  assign new_n34141_ = ~new_n34123_ & ~new_n34126_;
  assign new_n34142_ = ~new_n34140_ & ~new_n34141_;
  assign new_n34143_ = new_n34129_ & ~new_n34142_;
  assign new_n34144_ = ~new_n34138_ & ~new_n34143_;
  assign new_n34145_ = ~\b[28]  & ~new_n34144_;
  assign new_n34146_ = ~\b[27]  & ~new_n34137_;
  assign new_n34147_ = ~new_n33780_ & ~new_n34129_;
  assign new_n34148_ = ~new_n33790_ & new_n34116_;
  assign new_n34149_ = ~new_n34112_ & new_n34148_;
  assign new_n34150_ = ~new_n34113_ & ~new_n34116_;
  assign new_n34151_ = ~new_n34149_ & ~new_n34150_;
  assign new_n34152_ = new_n5926_ & ~new_n34151_;
  assign new_n34153_ = ~new_n34128_ & new_n34152_;
  assign new_n34154_ = ~new_n34147_ & ~new_n34153_;
  assign new_n34155_ = ~\b[26]  & ~new_n34154_;
  assign new_n34156_ = ~new_n33789_ & ~new_n34129_;
  assign new_n34157_ = ~new_n33799_ & new_n34111_;
  assign new_n34158_ = ~new_n34107_ & new_n34157_;
  assign new_n34159_ = ~new_n34108_ & ~new_n34111_;
  assign new_n34160_ = ~new_n34158_ & ~new_n34159_;
  assign new_n34161_ = new_n5926_ & ~new_n34160_;
  assign new_n34162_ = ~new_n34128_ & new_n34161_;
  assign new_n34163_ = ~new_n34156_ & ~new_n34162_;
  assign new_n34164_ = ~\b[25]  & ~new_n34163_;
  assign new_n34165_ = ~new_n33798_ & ~new_n34129_;
  assign new_n34166_ = ~new_n33808_ & new_n34106_;
  assign new_n34167_ = ~new_n34102_ & new_n34166_;
  assign new_n34168_ = ~new_n34103_ & ~new_n34106_;
  assign new_n34169_ = ~new_n34167_ & ~new_n34168_;
  assign new_n34170_ = new_n5926_ & ~new_n34169_;
  assign new_n34171_ = ~new_n34128_ & new_n34170_;
  assign new_n34172_ = ~new_n34165_ & ~new_n34171_;
  assign new_n34173_ = ~\b[24]  & ~new_n34172_;
  assign new_n34174_ = ~new_n33807_ & ~new_n34129_;
  assign new_n34175_ = ~new_n33817_ & new_n34101_;
  assign new_n34176_ = ~new_n34097_ & new_n34175_;
  assign new_n34177_ = ~new_n34098_ & ~new_n34101_;
  assign new_n34178_ = ~new_n34176_ & ~new_n34177_;
  assign new_n34179_ = new_n5926_ & ~new_n34178_;
  assign new_n34180_ = ~new_n34128_ & new_n34179_;
  assign new_n34181_ = ~new_n34174_ & ~new_n34180_;
  assign new_n34182_ = ~\b[23]  & ~new_n34181_;
  assign new_n34183_ = ~new_n33816_ & ~new_n34129_;
  assign new_n34184_ = ~new_n33826_ & new_n34096_;
  assign new_n34185_ = ~new_n34092_ & new_n34184_;
  assign new_n34186_ = ~new_n34093_ & ~new_n34096_;
  assign new_n34187_ = ~new_n34185_ & ~new_n34186_;
  assign new_n34188_ = new_n5926_ & ~new_n34187_;
  assign new_n34189_ = ~new_n34128_ & new_n34188_;
  assign new_n34190_ = ~new_n34183_ & ~new_n34189_;
  assign new_n34191_ = ~\b[22]  & ~new_n34190_;
  assign new_n34192_ = ~new_n33825_ & ~new_n34129_;
  assign new_n34193_ = ~new_n33835_ & new_n34091_;
  assign new_n34194_ = ~new_n34087_ & new_n34193_;
  assign new_n34195_ = ~new_n34088_ & ~new_n34091_;
  assign new_n34196_ = ~new_n34194_ & ~new_n34195_;
  assign new_n34197_ = new_n5926_ & ~new_n34196_;
  assign new_n34198_ = ~new_n34128_ & new_n34197_;
  assign new_n34199_ = ~new_n34192_ & ~new_n34198_;
  assign new_n34200_ = ~\b[21]  & ~new_n34199_;
  assign new_n34201_ = ~new_n33834_ & ~new_n34129_;
  assign new_n34202_ = ~new_n33844_ & new_n34086_;
  assign new_n34203_ = ~new_n34082_ & new_n34202_;
  assign new_n34204_ = ~new_n34083_ & ~new_n34086_;
  assign new_n34205_ = ~new_n34203_ & ~new_n34204_;
  assign new_n34206_ = new_n5926_ & ~new_n34205_;
  assign new_n34207_ = ~new_n34128_ & new_n34206_;
  assign new_n34208_ = ~new_n34201_ & ~new_n34207_;
  assign new_n34209_ = ~\b[20]  & ~new_n34208_;
  assign new_n34210_ = ~new_n33843_ & ~new_n34129_;
  assign new_n34211_ = ~new_n33853_ & new_n34081_;
  assign new_n34212_ = ~new_n34077_ & new_n34211_;
  assign new_n34213_ = ~new_n34078_ & ~new_n34081_;
  assign new_n34214_ = ~new_n34212_ & ~new_n34213_;
  assign new_n34215_ = new_n5926_ & ~new_n34214_;
  assign new_n34216_ = ~new_n34128_ & new_n34215_;
  assign new_n34217_ = ~new_n34210_ & ~new_n34216_;
  assign new_n34218_ = ~\b[19]  & ~new_n34217_;
  assign new_n34219_ = ~new_n33852_ & ~new_n34129_;
  assign new_n34220_ = ~new_n33862_ & new_n34076_;
  assign new_n34221_ = ~new_n34072_ & new_n34220_;
  assign new_n34222_ = ~new_n34073_ & ~new_n34076_;
  assign new_n34223_ = ~new_n34221_ & ~new_n34222_;
  assign new_n34224_ = new_n5926_ & ~new_n34223_;
  assign new_n34225_ = ~new_n34128_ & new_n34224_;
  assign new_n34226_ = ~new_n34219_ & ~new_n34225_;
  assign new_n34227_ = ~\b[18]  & ~new_n34226_;
  assign new_n34228_ = ~new_n33861_ & ~new_n34129_;
  assign new_n34229_ = ~new_n33871_ & new_n34071_;
  assign new_n34230_ = ~new_n34067_ & new_n34229_;
  assign new_n34231_ = ~new_n34068_ & ~new_n34071_;
  assign new_n34232_ = ~new_n34230_ & ~new_n34231_;
  assign new_n34233_ = new_n5926_ & ~new_n34232_;
  assign new_n34234_ = ~new_n34128_ & new_n34233_;
  assign new_n34235_ = ~new_n34228_ & ~new_n34234_;
  assign new_n34236_ = ~\b[17]  & ~new_n34235_;
  assign new_n34237_ = ~new_n33870_ & ~new_n34129_;
  assign new_n34238_ = ~new_n33880_ & new_n34066_;
  assign new_n34239_ = ~new_n34062_ & new_n34238_;
  assign new_n34240_ = ~new_n34063_ & ~new_n34066_;
  assign new_n34241_ = ~new_n34239_ & ~new_n34240_;
  assign new_n34242_ = new_n5926_ & ~new_n34241_;
  assign new_n34243_ = ~new_n34128_ & new_n34242_;
  assign new_n34244_ = ~new_n34237_ & ~new_n34243_;
  assign new_n34245_ = ~\b[16]  & ~new_n34244_;
  assign new_n34246_ = ~new_n33879_ & ~new_n34129_;
  assign new_n34247_ = ~new_n33889_ & new_n34061_;
  assign new_n34248_ = ~new_n34057_ & new_n34247_;
  assign new_n34249_ = ~new_n34058_ & ~new_n34061_;
  assign new_n34250_ = ~new_n34248_ & ~new_n34249_;
  assign new_n34251_ = new_n5926_ & ~new_n34250_;
  assign new_n34252_ = ~new_n34128_ & new_n34251_;
  assign new_n34253_ = ~new_n34246_ & ~new_n34252_;
  assign new_n34254_ = ~\b[15]  & ~new_n34253_;
  assign new_n34255_ = ~new_n33888_ & ~new_n34129_;
  assign new_n34256_ = ~new_n33898_ & new_n34056_;
  assign new_n34257_ = ~new_n34052_ & new_n34256_;
  assign new_n34258_ = ~new_n34053_ & ~new_n34056_;
  assign new_n34259_ = ~new_n34257_ & ~new_n34258_;
  assign new_n34260_ = new_n5926_ & ~new_n34259_;
  assign new_n34261_ = ~new_n34128_ & new_n34260_;
  assign new_n34262_ = ~new_n34255_ & ~new_n34261_;
  assign new_n34263_ = ~\b[14]  & ~new_n34262_;
  assign new_n34264_ = ~new_n33897_ & ~new_n34129_;
  assign new_n34265_ = ~new_n33907_ & new_n34051_;
  assign new_n34266_ = ~new_n34047_ & new_n34265_;
  assign new_n34267_ = ~new_n34048_ & ~new_n34051_;
  assign new_n34268_ = ~new_n34266_ & ~new_n34267_;
  assign new_n34269_ = new_n5926_ & ~new_n34268_;
  assign new_n34270_ = ~new_n34128_ & new_n34269_;
  assign new_n34271_ = ~new_n34264_ & ~new_n34270_;
  assign new_n34272_ = ~\b[13]  & ~new_n34271_;
  assign new_n34273_ = ~new_n33906_ & ~new_n34129_;
  assign new_n34274_ = ~new_n33916_ & new_n34046_;
  assign new_n34275_ = ~new_n34042_ & new_n34274_;
  assign new_n34276_ = ~new_n34043_ & ~new_n34046_;
  assign new_n34277_ = ~new_n34275_ & ~new_n34276_;
  assign new_n34278_ = new_n5926_ & ~new_n34277_;
  assign new_n34279_ = ~new_n34128_ & new_n34278_;
  assign new_n34280_ = ~new_n34273_ & ~new_n34279_;
  assign new_n34281_ = ~\b[12]  & ~new_n34280_;
  assign new_n34282_ = ~new_n33915_ & ~new_n34129_;
  assign new_n34283_ = ~new_n33925_ & new_n34041_;
  assign new_n34284_ = ~new_n34037_ & new_n34283_;
  assign new_n34285_ = ~new_n34038_ & ~new_n34041_;
  assign new_n34286_ = ~new_n34284_ & ~new_n34285_;
  assign new_n34287_ = new_n5926_ & ~new_n34286_;
  assign new_n34288_ = ~new_n34128_ & new_n34287_;
  assign new_n34289_ = ~new_n34282_ & ~new_n34288_;
  assign new_n34290_ = ~\b[11]  & ~new_n34289_;
  assign new_n34291_ = ~new_n33924_ & ~new_n34129_;
  assign new_n34292_ = ~new_n33934_ & new_n34036_;
  assign new_n34293_ = ~new_n34032_ & new_n34292_;
  assign new_n34294_ = ~new_n34033_ & ~new_n34036_;
  assign new_n34295_ = ~new_n34293_ & ~new_n34294_;
  assign new_n34296_ = new_n5926_ & ~new_n34295_;
  assign new_n34297_ = ~new_n34128_ & new_n34296_;
  assign new_n34298_ = ~new_n34291_ & ~new_n34297_;
  assign new_n34299_ = ~\b[10]  & ~new_n34298_;
  assign new_n34300_ = ~new_n33933_ & ~new_n34129_;
  assign new_n34301_ = ~new_n33943_ & new_n34031_;
  assign new_n34302_ = ~new_n34027_ & new_n34301_;
  assign new_n34303_ = ~new_n34028_ & ~new_n34031_;
  assign new_n34304_ = ~new_n34302_ & ~new_n34303_;
  assign new_n34305_ = new_n5926_ & ~new_n34304_;
  assign new_n34306_ = ~new_n34128_ & new_n34305_;
  assign new_n34307_ = ~new_n34300_ & ~new_n34306_;
  assign new_n34308_ = ~\b[9]  & ~new_n34307_;
  assign new_n34309_ = ~new_n33942_ & ~new_n34129_;
  assign new_n34310_ = ~new_n33952_ & new_n34026_;
  assign new_n34311_ = ~new_n34022_ & new_n34310_;
  assign new_n34312_ = ~new_n34023_ & ~new_n34026_;
  assign new_n34313_ = ~new_n34311_ & ~new_n34312_;
  assign new_n34314_ = new_n5926_ & ~new_n34313_;
  assign new_n34315_ = ~new_n34128_ & new_n34314_;
  assign new_n34316_ = ~new_n34309_ & ~new_n34315_;
  assign new_n34317_ = ~\b[8]  & ~new_n34316_;
  assign new_n34318_ = ~new_n33951_ & ~new_n34129_;
  assign new_n34319_ = ~new_n33961_ & new_n34021_;
  assign new_n34320_ = ~new_n34017_ & new_n34319_;
  assign new_n34321_ = ~new_n34018_ & ~new_n34021_;
  assign new_n34322_ = ~new_n34320_ & ~new_n34321_;
  assign new_n34323_ = new_n5926_ & ~new_n34322_;
  assign new_n34324_ = ~new_n34128_ & new_n34323_;
  assign new_n34325_ = ~new_n34318_ & ~new_n34324_;
  assign new_n34326_ = ~\b[7]  & ~new_n34325_;
  assign new_n34327_ = ~new_n33960_ & ~new_n34129_;
  assign new_n34328_ = ~new_n33970_ & new_n34016_;
  assign new_n34329_ = ~new_n34012_ & new_n34328_;
  assign new_n34330_ = ~new_n34013_ & ~new_n34016_;
  assign new_n34331_ = ~new_n34329_ & ~new_n34330_;
  assign new_n34332_ = new_n5926_ & ~new_n34331_;
  assign new_n34333_ = ~new_n34128_ & new_n34332_;
  assign new_n34334_ = ~new_n34327_ & ~new_n34333_;
  assign new_n34335_ = ~\b[6]  & ~new_n34334_;
  assign new_n34336_ = ~new_n33969_ & ~new_n34129_;
  assign new_n34337_ = ~new_n33979_ & new_n34011_;
  assign new_n34338_ = ~new_n34007_ & new_n34337_;
  assign new_n34339_ = ~new_n34008_ & ~new_n34011_;
  assign new_n34340_ = ~new_n34338_ & ~new_n34339_;
  assign new_n34341_ = new_n5926_ & ~new_n34340_;
  assign new_n34342_ = ~new_n34128_ & new_n34341_;
  assign new_n34343_ = ~new_n34336_ & ~new_n34342_;
  assign new_n34344_ = ~\b[5]  & ~new_n34343_;
  assign new_n34345_ = ~new_n33978_ & ~new_n34129_;
  assign new_n34346_ = ~new_n33987_ & new_n34006_;
  assign new_n34347_ = ~new_n34002_ & new_n34346_;
  assign new_n34348_ = ~new_n34003_ & ~new_n34006_;
  assign new_n34349_ = ~new_n34347_ & ~new_n34348_;
  assign new_n34350_ = new_n5926_ & ~new_n34349_;
  assign new_n34351_ = ~new_n34128_ & new_n34350_;
  assign new_n34352_ = ~new_n34345_ & ~new_n34351_;
  assign new_n34353_ = ~\b[4]  & ~new_n34352_;
  assign new_n34354_ = ~new_n33986_ & ~new_n34129_;
  assign new_n34355_ = ~new_n33997_ & new_n34001_;
  assign new_n34356_ = ~new_n33996_ & new_n34355_;
  assign new_n34357_ = ~new_n33998_ & ~new_n34001_;
  assign new_n34358_ = ~new_n34356_ & ~new_n34357_;
  assign new_n34359_ = new_n5926_ & ~new_n34358_;
  assign new_n34360_ = ~new_n34128_ & new_n34359_;
  assign new_n34361_ = ~new_n34354_ & ~new_n34360_;
  assign new_n34362_ = ~\b[3]  & ~new_n34361_;
  assign new_n34363_ = ~new_n33991_ & ~new_n34129_;
  assign new_n34364_ = new_n5791_ & ~new_n33994_;
  assign new_n34365_ = ~new_n33992_ & new_n34364_;
  assign new_n34366_ = new_n5926_ & ~new_n34365_;
  assign new_n34367_ = ~new_n33996_ & new_n34366_;
  assign new_n34368_ = ~new_n34128_ & new_n34367_;
  assign new_n34369_ = ~new_n34363_ & ~new_n34368_;
  assign new_n34370_ = ~\b[2]  & ~new_n34369_;
  assign new_n34371_ = new_n6172_ & ~new_n34128_;
  assign new_n34372_ = \a[36]  & ~new_n34371_;
  assign new_n34373_ = new_n6177_ & ~new_n34128_;
  assign new_n34374_ = ~new_n34372_ & ~new_n34373_;
  assign new_n34375_ = \b[1]  & ~new_n34374_;
  assign new_n34376_ = ~\b[1]  & ~new_n34373_;
  assign new_n34377_ = ~new_n34372_ & new_n34376_;
  assign new_n34378_ = ~new_n34375_ & ~new_n34377_;
  assign new_n34379_ = ~new_n6184_ & ~new_n34378_;
  assign new_n34380_ = ~\b[1]  & ~new_n34374_;
  assign new_n34381_ = ~new_n34379_ & ~new_n34380_;
  assign new_n34382_ = \b[2]  & ~new_n34368_;
  assign new_n34383_ = ~new_n34363_ & new_n34382_;
  assign new_n34384_ = ~new_n34370_ & ~new_n34383_;
  assign new_n34385_ = ~new_n34381_ & new_n34384_;
  assign new_n34386_ = ~new_n34370_ & ~new_n34385_;
  assign new_n34387_ = \b[3]  & ~new_n34360_;
  assign new_n34388_ = ~new_n34354_ & new_n34387_;
  assign new_n34389_ = ~new_n34362_ & ~new_n34388_;
  assign new_n34390_ = ~new_n34386_ & new_n34389_;
  assign new_n34391_ = ~new_n34362_ & ~new_n34390_;
  assign new_n34392_ = \b[4]  & ~new_n34351_;
  assign new_n34393_ = ~new_n34345_ & new_n34392_;
  assign new_n34394_ = ~new_n34353_ & ~new_n34393_;
  assign new_n34395_ = ~new_n34391_ & new_n34394_;
  assign new_n34396_ = ~new_n34353_ & ~new_n34395_;
  assign new_n34397_ = \b[5]  & ~new_n34342_;
  assign new_n34398_ = ~new_n34336_ & new_n34397_;
  assign new_n34399_ = ~new_n34344_ & ~new_n34398_;
  assign new_n34400_ = ~new_n34396_ & new_n34399_;
  assign new_n34401_ = ~new_n34344_ & ~new_n34400_;
  assign new_n34402_ = \b[6]  & ~new_n34333_;
  assign new_n34403_ = ~new_n34327_ & new_n34402_;
  assign new_n34404_ = ~new_n34335_ & ~new_n34403_;
  assign new_n34405_ = ~new_n34401_ & new_n34404_;
  assign new_n34406_ = ~new_n34335_ & ~new_n34405_;
  assign new_n34407_ = \b[7]  & ~new_n34324_;
  assign new_n34408_ = ~new_n34318_ & new_n34407_;
  assign new_n34409_ = ~new_n34326_ & ~new_n34408_;
  assign new_n34410_ = ~new_n34406_ & new_n34409_;
  assign new_n34411_ = ~new_n34326_ & ~new_n34410_;
  assign new_n34412_ = \b[8]  & ~new_n34315_;
  assign new_n34413_ = ~new_n34309_ & new_n34412_;
  assign new_n34414_ = ~new_n34317_ & ~new_n34413_;
  assign new_n34415_ = ~new_n34411_ & new_n34414_;
  assign new_n34416_ = ~new_n34317_ & ~new_n34415_;
  assign new_n34417_ = \b[9]  & ~new_n34306_;
  assign new_n34418_ = ~new_n34300_ & new_n34417_;
  assign new_n34419_ = ~new_n34308_ & ~new_n34418_;
  assign new_n34420_ = ~new_n34416_ & new_n34419_;
  assign new_n34421_ = ~new_n34308_ & ~new_n34420_;
  assign new_n34422_ = \b[10]  & ~new_n34297_;
  assign new_n34423_ = ~new_n34291_ & new_n34422_;
  assign new_n34424_ = ~new_n34299_ & ~new_n34423_;
  assign new_n34425_ = ~new_n34421_ & new_n34424_;
  assign new_n34426_ = ~new_n34299_ & ~new_n34425_;
  assign new_n34427_ = \b[11]  & ~new_n34288_;
  assign new_n34428_ = ~new_n34282_ & new_n34427_;
  assign new_n34429_ = ~new_n34290_ & ~new_n34428_;
  assign new_n34430_ = ~new_n34426_ & new_n34429_;
  assign new_n34431_ = ~new_n34290_ & ~new_n34430_;
  assign new_n34432_ = \b[12]  & ~new_n34279_;
  assign new_n34433_ = ~new_n34273_ & new_n34432_;
  assign new_n34434_ = ~new_n34281_ & ~new_n34433_;
  assign new_n34435_ = ~new_n34431_ & new_n34434_;
  assign new_n34436_ = ~new_n34281_ & ~new_n34435_;
  assign new_n34437_ = \b[13]  & ~new_n34270_;
  assign new_n34438_ = ~new_n34264_ & new_n34437_;
  assign new_n34439_ = ~new_n34272_ & ~new_n34438_;
  assign new_n34440_ = ~new_n34436_ & new_n34439_;
  assign new_n34441_ = ~new_n34272_ & ~new_n34440_;
  assign new_n34442_ = \b[14]  & ~new_n34261_;
  assign new_n34443_ = ~new_n34255_ & new_n34442_;
  assign new_n34444_ = ~new_n34263_ & ~new_n34443_;
  assign new_n34445_ = ~new_n34441_ & new_n34444_;
  assign new_n34446_ = ~new_n34263_ & ~new_n34445_;
  assign new_n34447_ = \b[15]  & ~new_n34252_;
  assign new_n34448_ = ~new_n34246_ & new_n34447_;
  assign new_n34449_ = ~new_n34254_ & ~new_n34448_;
  assign new_n34450_ = ~new_n34446_ & new_n34449_;
  assign new_n34451_ = ~new_n34254_ & ~new_n34450_;
  assign new_n34452_ = \b[16]  & ~new_n34243_;
  assign new_n34453_ = ~new_n34237_ & new_n34452_;
  assign new_n34454_ = ~new_n34245_ & ~new_n34453_;
  assign new_n34455_ = ~new_n34451_ & new_n34454_;
  assign new_n34456_ = ~new_n34245_ & ~new_n34455_;
  assign new_n34457_ = \b[17]  & ~new_n34234_;
  assign new_n34458_ = ~new_n34228_ & new_n34457_;
  assign new_n34459_ = ~new_n34236_ & ~new_n34458_;
  assign new_n34460_ = ~new_n34456_ & new_n34459_;
  assign new_n34461_ = ~new_n34236_ & ~new_n34460_;
  assign new_n34462_ = \b[18]  & ~new_n34225_;
  assign new_n34463_ = ~new_n34219_ & new_n34462_;
  assign new_n34464_ = ~new_n34227_ & ~new_n34463_;
  assign new_n34465_ = ~new_n34461_ & new_n34464_;
  assign new_n34466_ = ~new_n34227_ & ~new_n34465_;
  assign new_n34467_ = \b[19]  & ~new_n34216_;
  assign new_n34468_ = ~new_n34210_ & new_n34467_;
  assign new_n34469_ = ~new_n34218_ & ~new_n34468_;
  assign new_n34470_ = ~new_n34466_ & new_n34469_;
  assign new_n34471_ = ~new_n34218_ & ~new_n34470_;
  assign new_n34472_ = \b[20]  & ~new_n34207_;
  assign new_n34473_ = ~new_n34201_ & new_n34472_;
  assign new_n34474_ = ~new_n34209_ & ~new_n34473_;
  assign new_n34475_ = ~new_n34471_ & new_n34474_;
  assign new_n34476_ = ~new_n34209_ & ~new_n34475_;
  assign new_n34477_ = \b[21]  & ~new_n34198_;
  assign new_n34478_ = ~new_n34192_ & new_n34477_;
  assign new_n34479_ = ~new_n34200_ & ~new_n34478_;
  assign new_n34480_ = ~new_n34476_ & new_n34479_;
  assign new_n34481_ = ~new_n34200_ & ~new_n34480_;
  assign new_n34482_ = \b[22]  & ~new_n34189_;
  assign new_n34483_ = ~new_n34183_ & new_n34482_;
  assign new_n34484_ = ~new_n34191_ & ~new_n34483_;
  assign new_n34485_ = ~new_n34481_ & new_n34484_;
  assign new_n34486_ = ~new_n34191_ & ~new_n34485_;
  assign new_n34487_ = \b[23]  & ~new_n34180_;
  assign new_n34488_ = ~new_n34174_ & new_n34487_;
  assign new_n34489_ = ~new_n34182_ & ~new_n34488_;
  assign new_n34490_ = ~new_n34486_ & new_n34489_;
  assign new_n34491_ = ~new_n34182_ & ~new_n34490_;
  assign new_n34492_ = \b[24]  & ~new_n34171_;
  assign new_n34493_ = ~new_n34165_ & new_n34492_;
  assign new_n34494_ = ~new_n34173_ & ~new_n34493_;
  assign new_n34495_ = ~new_n34491_ & new_n34494_;
  assign new_n34496_ = ~new_n34173_ & ~new_n34495_;
  assign new_n34497_ = \b[25]  & ~new_n34162_;
  assign new_n34498_ = ~new_n34156_ & new_n34497_;
  assign new_n34499_ = ~new_n34164_ & ~new_n34498_;
  assign new_n34500_ = ~new_n34496_ & new_n34499_;
  assign new_n34501_ = ~new_n34164_ & ~new_n34500_;
  assign new_n34502_ = \b[26]  & ~new_n34153_;
  assign new_n34503_ = ~new_n34147_ & new_n34502_;
  assign new_n34504_ = ~new_n34155_ & ~new_n34503_;
  assign new_n34505_ = ~new_n34501_ & new_n34504_;
  assign new_n34506_ = ~new_n34155_ & ~new_n34505_;
  assign new_n34507_ = \b[27]  & ~new_n34136_;
  assign new_n34508_ = ~new_n34130_ & new_n34507_;
  assign new_n34509_ = ~new_n34146_ & ~new_n34508_;
  assign new_n34510_ = ~new_n34506_ & new_n34509_;
  assign new_n34511_ = ~new_n34146_ & ~new_n34510_;
  assign new_n34512_ = \b[28]  & ~new_n34138_;
  assign new_n34513_ = ~new_n34143_ & new_n34512_;
  assign new_n34514_ = ~new_n34145_ & ~new_n34513_;
  assign new_n34515_ = ~new_n34511_ & new_n34514_;
  assign new_n34516_ = ~new_n34145_ & ~new_n34515_;
  assign new_n34517_ = new_n6324_ & ~new_n34516_;
  assign new_n34518_ = ~new_n34137_ & ~new_n34517_;
  assign new_n34519_ = ~new_n34155_ & new_n34509_;
  assign new_n34520_ = ~new_n34505_ & new_n34519_;
  assign new_n34521_ = ~new_n34506_ & ~new_n34509_;
  assign new_n34522_ = ~new_n34520_ & ~new_n34521_;
  assign new_n34523_ = new_n6324_ & ~new_n34522_;
  assign new_n34524_ = ~new_n34516_ & new_n34523_;
  assign new_n34525_ = ~new_n34518_ & ~new_n34524_;
  assign new_n34526_ = ~\b[28]  & ~new_n34525_;
  assign new_n34527_ = ~new_n34154_ & ~new_n34517_;
  assign new_n34528_ = ~new_n34164_ & new_n34504_;
  assign new_n34529_ = ~new_n34500_ & new_n34528_;
  assign new_n34530_ = ~new_n34501_ & ~new_n34504_;
  assign new_n34531_ = ~new_n34529_ & ~new_n34530_;
  assign new_n34532_ = new_n6324_ & ~new_n34531_;
  assign new_n34533_ = ~new_n34516_ & new_n34532_;
  assign new_n34534_ = ~new_n34527_ & ~new_n34533_;
  assign new_n34535_ = ~\b[27]  & ~new_n34534_;
  assign new_n34536_ = ~new_n34163_ & ~new_n34517_;
  assign new_n34537_ = ~new_n34173_ & new_n34499_;
  assign new_n34538_ = ~new_n34495_ & new_n34537_;
  assign new_n34539_ = ~new_n34496_ & ~new_n34499_;
  assign new_n34540_ = ~new_n34538_ & ~new_n34539_;
  assign new_n34541_ = new_n6324_ & ~new_n34540_;
  assign new_n34542_ = ~new_n34516_ & new_n34541_;
  assign new_n34543_ = ~new_n34536_ & ~new_n34542_;
  assign new_n34544_ = ~\b[26]  & ~new_n34543_;
  assign new_n34545_ = ~new_n34172_ & ~new_n34517_;
  assign new_n34546_ = ~new_n34182_ & new_n34494_;
  assign new_n34547_ = ~new_n34490_ & new_n34546_;
  assign new_n34548_ = ~new_n34491_ & ~new_n34494_;
  assign new_n34549_ = ~new_n34547_ & ~new_n34548_;
  assign new_n34550_ = new_n6324_ & ~new_n34549_;
  assign new_n34551_ = ~new_n34516_ & new_n34550_;
  assign new_n34552_ = ~new_n34545_ & ~new_n34551_;
  assign new_n34553_ = ~\b[25]  & ~new_n34552_;
  assign new_n34554_ = ~new_n34181_ & ~new_n34517_;
  assign new_n34555_ = ~new_n34191_ & new_n34489_;
  assign new_n34556_ = ~new_n34485_ & new_n34555_;
  assign new_n34557_ = ~new_n34486_ & ~new_n34489_;
  assign new_n34558_ = ~new_n34556_ & ~new_n34557_;
  assign new_n34559_ = new_n6324_ & ~new_n34558_;
  assign new_n34560_ = ~new_n34516_ & new_n34559_;
  assign new_n34561_ = ~new_n34554_ & ~new_n34560_;
  assign new_n34562_ = ~\b[24]  & ~new_n34561_;
  assign new_n34563_ = ~new_n34190_ & ~new_n34517_;
  assign new_n34564_ = ~new_n34200_ & new_n34484_;
  assign new_n34565_ = ~new_n34480_ & new_n34564_;
  assign new_n34566_ = ~new_n34481_ & ~new_n34484_;
  assign new_n34567_ = ~new_n34565_ & ~new_n34566_;
  assign new_n34568_ = new_n6324_ & ~new_n34567_;
  assign new_n34569_ = ~new_n34516_ & new_n34568_;
  assign new_n34570_ = ~new_n34563_ & ~new_n34569_;
  assign new_n34571_ = ~\b[23]  & ~new_n34570_;
  assign new_n34572_ = ~new_n34199_ & ~new_n34517_;
  assign new_n34573_ = ~new_n34209_ & new_n34479_;
  assign new_n34574_ = ~new_n34475_ & new_n34573_;
  assign new_n34575_ = ~new_n34476_ & ~new_n34479_;
  assign new_n34576_ = ~new_n34574_ & ~new_n34575_;
  assign new_n34577_ = new_n6324_ & ~new_n34576_;
  assign new_n34578_ = ~new_n34516_ & new_n34577_;
  assign new_n34579_ = ~new_n34572_ & ~new_n34578_;
  assign new_n34580_ = ~\b[22]  & ~new_n34579_;
  assign new_n34581_ = ~new_n34208_ & ~new_n34517_;
  assign new_n34582_ = ~new_n34218_ & new_n34474_;
  assign new_n34583_ = ~new_n34470_ & new_n34582_;
  assign new_n34584_ = ~new_n34471_ & ~new_n34474_;
  assign new_n34585_ = ~new_n34583_ & ~new_n34584_;
  assign new_n34586_ = new_n6324_ & ~new_n34585_;
  assign new_n34587_ = ~new_n34516_ & new_n34586_;
  assign new_n34588_ = ~new_n34581_ & ~new_n34587_;
  assign new_n34589_ = ~\b[21]  & ~new_n34588_;
  assign new_n34590_ = ~new_n34217_ & ~new_n34517_;
  assign new_n34591_ = ~new_n34227_ & new_n34469_;
  assign new_n34592_ = ~new_n34465_ & new_n34591_;
  assign new_n34593_ = ~new_n34466_ & ~new_n34469_;
  assign new_n34594_ = ~new_n34592_ & ~new_n34593_;
  assign new_n34595_ = new_n6324_ & ~new_n34594_;
  assign new_n34596_ = ~new_n34516_ & new_n34595_;
  assign new_n34597_ = ~new_n34590_ & ~new_n34596_;
  assign new_n34598_ = ~\b[20]  & ~new_n34597_;
  assign new_n34599_ = ~new_n34226_ & ~new_n34517_;
  assign new_n34600_ = ~new_n34236_ & new_n34464_;
  assign new_n34601_ = ~new_n34460_ & new_n34600_;
  assign new_n34602_ = ~new_n34461_ & ~new_n34464_;
  assign new_n34603_ = ~new_n34601_ & ~new_n34602_;
  assign new_n34604_ = new_n6324_ & ~new_n34603_;
  assign new_n34605_ = ~new_n34516_ & new_n34604_;
  assign new_n34606_ = ~new_n34599_ & ~new_n34605_;
  assign new_n34607_ = ~\b[19]  & ~new_n34606_;
  assign new_n34608_ = ~new_n34235_ & ~new_n34517_;
  assign new_n34609_ = ~new_n34245_ & new_n34459_;
  assign new_n34610_ = ~new_n34455_ & new_n34609_;
  assign new_n34611_ = ~new_n34456_ & ~new_n34459_;
  assign new_n34612_ = ~new_n34610_ & ~new_n34611_;
  assign new_n34613_ = new_n6324_ & ~new_n34612_;
  assign new_n34614_ = ~new_n34516_ & new_n34613_;
  assign new_n34615_ = ~new_n34608_ & ~new_n34614_;
  assign new_n34616_ = ~\b[18]  & ~new_n34615_;
  assign new_n34617_ = ~new_n34244_ & ~new_n34517_;
  assign new_n34618_ = ~new_n34254_ & new_n34454_;
  assign new_n34619_ = ~new_n34450_ & new_n34618_;
  assign new_n34620_ = ~new_n34451_ & ~new_n34454_;
  assign new_n34621_ = ~new_n34619_ & ~new_n34620_;
  assign new_n34622_ = new_n6324_ & ~new_n34621_;
  assign new_n34623_ = ~new_n34516_ & new_n34622_;
  assign new_n34624_ = ~new_n34617_ & ~new_n34623_;
  assign new_n34625_ = ~\b[17]  & ~new_n34624_;
  assign new_n34626_ = ~new_n34253_ & ~new_n34517_;
  assign new_n34627_ = ~new_n34263_ & new_n34449_;
  assign new_n34628_ = ~new_n34445_ & new_n34627_;
  assign new_n34629_ = ~new_n34446_ & ~new_n34449_;
  assign new_n34630_ = ~new_n34628_ & ~new_n34629_;
  assign new_n34631_ = new_n6324_ & ~new_n34630_;
  assign new_n34632_ = ~new_n34516_ & new_n34631_;
  assign new_n34633_ = ~new_n34626_ & ~new_n34632_;
  assign new_n34634_ = ~\b[16]  & ~new_n34633_;
  assign new_n34635_ = ~new_n34262_ & ~new_n34517_;
  assign new_n34636_ = ~new_n34272_ & new_n34444_;
  assign new_n34637_ = ~new_n34440_ & new_n34636_;
  assign new_n34638_ = ~new_n34441_ & ~new_n34444_;
  assign new_n34639_ = ~new_n34637_ & ~new_n34638_;
  assign new_n34640_ = new_n6324_ & ~new_n34639_;
  assign new_n34641_ = ~new_n34516_ & new_n34640_;
  assign new_n34642_ = ~new_n34635_ & ~new_n34641_;
  assign new_n34643_ = ~\b[15]  & ~new_n34642_;
  assign new_n34644_ = ~new_n34271_ & ~new_n34517_;
  assign new_n34645_ = ~new_n34281_ & new_n34439_;
  assign new_n34646_ = ~new_n34435_ & new_n34645_;
  assign new_n34647_ = ~new_n34436_ & ~new_n34439_;
  assign new_n34648_ = ~new_n34646_ & ~new_n34647_;
  assign new_n34649_ = new_n6324_ & ~new_n34648_;
  assign new_n34650_ = ~new_n34516_ & new_n34649_;
  assign new_n34651_ = ~new_n34644_ & ~new_n34650_;
  assign new_n34652_ = ~\b[14]  & ~new_n34651_;
  assign new_n34653_ = ~new_n34280_ & ~new_n34517_;
  assign new_n34654_ = ~new_n34290_ & new_n34434_;
  assign new_n34655_ = ~new_n34430_ & new_n34654_;
  assign new_n34656_ = ~new_n34431_ & ~new_n34434_;
  assign new_n34657_ = ~new_n34655_ & ~new_n34656_;
  assign new_n34658_ = new_n6324_ & ~new_n34657_;
  assign new_n34659_ = ~new_n34516_ & new_n34658_;
  assign new_n34660_ = ~new_n34653_ & ~new_n34659_;
  assign new_n34661_ = ~\b[13]  & ~new_n34660_;
  assign new_n34662_ = ~new_n34289_ & ~new_n34517_;
  assign new_n34663_ = ~new_n34299_ & new_n34429_;
  assign new_n34664_ = ~new_n34425_ & new_n34663_;
  assign new_n34665_ = ~new_n34426_ & ~new_n34429_;
  assign new_n34666_ = ~new_n34664_ & ~new_n34665_;
  assign new_n34667_ = new_n6324_ & ~new_n34666_;
  assign new_n34668_ = ~new_n34516_ & new_n34667_;
  assign new_n34669_ = ~new_n34662_ & ~new_n34668_;
  assign new_n34670_ = ~\b[12]  & ~new_n34669_;
  assign new_n34671_ = ~new_n34298_ & ~new_n34517_;
  assign new_n34672_ = ~new_n34308_ & new_n34424_;
  assign new_n34673_ = ~new_n34420_ & new_n34672_;
  assign new_n34674_ = ~new_n34421_ & ~new_n34424_;
  assign new_n34675_ = ~new_n34673_ & ~new_n34674_;
  assign new_n34676_ = new_n6324_ & ~new_n34675_;
  assign new_n34677_ = ~new_n34516_ & new_n34676_;
  assign new_n34678_ = ~new_n34671_ & ~new_n34677_;
  assign new_n34679_ = ~\b[11]  & ~new_n34678_;
  assign new_n34680_ = ~new_n34307_ & ~new_n34517_;
  assign new_n34681_ = ~new_n34317_ & new_n34419_;
  assign new_n34682_ = ~new_n34415_ & new_n34681_;
  assign new_n34683_ = ~new_n34416_ & ~new_n34419_;
  assign new_n34684_ = ~new_n34682_ & ~new_n34683_;
  assign new_n34685_ = new_n6324_ & ~new_n34684_;
  assign new_n34686_ = ~new_n34516_ & new_n34685_;
  assign new_n34687_ = ~new_n34680_ & ~new_n34686_;
  assign new_n34688_ = ~\b[10]  & ~new_n34687_;
  assign new_n34689_ = ~new_n34316_ & ~new_n34517_;
  assign new_n34690_ = ~new_n34326_ & new_n34414_;
  assign new_n34691_ = ~new_n34410_ & new_n34690_;
  assign new_n34692_ = ~new_n34411_ & ~new_n34414_;
  assign new_n34693_ = ~new_n34691_ & ~new_n34692_;
  assign new_n34694_ = new_n6324_ & ~new_n34693_;
  assign new_n34695_ = ~new_n34516_ & new_n34694_;
  assign new_n34696_ = ~new_n34689_ & ~new_n34695_;
  assign new_n34697_ = ~\b[9]  & ~new_n34696_;
  assign new_n34698_ = ~new_n34325_ & ~new_n34517_;
  assign new_n34699_ = ~new_n34335_ & new_n34409_;
  assign new_n34700_ = ~new_n34405_ & new_n34699_;
  assign new_n34701_ = ~new_n34406_ & ~new_n34409_;
  assign new_n34702_ = ~new_n34700_ & ~new_n34701_;
  assign new_n34703_ = new_n6324_ & ~new_n34702_;
  assign new_n34704_ = ~new_n34516_ & new_n34703_;
  assign new_n34705_ = ~new_n34698_ & ~new_n34704_;
  assign new_n34706_ = ~\b[8]  & ~new_n34705_;
  assign new_n34707_ = ~new_n34334_ & ~new_n34517_;
  assign new_n34708_ = ~new_n34344_ & new_n34404_;
  assign new_n34709_ = ~new_n34400_ & new_n34708_;
  assign new_n34710_ = ~new_n34401_ & ~new_n34404_;
  assign new_n34711_ = ~new_n34709_ & ~new_n34710_;
  assign new_n34712_ = new_n6324_ & ~new_n34711_;
  assign new_n34713_ = ~new_n34516_ & new_n34712_;
  assign new_n34714_ = ~new_n34707_ & ~new_n34713_;
  assign new_n34715_ = ~\b[7]  & ~new_n34714_;
  assign new_n34716_ = ~new_n34343_ & ~new_n34517_;
  assign new_n34717_ = ~new_n34353_ & new_n34399_;
  assign new_n34718_ = ~new_n34395_ & new_n34717_;
  assign new_n34719_ = ~new_n34396_ & ~new_n34399_;
  assign new_n34720_ = ~new_n34718_ & ~new_n34719_;
  assign new_n34721_ = new_n6324_ & ~new_n34720_;
  assign new_n34722_ = ~new_n34516_ & new_n34721_;
  assign new_n34723_ = ~new_n34716_ & ~new_n34722_;
  assign new_n34724_ = ~\b[6]  & ~new_n34723_;
  assign new_n34725_ = ~new_n34352_ & ~new_n34517_;
  assign new_n34726_ = ~new_n34362_ & new_n34394_;
  assign new_n34727_ = ~new_n34390_ & new_n34726_;
  assign new_n34728_ = ~new_n34391_ & ~new_n34394_;
  assign new_n34729_ = ~new_n34727_ & ~new_n34728_;
  assign new_n34730_ = new_n6324_ & ~new_n34729_;
  assign new_n34731_ = ~new_n34516_ & new_n34730_;
  assign new_n34732_ = ~new_n34725_ & ~new_n34731_;
  assign new_n34733_ = ~\b[5]  & ~new_n34732_;
  assign new_n34734_ = ~new_n34361_ & ~new_n34517_;
  assign new_n34735_ = ~new_n34370_ & new_n34389_;
  assign new_n34736_ = ~new_n34385_ & new_n34735_;
  assign new_n34737_ = ~new_n34386_ & ~new_n34389_;
  assign new_n34738_ = ~new_n34736_ & ~new_n34737_;
  assign new_n34739_ = new_n6324_ & ~new_n34738_;
  assign new_n34740_ = ~new_n34516_ & new_n34739_;
  assign new_n34741_ = ~new_n34734_ & ~new_n34740_;
  assign new_n34742_ = ~\b[4]  & ~new_n34741_;
  assign new_n34743_ = ~new_n34369_ & ~new_n34517_;
  assign new_n34744_ = ~new_n34380_ & new_n34384_;
  assign new_n34745_ = ~new_n34379_ & new_n34744_;
  assign new_n34746_ = ~new_n34381_ & ~new_n34384_;
  assign new_n34747_ = ~new_n34745_ & ~new_n34746_;
  assign new_n34748_ = new_n6324_ & ~new_n34747_;
  assign new_n34749_ = ~new_n34516_ & new_n34748_;
  assign new_n34750_ = ~new_n34743_ & ~new_n34749_;
  assign new_n34751_ = ~\b[3]  & ~new_n34750_;
  assign new_n34752_ = ~new_n34374_ & ~new_n34517_;
  assign new_n34753_ = new_n6184_ & ~new_n34377_;
  assign new_n34754_ = ~new_n34375_ & new_n34753_;
  assign new_n34755_ = new_n6324_ & ~new_n34754_;
  assign new_n34756_ = ~new_n34379_ & new_n34755_;
  assign new_n34757_ = ~new_n34516_ & new_n34756_;
  assign new_n34758_ = ~new_n34752_ & ~new_n34757_;
  assign new_n34759_ = ~\b[2]  & ~new_n34758_;
  assign new_n34760_ = new_n6572_ & ~new_n34516_;
  assign new_n34761_ = \a[35]  & ~new_n34760_;
  assign new_n34762_ = new_n6577_ & ~new_n34516_;
  assign new_n34763_ = ~new_n34761_ & ~new_n34762_;
  assign new_n34764_ = \b[1]  & ~new_n34763_;
  assign new_n34765_ = ~\b[1]  & ~new_n34762_;
  assign new_n34766_ = ~new_n34761_ & new_n34765_;
  assign new_n34767_ = ~new_n34764_ & ~new_n34766_;
  assign new_n34768_ = ~new_n6584_ & ~new_n34767_;
  assign new_n34769_ = ~\b[1]  & ~new_n34763_;
  assign new_n34770_ = ~new_n34768_ & ~new_n34769_;
  assign new_n34771_ = \b[2]  & ~new_n34757_;
  assign new_n34772_ = ~new_n34752_ & new_n34771_;
  assign new_n34773_ = ~new_n34759_ & ~new_n34772_;
  assign new_n34774_ = ~new_n34770_ & new_n34773_;
  assign new_n34775_ = ~new_n34759_ & ~new_n34774_;
  assign new_n34776_ = \b[3]  & ~new_n34749_;
  assign new_n34777_ = ~new_n34743_ & new_n34776_;
  assign new_n34778_ = ~new_n34751_ & ~new_n34777_;
  assign new_n34779_ = ~new_n34775_ & new_n34778_;
  assign new_n34780_ = ~new_n34751_ & ~new_n34779_;
  assign new_n34781_ = \b[4]  & ~new_n34740_;
  assign new_n34782_ = ~new_n34734_ & new_n34781_;
  assign new_n34783_ = ~new_n34742_ & ~new_n34782_;
  assign new_n34784_ = ~new_n34780_ & new_n34783_;
  assign new_n34785_ = ~new_n34742_ & ~new_n34784_;
  assign new_n34786_ = \b[5]  & ~new_n34731_;
  assign new_n34787_ = ~new_n34725_ & new_n34786_;
  assign new_n34788_ = ~new_n34733_ & ~new_n34787_;
  assign new_n34789_ = ~new_n34785_ & new_n34788_;
  assign new_n34790_ = ~new_n34733_ & ~new_n34789_;
  assign new_n34791_ = \b[6]  & ~new_n34722_;
  assign new_n34792_ = ~new_n34716_ & new_n34791_;
  assign new_n34793_ = ~new_n34724_ & ~new_n34792_;
  assign new_n34794_ = ~new_n34790_ & new_n34793_;
  assign new_n34795_ = ~new_n34724_ & ~new_n34794_;
  assign new_n34796_ = \b[7]  & ~new_n34713_;
  assign new_n34797_ = ~new_n34707_ & new_n34796_;
  assign new_n34798_ = ~new_n34715_ & ~new_n34797_;
  assign new_n34799_ = ~new_n34795_ & new_n34798_;
  assign new_n34800_ = ~new_n34715_ & ~new_n34799_;
  assign new_n34801_ = \b[8]  & ~new_n34704_;
  assign new_n34802_ = ~new_n34698_ & new_n34801_;
  assign new_n34803_ = ~new_n34706_ & ~new_n34802_;
  assign new_n34804_ = ~new_n34800_ & new_n34803_;
  assign new_n34805_ = ~new_n34706_ & ~new_n34804_;
  assign new_n34806_ = \b[9]  & ~new_n34695_;
  assign new_n34807_ = ~new_n34689_ & new_n34806_;
  assign new_n34808_ = ~new_n34697_ & ~new_n34807_;
  assign new_n34809_ = ~new_n34805_ & new_n34808_;
  assign new_n34810_ = ~new_n34697_ & ~new_n34809_;
  assign new_n34811_ = \b[10]  & ~new_n34686_;
  assign new_n34812_ = ~new_n34680_ & new_n34811_;
  assign new_n34813_ = ~new_n34688_ & ~new_n34812_;
  assign new_n34814_ = ~new_n34810_ & new_n34813_;
  assign new_n34815_ = ~new_n34688_ & ~new_n34814_;
  assign new_n34816_ = \b[11]  & ~new_n34677_;
  assign new_n34817_ = ~new_n34671_ & new_n34816_;
  assign new_n34818_ = ~new_n34679_ & ~new_n34817_;
  assign new_n34819_ = ~new_n34815_ & new_n34818_;
  assign new_n34820_ = ~new_n34679_ & ~new_n34819_;
  assign new_n34821_ = \b[12]  & ~new_n34668_;
  assign new_n34822_ = ~new_n34662_ & new_n34821_;
  assign new_n34823_ = ~new_n34670_ & ~new_n34822_;
  assign new_n34824_ = ~new_n34820_ & new_n34823_;
  assign new_n34825_ = ~new_n34670_ & ~new_n34824_;
  assign new_n34826_ = \b[13]  & ~new_n34659_;
  assign new_n34827_ = ~new_n34653_ & new_n34826_;
  assign new_n34828_ = ~new_n34661_ & ~new_n34827_;
  assign new_n34829_ = ~new_n34825_ & new_n34828_;
  assign new_n34830_ = ~new_n34661_ & ~new_n34829_;
  assign new_n34831_ = \b[14]  & ~new_n34650_;
  assign new_n34832_ = ~new_n34644_ & new_n34831_;
  assign new_n34833_ = ~new_n34652_ & ~new_n34832_;
  assign new_n34834_ = ~new_n34830_ & new_n34833_;
  assign new_n34835_ = ~new_n34652_ & ~new_n34834_;
  assign new_n34836_ = \b[15]  & ~new_n34641_;
  assign new_n34837_ = ~new_n34635_ & new_n34836_;
  assign new_n34838_ = ~new_n34643_ & ~new_n34837_;
  assign new_n34839_ = ~new_n34835_ & new_n34838_;
  assign new_n34840_ = ~new_n34643_ & ~new_n34839_;
  assign new_n34841_ = \b[16]  & ~new_n34632_;
  assign new_n34842_ = ~new_n34626_ & new_n34841_;
  assign new_n34843_ = ~new_n34634_ & ~new_n34842_;
  assign new_n34844_ = ~new_n34840_ & new_n34843_;
  assign new_n34845_ = ~new_n34634_ & ~new_n34844_;
  assign new_n34846_ = \b[17]  & ~new_n34623_;
  assign new_n34847_ = ~new_n34617_ & new_n34846_;
  assign new_n34848_ = ~new_n34625_ & ~new_n34847_;
  assign new_n34849_ = ~new_n34845_ & new_n34848_;
  assign new_n34850_ = ~new_n34625_ & ~new_n34849_;
  assign new_n34851_ = \b[18]  & ~new_n34614_;
  assign new_n34852_ = ~new_n34608_ & new_n34851_;
  assign new_n34853_ = ~new_n34616_ & ~new_n34852_;
  assign new_n34854_ = ~new_n34850_ & new_n34853_;
  assign new_n34855_ = ~new_n34616_ & ~new_n34854_;
  assign new_n34856_ = \b[19]  & ~new_n34605_;
  assign new_n34857_ = ~new_n34599_ & new_n34856_;
  assign new_n34858_ = ~new_n34607_ & ~new_n34857_;
  assign new_n34859_ = ~new_n34855_ & new_n34858_;
  assign new_n34860_ = ~new_n34607_ & ~new_n34859_;
  assign new_n34861_ = \b[20]  & ~new_n34596_;
  assign new_n34862_ = ~new_n34590_ & new_n34861_;
  assign new_n34863_ = ~new_n34598_ & ~new_n34862_;
  assign new_n34864_ = ~new_n34860_ & new_n34863_;
  assign new_n34865_ = ~new_n34598_ & ~new_n34864_;
  assign new_n34866_ = \b[21]  & ~new_n34587_;
  assign new_n34867_ = ~new_n34581_ & new_n34866_;
  assign new_n34868_ = ~new_n34589_ & ~new_n34867_;
  assign new_n34869_ = ~new_n34865_ & new_n34868_;
  assign new_n34870_ = ~new_n34589_ & ~new_n34869_;
  assign new_n34871_ = \b[22]  & ~new_n34578_;
  assign new_n34872_ = ~new_n34572_ & new_n34871_;
  assign new_n34873_ = ~new_n34580_ & ~new_n34872_;
  assign new_n34874_ = ~new_n34870_ & new_n34873_;
  assign new_n34875_ = ~new_n34580_ & ~new_n34874_;
  assign new_n34876_ = \b[23]  & ~new_n34569_;
  assign new_n34877_ = ~new_n34563_ & new_n34876_;
  assign new_n34878_ = ~new_n34571_ & ~new_n34877_;
  assign new_n34879_ = ~new_n34875_ & new_n34878_;
  assign new_n34880_ = ~new_n34571_ & ~new_n34879_;
  assign new_n34881_ = \b[24]  & ~new_n34560_;
  assign new_n34882_ = ~new_n34554_ & new_n34881_;
  assign new_n34883_ = ~new_n34562_ & ~new_n34882_;
  assign new_n34884_ = ~new_n34880_ & new_n34883_;
  assign new_n34885_ = ~new_n34562_ & ~new_n34884_;
  assign new_n34886_ = \b[25]  & ~new_n34551_;
  assign new_n34887_ = ~new_n34545_ & new_n34886_;
  assign new_n34888_ = ~new_n34553_ & ~new_n34887_;
  assign new_n34889_ = ~new_n34885_ & new_n34888_;
  assign new_n34890_ = ~new_n34553_ & ~new_n34889_;
  assign new_n34891_ = \b[26]  & ~new_n34542_;
  assign new_n34892_ = ~new_n34536_ & new_n34891_;
  assign new_n34893_ = ~new_n34544_ & ~new_n34892_;
  assign new_n34894_ = ~new_n34890_ & new_n34893_;
  assign new_n34895_ = ~new_n34544_ & ~new_n34894_;
  assign new_n34896_ = \b[27]  & ~new_n34533_;
  assign new_n34897_ = ~new_n34527_ & new_n34896_;
  assign new_n34898_ = ~new_n34535_ & ~new_n34897_;
  assign new_n34899_ = ~new_n34895_ & new_n34898_;
  assign new_n34900_ = ~new_n34535_ & ~new_n34899_;
  assign new_n34901_ = \b[28]  & ~new_n34524_;
  assign new_n34902_ = ~new_n34518_ & new_n34901_;
  assign new_n34903_ = ~new_n34526_ & ~new_n34902_;
  assign new_n34904_ = ~new_n34900_ & new_n34903_;
  assign new_n34905_ = ~new_n34526_ & ~new_n34904_;
  assign new_n34906_ = ~new_n34144_ & ~new_n34517_;
  assign new_n34907_ = ~new_n34146_ & new_n34514_;
  assign new_n34908_ = ~new_n34510_ & new_n34907_;
  assign new_n34909_ = ~new_n34511_ & ~new_n34514_;
  assign new_n34910_ = ~new_n34908_ & ~new_n34909_;
  assign new_n34911_ = new_n34517_ & ~new_n34910_;
  assign new_n34912_ = ~new_n34906_ & ~new_n34911_;
  assign new_n34913_ = ~\b[29]  & ~new_n34912_;
  assign new_n34914_ = \b[29]  & ~new_n34906_;
  assign new_n34915_ = ~new_n34911_ & new_n34914_;
  assign new_n34916_ = new_n6735_ & ~new_n34915_;
  assign new_n34917_ = ~new_n34913_ & new_n34916_;
  assign new_n34918_ = ~new_n34905_ & new_n34917_;
  assign new_n34919_ = new_n6324_ & ~new_n34912_;
  assign new_n34920_ = ~new_n34918_ & ~new_n34919_;
  assign new_n34921_ = ~new_n34535_ & new_n34903_;
  assign new_n34922_ = ~new_n34899_ & new_n34921_;
  assign new_n34923_ = ~new_n34900_ & ~new_n34903_;
  assign new_n34924_ = ~new_n34922_ & ~new_n34923_;
  assign new_n34925_ = ~new_n34920_ & ~new_n34924_;
  assign new_n34926_ = ~new_n34525_ & ~new_n34919_;
  assign new_n34927_ = ~new_n34918_ & new_n34926_;
  assign new_n34928_ = ~new_n34925_ & ~new_n34927_;
  assign new_n34929_ = ~new_n34526_ & ~new_n34915_;
  assign new_n34930_ = ~new_n34913_ & new_n34929_;
  assign new_n34931_ = ~new_n34904_ & new_n34930_;
  assign new_n34932_ = ~new_n34913_ & ~new_n34915_;
  assign new_n34933_ = ~new_n34905_ & ~new_n34932_;
  assign new_n34934_ = ~new_n34931_ & ~new_n34933_;
  assign new_n34935_ = ~new_n34920_ & ~new_n34934_;
  assign new_n34936_ = ~new_n34912_ & ~new_n34919_;
  assign new_n34937_ = ~new_n34918_ & new_n34936_;
  assign new_n34938_ = ~new_n34935_ & ~new_n34937_;
  assign new_n34939_ = ~\b[30]  & ~new_n34938_;
  assign new_n34940_ = ~\b[29]  & ~new_n34928_;
  assign new_n34941_ = ~new_n34544_ & new_n34898_;
  assign new_n34942_ = ~new_n34894_ & new_n34941_;
  assign new_n34943_ = ~new_n34895_ & ~new_n34898_;
  assign new_n34944_ = ~new_n34942_ & ~new_n34943_;
  assign new_n34945_ = ~new_n34920_ & ~new_n34944_;
  assign new_n34946_ = ~new_n34534_ & ~new_n34919_;
  assign new_n34947_ = ~new_n34918_ & new_n34946_;
  assign new_n34948_ = ~new_n34945_ & ~new_n34947_;
  assign new_n34949_ = ~\b[28]  & ~new_n34948_;
  assign new_n34950_ = ~new_n34553_ & new_n34893_;
  assign new_n34951_ = ~new_n34889_ & new_n34950_;
  assign new_n34952_ = ~new_n34890_ & ~new_n34893_;
  assign new_n34953_ = ~new_n34951_ & ~new_n34952_;
  assign new_n34954_ = ~new_n34920_ & ~new_n34953_;
  assign new_n34955_ = ~new_n34543_ & ~new_n34919_;
  assign new_n34956_ = ~new_n34918_ & new_n34955_;
  assign new_n34957_ = ~new_n34954_ & ~new_n34956_;
  assign new_n34958_ = ~\b[27]  & ~new_n34957_;
  assign new_n34959_ = ~new_n34562_ & new_n34888_;
  assign new_n34960_ = ~new_n34884_ & new_n34959_;
  assign new_n34961_ = ~new_n34885_ & ~new_n34888_;
  assign new_n34962_ = ~new_n34960_ & ~new_n34961_;
  assign new_n34963_ = ~new_n34920_ & ~new_n34962_;
  assign new_n34964_ = ~new_n34552_ & ~new_n34919_;
  assign new_n34965_ = ~new_n34918_ & new_n34964_;
  assign new_n34966_ = ~new_n34963_ & ~new_n34965_;
  assign new_n34967_ = ~\b[26]  & ~new_n34966_;
  assign new_n34968_ = ~new_n34571_ & new_n34883_;
  assign new_n34969_ = ~new_n34879_ & new_n34968_;
  assign new_n34970_ = ~new_n34880_ & ~new_n34883_;
  assign new_n34971_ = ~new_n34969_ & ~new_n34970_;
  assign new_n34972_ = ~new_n34920_ & ~new_n34971_;
  assign new_n34973_ = ~new_n34561_ & ~new_n34919_;
  assign new_n34974_ = ~new_n34918_ & new_n34973_;
  assign new_n34975_ = ~new_n34972_ & ~new_n34974_;
  assign new_n34976_ = ~\b[25]  & ~new_n34975_;
  assign new_n34977_ = ~new_n34580_ & new_n34878_;
  assign new_n34978_ = ~new_n34874_ & new_n34977_;
  assign new_n34979_ = ~new_n34875_ & ~new_n34878_;
  assign new_n34980_ = ~new_n34978_ & ~new_n34979_;
  assign new_n34981_ = ~new_n34920_ & ~new_n34980_;
  assign new_n34982_ = ~new_n34570_ & ~new_n34919_;
  assign new_n34983_ = ~new_n34918_ & new_n34982_;
  assign new_n34984_ = ~new_n34981_ & ~new_n34983_;
  assign new_n34985_ = ~\b[24]  & ~new_n34984_;
  assign new_n34986_ = ~new_n34589_ & new_n34873_;
  assign new_n34987_ = ~new_n34869_ & new_n34986_;
  assign new_n34988_ = ~new_n34870_ & ~new_n34873_;
  assign new_n34989_ = ~new_n34987_ & ~new_n34988_;
  assign new_n34990_ = ~new_n34920_ & ~new_n34989_;
  assign new_n34991_ = ~new_n34579_ & ~new_n34919_;
  assign new_n34992_ = ~new_n34918_ & new_n34991_;
  assign new_n34993_ = ~new_n34990_ & ~new_n34992_;
  assign new_n34994_ = ~\b[23]  & ~new_n34993_;
  assign new_n34995_ = ~new_n34598_ & new_n34868_;
  assign new_n34996_ = ~new_n34864_ & new_n34995_;
  assign new_n34997_ = ~new_n34865_ & ~new_n34868_;
  assign new_n34998_ = ~new_n34996_ & ~new_n34997_;
  assign new_n34999_ = ~new_n34920_ & ~new_n34998_;
  assign new_n35000_ = ~new_n34588_ & ~new_n34919_;
  assign new_n35001_ = ~new_n34918_ & new_n35000_;
  assign new_n35002_ = ~new_n34999_ & ~new_n35001_;
  assign new_n35003_ = ~\b[22]  & ~new_n35002_;
  assign new_n35004_ = ~new_n34607_ & new_n34863_;
  assign new_n35005_ = ~new_n34859_ & new_n35004_;
  assign new_n35006_ = ~new_n34860_ & ~new_n34863_;
  assign new_n35007_ = ~new_n35005_ & ~new_n35006_;
  assign new_n35008_ = ~new_n34920_ & ~new_n35007_;
  assign new_n35009_ = ~new_n34597_ & ~new_n34919_;
  assign new_n35010_ = ~new_n34918_ & new_n35009_;
  assign new_n35011_ = ~new_n35008_ & ~new_n35010_;
  assign new_n35012_ = ~\b[21]  & ~new_n35011_;
  assign new_n35013_ = ~new_n34616_ & new_n34858_;
  assign new_n35014_ = ~new_n34854_ & new_n35013_;
  assign new_n35015_ = ~new_n34855_ & ~new_n34858_;
  assign new_n35016_ = ~new_n35014_ & ~new_n35015_;
  assign new_n35017_ = ~new_n34920_ & ~new_n35016_;
  assign new_n35018_ = ~new_n34606_ & ~new_n34919_;
  assign new_n35019_ = ~new_n34918_ & new_n35018_;
  assign new_n35020_ = ~new_n35017_ & ~new_n35019_;
  assign new_n35021_ = ~\b[20]  & ~new_n35020_;
  assign new_n35022_ = ~new_n34625_ & new_n34853_;
  assign new_n35023_ = ~new_n34849_ & new_n35022_;
  assign new_n35024_ = ~new_n34850_ & ~new_n34853_;
  assign new_n35025_ = ~new_n35023_ & ~new_n35024_;
  assign new_n35026_ = ~new_n34920_ & ~new_n35025_;
  assign new_n35027_ = ~new_n34615_ & ~new_n34919_;
  assign new_n35028_ = ~new_n34918_ & new_n35027_;
  assign new_n35029_ = ~new_n35026_ & ~new_n35028_;
  assign new_n35030_ = ~\b[19]  & ~new_n35029_;
  assign new_n35031_ = ~new_n34634_ & new_n34848_;
  assign new_n35032_ = ~new_n34844_ & new_n35031_;
  assign new_n35033_ = ~new_n34845_ & ~new_n34848_;
  assign new_n35034_ = ~new_n35032_ & ~new_n35033_;
  assign new_n35035_ = ~new_n34920_ & ~new_n35034_;
  assign new_n35036_ = ~new_n34624_ & ~new_n34919_;
  assign new_n35037_ = ~new_n34918_ & new_n35036_;
  assign new_n35038_ = ~new_n35035_ & ~new_n35037_;
  assign new_n35039_ = ~\b[18]  & ~new_n35038_;
  assign new_n35040_ = ~new_n34643_ & new_n34843_;
  assign new_n35041_ = ~new_n34839_ & new_n35040_;
  assign new_n35042_ = ~new_n34840_ & ~new_n34843_;
  assign new_n35043_ = ~new_n35041_ & ~new_n35042_;
  assign new_n35044_ = ~new_n34920_ & ~new_n35043_;
  assign new_n35045_ = ~new_n34633_ & ~new_n34919_;
  assign new_n35046_ = ~new_n34918_ & new_n35045_;
  assign new_n35047_ = ~new_n35044_ & ~new_n35046_;
  assign new_n35048_ = ~\b[17]  & ~new_n35047_;
  assign new_n35049_ = ~new_n34652_ & new_n34838_;
  assign new_n35050_ = ~new_n34834_ & new_n35049_;
  assign new_n35051_ = ~new_n34835_ & ~new_n34838_;
  assign new_n35052_ = ~new_n35050_ & ~new_n35051_;
  assign new_n35053_ = ~new_n34920_ & ~new_n35052_;
  assign new_n35054_ = ~new_n34642_ & ~new_n34919_;
  assign new_n35055_ = ~new_n34918_ & new_n35054_;
  assign new_n35056_ = ~new_n35053_ & ~new_n35055_;
  assign new_n35057_ = ~\b[16]  & ~new_n35056_;
  assign new_n35058_ = ~new_n34661_ & new_n34833_;
  assign new_n35059_ = ~new_n34829_ & new_n35058_;
  assign new_n35060_ = ~new_n34830_ & ~new_n34833_;
  assign new_n35061_ = ~new_n35059_ & ~new_n35060_;
  assign new_n35062_ = ~new_n34920_ & ~new_n35061_;
  assign new_n35063_ = ~new_n34651_ & ~new_n34919_;
  assign new_n35064_ = ~new_n34918_ & new_n35063_;
  assign new_n35065_ = ~new_n35062_ & ~new_n35064_;
  assign new_n35066_ = ~\b[15]  & ~new_n35065_;
  assign new_n35067_ = ~new_n34670_ & new_n34828_;
  assign new_n35068_ = ~new_n34824_ & new_n35067_;
  assign new_n35069_ = ~new_n34825_ & ~new_n34828_;
  assign new_n35070_ = ~new_n35068_ & ~new_n35069_;
  assign new_n35071_ = ~new_n34920_ & ~new_n35070_;
  assign new_n35072_ = ~new_n34660_ & ~new_n34919_;
  assign new_n35073_ = ~new_n34918_ & new_n35072_;
  assign new_n35074_ = ~new_n35071_ & ~new_n35073_;
  assign new_n35075_ = ~\b[14]  & ~new_n35074_;
  assign new_n35076_ = ~new_n34679_ & new_n34823_;
  assign new_n35077_ = ~new_n34819_ & new_n35076_;
  assign new_n35078_ = ~new_n34820_ & ~new_n34823_;
  assign new_n35079_ = ~new_n35077_ & ~new_n35078_;
  assign new_n35080_ = ~new_n34920_ & ~new_n35079_;
  assign new_n35081_ = ~new_n34669_ & ~new_n34919_;
  assign new_n35082_ = ~new_n34918_ & new_n35081_;
  assign new_n35083_ = ~new_n35080_ & ~new_n35082_;
  assign new_n35084_ = ~\b[13]  & ~new_n35083_;
  assign new_n35085_ = ~new_n34688_ & new_n34818_;
  assign new_n35086_ = ~new_n34814_ & new_n35085_;
  assign new_n35087_ = ~new_n34815_ & ~new_n34818_;
  assign new_n35088_ = ~new_n35086_ & ~new_n35087_;
  assign new_n35089_ = ~new_n34920_ & ~new_n35088_;
  assign new_n35090_ = ~new_n34678_ & ~new_n34919_;
  assign new_n35091_ = ~new_n34918_ & new_n35090_;
  assign new_n35092_ = ~new_n35089_ & ~new_n35091_;
  assign new_n35093_ = ~\b[12]  & ~new_n35092_;
  assign new_n35094_ = ~new_n34697_ & new_n34813_;
  assign new_n35095_ = ~new_n34809_ & new_n35094_;
  assign new_n35096_ = ~new_n34810_ & ~new_n34813_;
  assign new_n35097_ = ~new_n35095_ & ~new_n35096_;
  assign new_n35098_ = ~new_n34920_ & ~new_n35097_;
  assign new_n35099_ = ~new_n34687_ & ~new_n34919_;
  assign new_n35100_ = ~new_n34918_ & new_n35099_;
  assign new_n35101_ = ~new_n35098_ & ~new_n35100_;
  assign new_n35102_ = ~\b[11]  & ~new_n35101_;
  assign new_n35103_ = ~new_n34706_ & new_n34808_;
  assign new_n35104_ = ~new_n34804_ & new_n35103_;
  assign new_n35105_ = ~new_n34805_ & ~new_n34808_;
  assign new_n35106_ = ~new_n35104_ & ~new_n35105_;
  assign new_n35107_ = ~new_n34920_ & ~new_n35106_;
  assign new_n35108_ = ~new_n34696_ & ~new_n34919_;
  assign new_n35109_ = ~new_n34918_ & new_n35108_;
  assign new_n35110_ = ~new_n35107_ & ~new_n35109_;
  assign new_n35111_ = ~\b[10]  & ~new_n35110_;
  assign new_n35112_ = ~new_n34715_ & new_n34803_;
  assign new_n35113_ = ~new_n34799_ & new_n35112_;
  assign new_n35114_ = ~new_n34800_ & ~new_n34803_;
  assign new_n35115_ = ~new_n35113_ & ~new_n35114_;
  assign new_n35116_ = ~new_n34920_ & ~new_n35115_;
  assign new_n35117_ = ~new_n34705_ & ~new_n34919_;
  assign new_n35118_ = ~new_n34918_ & new_n35117_;
  assign new_n35119_ = ~new_n35116_ & ~new_n35118_;
  assign new_n35120_ = ~\b[9]  & ~new_n35119_;
  assign new_n35121_ = ~new_n34724_ & new_n34798_;
  assign new_n35122_ = ~new_n34794_ & new_n35121_;
  assign new_n35123_ = ~new_n34795_ & ~new_n34798_;
  assign new_n35124_ = ~new_n35122_ & ~new_n35123_;
  assign new_n35125_ = ~new_n34920_ & ~new_n35124_;
  assign new_n35126_ = ~new_n34714_ & ~new_n34919_;
  assign new_n35127_ = ~new_n34918_ & new_n35126_;
  assign new_n35128_ = ~new_n35125_ & ~new_n35127_;
  assign new_n35129_ = ~\b[8]  & ~new_n35128_;
  assign new_n35130_ = ~new_n34733_ & new_n34793_;
  assign new_n35131_ = ~new_n34789_ & new_n35130_;
  assign new_n35132_ = ~new_n34790_ & ~new_n34793_;
  assign new_n35133_ = ~new_n35131_ & ~new_n35132_;
  assign new_n35134_ = ~new_n34920_ & ~new_n35133_;
  assign new_n35135_ = ~new_n34723_ & ~new_n34919_;
  assign new_n35136_ = ~new_n34918_ & new_n35135_;
  assign new_n35137_ = ~new_n35134_ & ~new_n35136_;
  assign new_n35138_ = ~\b[7]  & ~new_n35137_;
  assign new_n35139_ = ~new_n34742_ & new_n34788_;
  assign new_n35140_ = ~new_n34784_ & new_n35139_;
  assign new_n35141_ = ~new_n34785_ & ~new_n34788_;
  assign new_n35142_ = ~new_n35140_ & ~new_n35141_;
  assign new_n35143_ = ~new_n34920_ & ~new_n35142_;
  assign new_n35144_ = ~new_n34732_ & ~new_n34919_;
  assign new_n35145_ = ~new_n34918_ & new_n35144_;
  assign new_n35146_ = ~new_n35143_ & ~new_n35145_;
  assign new_n35147_ = ~\b[6]  & ~new_n35146_;
  assign new_n35148_ = ~new_n34751_ & new_n34783_;
  assign new_n35149_ = ~new_n34779_ & new_n35148_;
  assign new_n35150_ = ~new_n34780_ & ~new_n34783_;
  assign new_n35151_ = ~new_n35149_ & ~new_n35150_;
  assign new_n35152_ = ~new_n34920_ & ~new_n35151_;
  assign new_n35153_ = ~new_n34741_ & ~new_n34919_;
  assign new_n35154_ = ~new_n34918_ & new_n35153_;
  assign new_n35155_ = ~new_n35152_ & ~new_n35154_;
  assign new_n35156_ = ~\b[5]  & ~new_n35155_;
  assign new_n35157_ = ~new_n34759_ & new_n34778_;
  assign new_n35158_ = ~new_n34774_ & new_n35157_;
  assign new_n35159_ = ~new_n34775_ & ~new_n34778_;
  assign new_n35160_ = ~new_n35158_ & ~new_n35159_;
  assign new_n35161_ = ~new_n34920_ & ~new_n35160_;
  assign new_n35162_ = ~new_n34750_ & ~new_n34919_;
  assign new_n35163_ = ~new_n34918_ & new_n35162_;
  assign new_n35164_ = ~new_n35161_ & ~new_n35163_;
  assign new_n35165_ = ~\b[4]  & ~new_n35164_;
  assign new_n35166_ = ~new_n34769_ & new_n34773_;
  assign new_n35167_ = ~new_n34768_ & new_n35166_;
  assign new_n35168_ = ~new_n34770_ & ~new_n34773_;
  assign new_n35169_ = ~new_n35167_ & ~new_n35168_;
  assign new_n35170_ = ~new_n34920_ & ~new_n35169_;
  assign new_n35171_ = ~new_n34758_ & ~new_n34919_;
  assign new_n35172_ = ~new_n34918_ & new_n35171_;
  assign new_n35173_ = ~new_n35170_ & ~new_n35172_;
  assign new_n35174_ = ~\b[3]  & ~new_n35173_;
  assign new_n35175_ = new_n6584_ & ~new_n34766_;
  assign new_n35176_ = ~new_n34764_ & new_n35175_;
  assign new_n35177_ = ~new_n34768_ & ~new_n35176_;
  assign new_n35178_ = ~new_n34920_ & new_n35177_;
  assign new_n35179_ = ~new_n34763_ & ~new_n34919_;
  assign new_n35180_ = ~new_n34918_ & new_n35179_;
  assign new_n35181_ = ~new_n35178_ & ~new_n35180_;
  assign new_n35182_ = ~\b[2]  & ~new_n35181_;
  assign new_n35183_ = \b[0]  & ~new_n34920_;
  assign new_n35184_ = \a[34]  & ~new_n35183_;
  assign new_n35185_ = new_n6584_ & ~new_n34920_;
  assign new_n35186_ = ~new_n35184_ & ~new_n35185_;
  assign new_n35187_ = \b[1]  & ~new_n35186_;
  assign new_n35188_ = ~\b[1]  & ~new_n35185_;
  assign new_n35189_ = ~new_n35184_ & new_n35188_;
  assign new_n35190_ = ~new_n35187_ & ~new_n35189_;
  assign new_n35191_ = ~new_n7011_ & ~new_n35190_;
  assign new_n35192_ = ~\b[1]  & ~new_n35186_;
  assign new_n35193_ = ~new_n35191_ & ~new_n35192_;
  assign new_n35194_ = \b[2]  & ~new_n35180_;
  assign new_n35195_ = ~new_n35178_ & new_n35194_;
  assign new_n35196_ = ~new_n35182_ & ~new_n35195_;
  assign new_n35197_ = ~new_n35193_ & new_n35196_;
  assign new_n35198_ = ~new_n35182_ & ~new_n35197_;
  assign new_n35199_ = \b[3]  & ~new_n35172_;
  assign new_n35200_ = ~new_n35170_ & new_n35199_;
  assign new_n35201_ = ~new_n35174_ & ~new_n35200_;
  assign new_n35202_ = ~new_n35198_ & new_n35201_;
  assign new_n35203_ = ~new_n35174_ & ~new_n35202_;
  assign new_n35204_ = \b[4]  & ~new_n35163_;
  assign new_n35205_ = ~new_n35161_ & new_n35204_;
  assign new_n35206_ = ~new_n35165_ & ~new_n35205_;
  assign new_n35207_ = ~new_n35203_ & new_n35206_;
  assign new_n35208_ = ~new_n35165_ & ~new_n35207_;
  assign new_n35209_ = \b[5]  & ~new_n35154_;
  assign new_n35210_ = ~new_n35152_ & new_n35209_;
  assign new_n35211_ = ~new_n35156_ & ~new_n35210_;
  assign new_n35212_ = ~new_n35208_ & new_n35211_;
  assign new_n35213_ = ~new_n35156_ & ~new_n35212_;
  assign new_n35214_ = \b[6]  & ~new_n35145_;
  assign new_n35215_ = ~new_n35143_ & new_n35214_;
  assign new_n35216_ = ~new_n35147_ & ~new_n35215_;
  assign new_n35217_ = ~new_n35213_ & new_n35216_;
  assign new_n35218_ = ~new_n35147_ & ~new_n35217_;
  assign new_n35219_ = \b[7]  & ~new_n35136_;
  assign new_n35220_ = ~new_n35134_ & new_n35219_;
  assign new_n35221_ = ~new_n35138_ & ~new_n35220_;
  assign new_n35222_ = ~new_n35218_ & new_n35221_;
  assign new_n35223_ = ~new_n35138_ & ~new_n35222_;
  assign new_n35224_ = \b[8]  & ~new_n35127_;
  assign new_n35225_ = ~new_n35125_ & new_n35224_;
  assign new_n35226_ = ~new_n35129_ & ~new_n35225_;
  assign new_n35227_ = ~new_n35223_ & new_n35226_;
  assign new_n35228_ = ~new_n35129_ & ~new_n35227_;
  assign new_n35229_ = \b[9]  & ~new_n35118_;
  assign new_n35230_ = ~new_n35116_ & new_n35229_;
  assign new_n35231_ = ~new_n35120_ & ~new_n35230_;
  assign new_n35232_ = ~new_n35228_ & new_n35231_;
  assign new_n35233_ = ~new_n35120_ & ~new_n35232_;
  assign new_n35234_ = \b[10]  & ~new_n35109_;
  assign new_n35235_ = ~new_n35107_ & new_n35234_;
  assign new_n35236_ = ~new_n35111_ & ~new_n35235_;
  assign new_n35237_ = ~new_n35233_ & new_n35236_;
  assign new_n35238_ = ~new_n35111_ & ~new_n35237_;
  assign new_n35239_ = \b[11]  & ~new_n35100_;
  assign new_n35240_ = ~new_n35098_ & new_n35239_;
  assign new_n35241_ = ~new_n35102_ & ~new_n35240_;
  assign new_n35242_ = ~new_n35238_ & new_n35241_;
  assign new_n35243_ = ~new_n35102_ & ~new_n35242_;
  assign new_n35244_ = \b[12]  & ~new_n35091_;
  assign new_n35245_ = ~new_n35089_ & new_n35244_;
  assign new_n35246_ = ~new_n35093_ & ~new_n35245_;
  assign new_n35247_ = ~new_n35243_ & new_n35246_;
  assign new_n35248_ = ~new_n35093_ & ~new_n35247_;
  assign new_n35249_ = \b[13]  & ~new_n35082_;
  assign new_n35250_ = ~new_n35080_ & new_n35249_;
  assign new_n35251_ = ~new_n35084_ & ~new_n35250_;
  assign new_n35252_ = ~new_n35248_ & new_n35251_;
  assign new_n35253_ = ~new_n35084_ & ~new_n35252_;
  assign new_n35254_ = \b[14]  & ~new_n35073_;
  assign new_n35255_ = ~new_n35071_ & new_n35254_;
  assign new_n35256_ = ~new_n35075_ & ~new_n35255_;
  assign new_n35257_ = ~new_n35253_ & new_n35256_;
  assign new_n35258_ = ~new_n35075_ & ~new_n35257_;
  assign new_n35259_ = \b[15]  & ~new_n35064_;
  assign new_n35260_ = ~new_n35062_ & new_n35259_;
  assign new_n35261_ = ~new_n35066_ & ~new_n35260_;
  assign new_n35262_ = ~new_n35258_ & new_n35261_;
  assign new_n35263_ = ~new_n35066_ & ~new_n35262_;
  assign new_n35264_ = \b[16]  & ~new_n35055_;
  assign new_n35265_ = ~new_n35053_ & new_n35264_;
  assign new_n35266_ = ~new_n35057_ & ~new_n35265_;
  assign new_n35267_ = ~new_n35263_ & new_n35266_;
  assign new_n35268_ = ~new_n35057_ & ~new_n35267_;
  assign new_n35269_ = \b[17]  & ~new_n35046_;
  assign new_n35270_ = ~new_n35044_ & new_n35269_;
  assign new_n35271_ = ~new_n35048_ & ~new_n35270_;
  assign new_n35272_ = ~new_n35268_ & new_n35271_;
  assign new_n35273_ = ~new_n35048_ & ~new_n35272_;
  assign new_n35274_ = \b[18]  & ~new_n35037_;
  assign new_n35275_ = ~new_n35035_ & new_n35274_;
  assign new_n35276_ = ~new_n35039_ & ~new_n35275_;
  assign new_n35277_ = ~new_n35273_ & new_n35276_;
  assign new_n35278_ = ~new_n35039_ & ~new_n35277_;
  assign new_n35279_ = \b[19]  & ~new_n35028_;
  assign new_n35280_ = ~new_n35026_ & new_n35279_;
  assign new_n35281_ = ~new_n35030_ & ~new_n35280_;
  assign new_n35282_ = ~new_n35278_ & new_n35281_;
  assign new_n35283_ = ~new_n35030_ & ~new_n35282_;
  assign new_n35284_ = \b[20]  & ~new_n35019_;
  assign new_n35285_ = ~new_n35017_ & new_n35284_;
  assign new_n35286_ = ~new_n35021_ & ~new_n35285_;
  assign new_n35287_ = ~new_n35283_ & new_n35286_;
  assign new_n35288_ = ~new_n35021_ & ~new_n35287_;
  assign new_n35289_ = \b[21]  & ~new_n35010_;
  assign new_n35290_ = ~new_n35008_ & new_n35289_;
  assign new_n35291_ = ~new_n35012_ & ~new_n35290_;
  assign new_n35292_ = ~new_n35288_ & new_n35291_;
  assign new_n35293_ = ~new_n35012_ & ~new_n35292_;
  assign new_n35294_ = \b[22]  & ~new_n35001_;
  assign new_n35295_ = ~new_n34999_ & new_n35294_;
  assign new_n35296_ = ~new_n35003_ & ~new_n35295_;
  assign new_n35297_ = ~new_n35293_ & new_n35296_;
  assign new_n35298_ = ~new_n35003_ & ~new_n35297_;
  assign new_n35299_ = \b[23]  & ~new_n34992_;
  assign new_n35300_ = ~new_n34990_ & new_n35299_;
  assign new_n35301_ = ~new_n34994_ & ~new_n35300_;
  assign new_n35302_ = ~new_n35298_ & new_n35301_;
  assign new_n35303_ = ~new_n34994_ & ~new_n35302_;
  assign new_n35304_ = \b[24]  & ~new_n34983_;
  assign new_n35305_ = ~new_n34981_ & new_n35304_;
  assign new_n35306_ = ~new_n34985_ & ~new_n35305_;
  assign new_n35307_ = ~new_n35303_ & new_n35306_;
  assign new_n35308_ = ~new_n34985_ & ~new_n35307_;
  assign new_n35309_ = \b[25]  & ~new_n34974_;
  assign new_n35310_ = ~new_n34972_ & new_n35309_;
  assign new_n35311_ = ~new_n34976_ & ~new_n35310_;
  assign new_n35312_ = ~new_n35308_ & new_n35311_;
  assign new_n35313_ = ~new_n34976_ & ~new_n35312_;
  assign new_n35314_ = \b[26]  & ~new_n34965_;
  assign new_n35315_ = ~new_n34963_ & new_n35314_;
  assign new_n35316_ = ~new_n34967_ & ~new_n35315_;
  assign new_n35317_ = ~new_n35313_ & new_n35316_;
  assign new_n35318_ = ~new_n34967_ & ~new_n35317_;
  assign new_n35319_ = \b[27]  & ~new_n34956_;
  assign new_n35320_ = ~new_n34954_ & new_n35319_;
  assign new_n35321_ = ~new_n34958_ & ~new_n35320_;
  assign new_n35322_ = ~new_n35318_ & new_n35321_;
  assign new_n35323_ = ~new_n34958_ & ~new_n35322_;
  assign new_n35324_ = \b[28]  & ~new_n34947_;
  assign new_n35325_ = ~new_n34945_ & new_n35324_;
  assign new_n35326_ = ~new_n34949_ & ~new_n35325_;
  assign new_n35327_ = ~new_n35323_ & new_n35326_;
  assign new_n35328_ = ~new_n34949_ & ~new_n35327_;
  assign new_n35329_ = \b[29]  & ~new_n34927_;
  assign new_n35330_ = ~new_n34925_ & new_n35329_;
  assign new_n35331_ = ~new_n34940_ & ~new_n35330_;
  assign new_n35332_ = ~new_n35328_ & new_n35331_;
  assign new_n35333_ = ~new_n34940_ & ~new_n35332_;
  assign new_n35334_ = \b[30]  & ~new_n34937_;
  assign new_n35335_ = ~new_n34935_ & new_n35334_;
  assign new_n35336_ = ~new_n34939_ & ~new_n35335_;
  assign new_n35337_ = ~new_n35333_ & new_n35336_;
  assign new_n35338_ = ~new_n34939_ & ~new_n35337_;
  assign new_n35339_ = new_n7162_ & ~new_n35338_;
  assign new_n35340_ = ~new_n34928_ & ~new_n35339_;
  assign new_n35341_ = ~new_n34949_ & new_n35331_;
  assign new_n35342_ = ~new_n35327_ & new_n35341_;
  assign new_n35343_ = ~new_n35328_ & ~new_n35331_;
  assign new_n35344_ = ~new_n35342_ & ~new_n35343_;
  assign new_n35345_ = new_n7162_ & ~new_n35344_;
  assign new_n35346_ = ~new_n35338_ & new_n35345_;
  assign new_n35347_ = ~new_n35340_ & ~new_n35346_;
  assign new_n35348_ = ~new_n34938_ & ~new_n35339_;
  assign new_n35349_ = ~new_n34940_ & new_n35336_;
  assign new_n35350_ = ~new_n35332_ & new_n35349_;
  assign new_n35351_ = ~new_n35333_ & ~new_n35336_;
  assign new_n35352_ = ~new_n35350_ & ~new_n35351_;
  assign new_n35353_ = new_n35339_ & ~new_n35352_;
  assign new_n35354_ = ~new_n35348_ & ~new_n35353_;
  assign new_n35355_ = ~\b[31]  & ~new_n35354_;
  assign new_n35356_ = ~\b[30]  & ~new_n35347_;
  assign new_n35357_ = ~new_n34948_ & ~new_n35339_;
  assign new_n35358_ = ~new_n34958_ & new_n35326_;
  assign new_n35359_ = ~new_n35322_ & new_n35358_;
  assign new_n35360_ = ~new_n35323_ & ~new_n35326_;
  assign new_n35361_ = ~new_n35359_ & ~new_n35360_;
  assign new_n35362_ = new_n7162_ & ~new_n35361_;
  assign new_n35363_ = ~new_n35338_ & new_n35362_;
  assign new_n35364_ = ~new_n35357_ & ~new_n35363_;
  assign new_n35365_ = ~\b[29]  & ~new_n35364_;
  assign new_n35366_ = ~new_n34957_ & ~new_n35339_;
  assign new_n35367_ = ~new_n34967_ & new_n35321_;
  assign new_n35368_ = ~new_n35317_ & new_n35367_;
  assign new_n35369_ = ~new_n35318_ & ~new_n35321_;
  assign new_n35370_ = ~new_n35368_ & ~new_n35369_;
  assign new_n35371_ = new_n7162_ & ~new_n35370_;
  assign new_n35372_ = ~new_n35338_ & new_n35371_;
  assign new_n35373_ = ~new_n35366_ & ~new_n35372_;
  assign new_n35374_ = ~\b[28]  & ~new_n35373_;
  assign new_n35375_ = ~new_n34966_ & ~new_n35339_;
  assign new_n35376_ = ~new_n34976_ & new_n35316_;
  assign new_n35377_ = ~new_n35312_ & new_n35376_;
  assign new_n35378_ = ~new_n35313_ & ~new_n35316_;
  assign new_n35379_ = ~new_n35377_ & ~new_n35378_;
  assign new_n35380_ = new_n7162_ & ~new_n35379_;
  assign new_n35381_ = ~new_n35338_ & new_n35380_;
  assign new_n35382_ = ~new_n35375_ & ~new_n35381_;
  assign new_n35383_ = ~\b[27]  & ~new_n35382_;
  assign new_n35384_ = ~new_n34975_ & ~new_n35339_;
  assign new_n35385_ = ~new_n34985_ & new_n35311_;
  assign new_n35386_ = ~new_n35307_ & new_n35385_;
  assign new_n35387_ = ~new_n35308_ & ~new_n35311_;
  assign new_n35388_ = ~new_n35386_ & ~new_n35387_;
  assign new_n35389_ = new_n7162_ & ~new_n35388_;
  assign new_n35390_ = ~new_n35338_ & new_n35389_;
  assign new_n35391_ = ~new_n35384_ & ~new_n35390_;
  assign new_n35392_ = ~\b[26]  & ~new_n35391_;
  assign new_n35393_ = ~new_n34984_ & ~new_n35339_;
  assign new_n35394_ = ~new_n34994_ & new_n35306_;
  assign new_n35395_ = ~new_n35302_ & new_n35394_;
  assign new_n35396_ = ~new_n35303_ & ~new_n35306_;
  assign new_n35397_ = ~new_n35395_ & ~new_n35396_;
  assign new_n35398_ = new_n7162_ & ~new_n35397_;
  assign new_n35399_ = ~new_n35338_ & new_n35398_;
  assign new_n35400_ = ~new_n35393_ & ~new_n35399_;
  assign new_n35401_ = ~\b[25]  & ~new_n35400_;
  assign new_n35402_ = ~new_n34993_ & ~new_n35339_;
  assign new_n35403_ = ~new_n35003_ & new_n35301_;
  assign new_n35404_ = ~new_n35297_ & new_n35403_;
  assign new_n35405_ = ~new_n35298_ & ~new_n35301_;
  assign new_n35406_ = ~new_n35404_ & ~new_n35405_;
  assign new_n35407_ = new_n7162_ & ~new_n35406_;
  assign new_n35408_ = ~new_n35338_ & new_n35407_;
  assign new_n35409_ = ~new_n35402_ & ~new_n35408_;
  assign new_n35410_ = ~\b[24]  & ~new_n35409_;
  assign new_n35411_ = ~new_n35002_ & ~new_n35339_;
  assign new_n35412_ = ~new_n35012_ & new_n35296_;
  assign new_n35413_ = ~new_n35292_ & new_n35412_;
  assign new_n35414_ = ~new_n35293_ & ~new_n35296_;
  assign new_n35415_ = ~new_n35413_ & ~new_n35414_;
  assign new_n35416_ = new_n7162_ & ~new_n35415_;
  assign new_n35417_ = ~new_n35338_ & new_n35416_;
  assign new_n35418_ = ~new_n35411_ & ~new_n35417_;
  assign new_n35419_ = ~\b[23]  & ~new_n35418_;
  assign new_n35420_ = ~new_n35011_ & ~new_n35339_;
  assign new_n35421_ = ~new_n35021_ & new_n35291_;
  assign new_n35422_ = ~new_n35287_ & new_n35421_;
  assign new_n35423_ = ~new_n35288_ & ~new_n35291_;
  assign new_n35424_ = ~new_n35422_ & ~new_n35423_;
  assign new_n35425_ = new_n7162_ & ~new_n35424_;
  assign new_n35426_ = ~new_n35338_ & new_n35425_;
  assign new_n35427_ = ~new_n35420_ & ~new_n35426_;
  assign new_n35428_ = ~\b[22]  & ~new_n35427_;
  assign new_n35429_ = ~new_n35020_ & ~new_n35339_;
  assign new_n35430_ = ~new_n35030_ & new_n35286_;
  assign new_n35431_ = ~new_n35282_ & new_n35430_;
  assign new_n35432_ = ~new_n35283_ & ~new_n35286_;
  assign new_n35433_ = ~new_n35431_ & ~new_n35432_;
  assign new_n35434_ = new_n7162_ & ~new_n35433_;
  assign new_n35435_ = ~new_n35338_ & new_n35434_;
  assign new_n35436_ = ~new_n35429_ & ~new_n35435_;
  assign new_n35437_ = ~\b[21]  & ~new_n35436_;
  assign new_n35438_ = ~new_n35029_ & ~new_n35339_;
  assign new_n35439_ = ~new_n35039_ & new_n35281_;
  assign new_n35440_ = ~new_n35277_ & new_n35439_;
  assign new_n35441_ = ~new_n35278_ & ~new_n35281_;
  assign new_n35442_ = ~new_n35440_ & ~new_n35441_;
  assign new_n35443_ = new_n7162_ & ~new_n35442_;
  assign new_n35444_ = ~new_n35338_ & new_n35443_;
  assign new_n35445_ = ~new_n35438_ & ~new_n35444_;
  assign new_n35446_ = ~\b[20]  & ~new_n35445_;
  assign new_n35447_ = ~new_n35038_ & ~new_n35339_;
  assign new_n35448_ = ~new_n35048_ & new_n35276_;
  assign new_n35449_ = ~new_n35272_ & new_n35448_;
  assign new_n35450_ = ~new_n35273_ & ~new_n35276_;
  assign new_n35451_ = ~new_n35449_ & ~new_n35450_;
  assign new_n35452_ = new_n7162_ & ~new_n35451_;
  assign new_n35453_ = ~new_n35338_ & new_n35452_;
  assign new_n35454_ = ~new_n35447_ & ~new_n35453_;
  assign new_n35455_ = ~\b[19]  & ~new_n35454_;
  assign new_n35456_ = ~new_n35047_ & ~new_n35339_;
  assign new_n35457_ = ~new_n35057_ & new_n35271_;
  assign new_n35458_ = ~new_n35267_ & new_n35457_;
  assign new_n35459_ = ~new_n35268_ & ~new_n35271_;
  assign new_n35460_ = ~new_n35458_ & ~new_n35459_;
  assign new_n35461_ = new_n7162_ & ~new_n35460_;
  assign new_n35462_ = ~new_n35338_ & new_n35461_;
  assign new_n35463_ = ~new_n35456_ & ~new_n35462_;
  assign new_n35464_ = ~\b[18]  & ~new_n35463_;
  assign new_n35465_ = ~new_n35056_ & ~new_n35339_;
  assign new_n35466_ = ~new_n35066_ & new_n35266_;
  assign new_n35467_ = ~new_n35262_ & new_n35466_;
  assign new_n35468_ = ~new_n35263_ & ~new_n35266_;
  assign new_n35469_ = ~new_n35467_ & ~new_n35468_;
  assign new_n35470_ = new_n7162_ & ~new_n35469_;
  assign new_n35471_ = ~new_n35338_ & new_n35470_;
  assign new_n35472_ = ~new_n35465_ & ~new_n35471_;
  assign new_n35473_ = ~\b[17]  & ~new_n35472_;
  assign new_n35474_ = ~new_n35065_ & ~new_n35339_;
  assign new_n35475_ = ~new_n35075_ & new_n35261_;
  assign new_n35476_ = ~new_n35257_ & new_n35475_;
  assign new_n35477_ = ~new_n35258_ & ~new_n35261_;
  assign new_n35478_ = ~new_n35476_ & ~new_n35477_;
  assign new_n35479_ = new_n7162_ & ~new_n35478_;
  assign new_n35480_ = ~new_n35338_ & new_n35479_;
  assign new_n35481_ = ~new_n35474_ & ~new_n35480_;
  assign new_n35482_ = ~\b[16]  & ~new_n35481_;
  assign new_n35483_ = ~new_n35074_ & ~new_n35339_;
  assign new_n35484_ = ~new_n35084_ & new_n35256_;
  assign new_n35485_ = ~new_n35252_ & new_n35484_;
  assign new_n35486_ = ~new_n35253_ & ~new_n35256_;
  assign new_n35487_ = ~new_n35485_ & ~new_n35486_;
  assign new_n35488_ = new_n7162_ & ~new_n35487_;
  assign new_n35489_ = ~new_n35338_ & new_n35488_;
  assign new_n35490_ = ~new_n35483_ & ~new_n35489_;
  assign new_n35491_ = ~\b[15]  & ~new_n35490_;
  assign new_n35492_ = ~new_n35083_ & ~new_n35339_;
  assign new_n35493_ = ~new_n35093_ & new_n35251_;
  assign new_n35494_ = ~new_n35247_ & new_n35493_;
  assign new_n35495_ = ~new_n35248_ & ~new_n35251_;
  assign new_n35496_ = ~new_n35494_ & ~new_n35495_;
  assign new_n35497_ = new_n7162_ & ~new_n35496_;
  assign new_n35498_ = ~new_n35338_ & new_n35497_;
  assign new_n35499_ = ~new_n35492_ & ~new_n35498_;
  assign new_n35500_ = ~\b[14]  & ~new_n35499_;
  assign new_n35501_ = ~new_n35092_ & ~new_n35339_;
  assign new_n35502_ = ~new_n35102_ & new_n35246_;
  assign new_n35503_ = ~new_n35242_ & new_n35502_;
  assign new_n35504_ = ~new_n35243_ & ~new_n35246_;
  assign new_n35505_ = ~new_n35503_ & ~new_n35504_;
  assign new_n35506_ = new_n7162_ & ~new_n35505_;
  assign new_n35507_ = ~new_n35338_ & new_n35506_;
  assign new_n35508_ = ~new_n35501_ & ~new_n35507_;
  assign new_n35509_ = ~\b[13]  & ~new_n35508_;
  assign new_n35510_ = ~new_n35101_ & ~new_n35339_;
  assign new_n35511_ = ~new_n35111_ & new_n35241_;
  assign new_n35512_ = ~new_n35237_ & new_n35511_;
  assign new_n35513_ = ~new_n35238_ & ~new_n35241_;
  assign new_n35514_ = ~new_n35512_ & ~new_n35513_;
  assign new_n35515_ = new_n7162_ & ~new_n35514_;
  assign new_n35516_ = ~new_n35338_ & new_n35515_;
  assign new_n35517_ = ~new_n35510_ & ~new_n35516_;
  assign new_n35518_ = ~\b[12]  & ~new_n35517_;
  assign new_n35519_ = ~new_n35110_ & ~new_n35339_;
  assign new_n35520_ = ~new_n35120_ & new_n35236_;
  assign new_n35521_ = ~new_n35232_ & new_n35520_;
  assign new_n35522_ = ~new_n35233_ & ~new_n35236_;
  assign new_n35523_ = ~new_n35521_ & ~new_n35522_;
  assign new_n35524_ = new_n7162_ & ~new_n35523_;
  assign new_n35525_ = ~new_n35338_ & new_n35524_;
  assign new_n35526_ = ~new_n35519_ & ~new_n35525_;
  assign new_n35527_ = ~\b[11]  & ~new_n35526_;
  assign new_n35528_ = ~new_n35119_ & ~new_n35339_;
  assign new_n35529_ = ~new_n35129_ & new_n35231_;
  assign new_n35530_ = ~new_n35227_ & new_n35529_;
  assign new_n35531_ = ~new_n35228_ & ~new_n35231_;
  assign new_n35532_ = ~new_n35530_ & ~new_n35531_;
  assign new_n35533_ = new_n7162_ & ~new_n35532_;
  assign new_n35534_ = ~new_n35338_ & new_n35533_;
  assign new_n35535_ = ~new_n35528_ & ~new_n35534_;
  assign new_n35536_ = ~\b[10]  & ~new_n35535_;
  assign new_n35537_ = ~new_n35128_ & ~new_n35339_;
  assign new_n35538_ = ~new_n35138_ & new_n35226_;
  assign new_n35539_ = ~new_n35222_ & new_n35538_;
  assign new_n35540_ = ~new_n35223_ & ~new_n35226_;
  assign new_n35541_ = ~new_n35539_ & ~new_n35540_;
  assign new_n35542_ = new_n7162_ & ~new_n35541_;
  assign new_n35543_ = ~new_n35338_ & new_n35542_;
  assign new_n35544_ = ~new_n35537_ & ~new_n35543_;
  assign new_n35545_ = ~\b[9]  & ~new_n35544_;
  assign new_n35546_ = ~new_n35137_ & ~new_n35339_;
  assign new_n35547_ = ~new_n35147_ & new_n35221_;
  assign new_n35548_ = ~new_n35217_ & new_n35547_;
  assign new_n35549_ = ~new_n35218_ & ~new_n35221_;
  assign new_n35550_ = ~new_n35548_ & ~new_n35549_;
  assign new_n35551_ = new_n7162_ & ~new_n35550_;
  assign new_n35552_ = ~new_n35338_ & new_n35551_;
  assign new_n35553_ = ~new_n35546_ & ~new_n35552_;
  assign new_n35554_ = ~\b[8]  & ~new_n35553_;
  assign new_n35555_ = ~new_n35146_ & ~new_n35339_;
  assign new_n35556_ = ~new_n35156_ & new_n35216_;
  assign new_n35557_ = ~new_n35212_ & new_n35556_;
  assign new_n35558_ = ~new_n35213_ & ~new_n35216_;
  assign new_n35559_ = ~new_n35557_ & ~new_n35558_;
  assign new_n35560_ = new_n7162_ & ~new_n35559_;
  assign new_n35561_ = ~new_n35338_ & new_n35560_;
  assign new_n35562_ = ~new_n35555_ & ~new_n35561_;
  assign new_n35563_ = ~\b[7]  & ~new_n35562_;
  assign new_n35564_ = ~new_n35155_ & ~new_n35339_;
  assign new_n35565_ = ~new_n35165_ & new_n35211_;
  assign new_n35566_ = ~new_n35207_ & new_n35565_;
  assign new_n35567_ = ~new_n35208_ & ~new_n35211_;
  assign new_n35568_ = ~new_n35566_ & ~new_n35567_;
  assign new_n35569_ = new_n7162_ & ~new_n35568_;
  assign new_n35570_ = ~new_n35338_ & new_n35569_;
  assign new_n35571_ = ~new_n35564_ & ~new_n35570_;
  assign new_n35572_ = ~\b[6]  & ~new_n35571_;
  assign new_n35573_ = ~new_n35164_ & ~new_n35339_;
  assign new_n35574_ = ~new_n35174_ & new_n35206_;
  assign new_n35575_ = ~new_n35202_ & new_n35574_;
  assign new_n35576_ = ~new_n35203_ & ~new_n35206_;
  assign new_n35577_ = ~new_n35575_ & ~new_n35576_;
  assign new_n35578_ = new_n7162_ & ~new_n35577_;
  assign new_n35579_ = ~new_n35338_ & new_n35578_;
  assign new_n35580_ = ~new_n35573_ & ~new_n35579_;
  assign new_n35581_ = ~\b[5]  & ~new_n35580_;
  assign new_n35582_ = ~new_n35173_ & ~new_n35339_;
  assign new_n35583_ = ~new_n35182_ & new_n35201_;
  assign new_n35584_ = ~new_n35197_ & new_n35583_;
  assign new_n35585_ = ~new_n35198_ & ~new_n35201_;
  assign new_n35586_ = ~new_n35584_ & ~new_n35585_;
  assign new_n35587_ = new_n7162_ & ~new_n35586_;
  assign new_n35588_ = ~new_n35338_ & new_n35587_;
  assign new_n35589_ = ~new_n35582_ & ~new_n35588_;
  assign new_n35590_ = ~\b[4]  & ~new_n35589_;
  assign new_n35591_ = ~new_n35181_ & ~new_n35339_;
  assign new_n35592_ = ~new_n35192_ & new_n35196_;
  assign new_n35593_ = ~new_n35191_ & new_n35592_;
  assign new_n35594_ = ~new_n35193_ & ~new_n35196_;
  assign new_n35595_ = ~new_n35593_ & ~new_n35594_;
  assign new_n35596_ = new_n7162_ & ~new_n35595_;
  assign new_n35597_ = ~new_n35338_ & new_n35596_;
  assign new_n35598_ = ~new_n35591_ & ~new_n35597_;
  assign new_n35599_ = ~\b[3]  & ~new_n35598_;
  assign new_n35600_ = ~new_n35186_ & ~new_n35339_;
  assign new_n35601_ = new_n7011_ & ~new_n35189_;
  assign new_n35602_ = ~new_n35187_ & new_n35601_;
  assign new_n35603_ = new_n7162_ & ~new_n35602_;
  assign new_n35604_ = ~new_n35191_ & new_n35603_;
  assign new_n35605_ = ~new_n35338_ & new_n35604_;
  assign new_n35606_ = ~new_n35600_ & ~new_n35605_;
  assign new_n35607_ = ~\b[2]  & ~new_n35606_;
  assign new_n35608_ = new_n7435_ & ~new_n35338_;
  assign new_n35609_ = \a[33]  & ~new_n35608_;
  assign new_n35610_ = new_n7441_ & ~new_n35338_;
  assign new_n35611_ = ~new_n35609_ & ~new_n35610_;
  assign new_n35612_ = \b[1]  & ~new_n35611_;
  assign new_n35613_ = ~\b[1]  & ~new_n35610_;
  assign new_n35614_ = ~new_n35609_ & new_n35613_;
  assign new_n35615_ = ~new_n35612_ & ~new_n35614_;
  assign new_n35616_ = ~new_n7448_ & ~new_n35615_;
  assign new_n35617_ = ~\b[1]  & ~new_n35611_;
  assign new_n35618_ = ~new_n35616_ & ~new_n35617_;
  assign new_n35619_ = \b[2]  & ~new_n35605_;
  assign new_n35620_ = ~new_n35600_ & new_n35619_;
  assign new_n35621_ = ~new_n35607_ & ~new_n35620_;
  assign new_n35622_ = ~new_n35618_ & new_n35621_;
  assign new_n35623_ = ~new_n35607_ & ~new_n35622_;
  assign new_n35624_ = \b[3]  & ~new_n35597_;
  assign new_n35625_ = ~new_n35591_ & new_n35624_;
  assign new_n35626_ = ~new_n35599_ & ~new_n35625_;
  assign new_n35627_ = ~new_n35623_ & new_n35626_;
  assign new_n35628_ = ~new_n35599_ & ~new_n35627_;
  assign new_n35629_ = \b[4]  & ~new_n35588_;
  assign new_n35630_ = ~new_n35582_ & new_n35629_;
  assign new_n35631_ = ~new_n35590_ & ~new_n35630_;
  assign new_n35632_ = ~new_n35628_ & new_n35631_;
  assign new_n35633_ = ~new_n35590_ & ~new_n35632_;
  assign new_n35634_ = \b[5]  & ~new_n35579_;
  assign new_n35635_ = ~new_n35573_ & new_n35634_;
  assign new_n35636_ = ~new_n35581_ & ~new_n35635_;
  assign new_n35637_ = ~new_n35633_ & new_n35636_;
  assign new_n35638_ = ~new_n35581_ & ~new_n35637_;
  assign new_n35639_ = \b[6]  & ~new_n35570_;
  assign new_n35640_ = ~new_n35564_ & new_n35639_;
  assign new_n35641_ = ~new_n35572_ & ~new_n35640_;
  assign new_n35642_ = ~new_n35638_ & new_n35641_;
  assign new_n35643_ = ~new_n35572_ & ~new_n35642_;
  assign new_n35644_ = \b[7]  & ~new_n35561_;
  assign new_n35645_ = ~new_n35555_ & new_n35644_;
  assign new_n35646_ = ~new_n35563_ & ~new_n35645_;
  assign new_n35647_ = ~new_n35643_ & new_n35646_;
  assign new_n35648_ = ~new_n35563_ & ~new_n35647_;
  assign new_n35649_ = \b[8]  & ~new_n35552_;
  assign new_n35650_ = ~new_n35546_ & new_n35649_;
  assign new_n35651_ = ~new_n35554_ & ~new_n35650_;
  assign new_n35652_ = ~new_n35648_ & new_n35651_;
  assign new_n35653_ = ~new_n35554_ & ~new_n35652_;
  assign new_n35654_ = \b[9]  & ~new_n35543_;
  assign new_n35655_ = ~new_n35537_ & new_n35654_;
  assign new_n35656_ = ~new_n35545_ & ~new_n35655_;
  assign new_n35657_ = ~new_n35653_ & new_n35656_;
  assign new_n35658_ = ~new_n35545_ & ~new_n35657_;
  assign new_n35659_ = \b[10]  & ~new_n35534_;
  assign new_n35660_ = ~new_n35528_ & new_n35659_;
  assign new_n35661_ = ~new_n35536_ & ~new_n35660_;
  assign new_n35662_ = ~new_n35658_ & new_n35661_;
  assign new_n35663_ = ~new_n35536_ & ~new_n35662_;
  assign new_n35664_ = \b[11]  & ~new_n35525_;
  assign new_n35665_ = ~new_n35519_ & new_n35664_;
  assign new_n35666_ = ~new_n35527_ & ~new_n35665_;
  assign new_n35667_ = ~new_n35663_ & new_n35666_;
  assign new_n35668_ = ~new_n35527_ & ~new_n35667_;
  assign new_n35669_ = \b[12]  & ~new_n35516_;
  assign new_n35670_ = ~new_n35510_ & new_n35669_;
  assign new_n35671_ = ~new_n35518_ & ~new_n35670_;
  assign new_n35672_ = ~new_n35668_ & new_n35671_;
  assign new_n35673_ = ~new_n35518_ & ~new_n35672_;
  assign new_n35674_ = \b[13]  & ~new_n35507_;
  assign new_n35675_ = ~new_n35501_ & new_n35674_;
  assign new_n35676_ = ~new_n35509_ & ~new_n35675_;
  assign new_n35677_ = ~new_n35673_ & new_n35676_;
  assign new_n35678_ = ~new_n35509_ & ~new_n35677_;
  assign new_n35679_ = \b[14]  & ~new_n35498_;
  assign new_n35680_ = ~new_n35492_ & new_n35679_;
  assign new_n35681_ = ~new_n35500_ & ~new_n35680_;
  assign new_n35682_ = ~new_n35678_ & new_n35681_;
  assign new_n35683_ = ~new_n35500_ & ~new_n35682_;
  assign new_n35684_ = \b[15]  & ~new_n35489_;
  assign new_n35685_ = ~new_n35483_ & new_n35684_;
  assign new_n35686_ = ~new_n35491_ & ~new_n35685_;
  assign new_n35687_ = ~new_n35683_ & new_n35686_;
  assign new_n35688_ = ~new_n35491_ & ~new_n35687_;
  assign new_n35689_ = \b[16]  & ~new_n35480_;
  assign new_n35690_ = ~new_n35474_ & new_n35689_;
  assign new_n35691_ = ~new_n35482_ & ~new_n35690_;
  assign new_n35692_ = ~new_n35688_ & new_n35691_;
  assign new_n35693_ = ~new_n35482_ & ~new_n35692_;
  assign new_n35694_ = \b[17]  & ~new_n35471_;
  assign new_n35695_ = ~new_n35465_ & new_n35694_;
  assign new_n35696_ = ~new_n35473_ & ~new_n35695_;
  assign new_n35697_ = ~new_n35693_ & new_n35696_;
  assign new_n35698_ = ~new_n35473_ & ~new_n35697_;
  assign new_n35699_ = \b[18]  & ~new_n35462_;
  assign new_n35700_ = ~new_n35456_ & new_n35699_;
  assign new_n35701_ = ~new_n35464_ & ~new_n35700_;
  assign new_n35702_ = ~new_n35698_ & new_n35701_;
  assign new_n35703_ = ~new_n35464_ & ~new_n35702_;
  assign new_n35704_ = \b[19]  & ~new_n35453_;
  assign new_n35705_ = ~new_n35447_ & new_n35704_;
  assign new_n35706_ = ~new_n35455_ & ~new_n35705_;
  assign new_n35707_ = ~new_n35703_ & new_n35706_;
  assign new_n35708_ = ~new_n35455_ & ~new_n35707_;
  assign new_n35709_ = \b[20]  & ~new_n35444_;
  assign new_n35710_ = ~new_n35438_ & new_n35709_;
  assign new_n35711_ = ~new_n35446_ & ~new_n35710_;
  assign new_n35712_ = ~new_n35708_ & new_n35711_;
  assign new_n35713_ = ~new_n35446_ & ~new_n35712_;
  assign new_n35714_ = \b[21]  & ~new_n35435_;
  assign new_n35715_ = ~new_n35429_ & new_n35714_;
  assign new_n35716_ = ~new_n35437_ & ~new_n35715_;
  assign new_n35717_ = ~new_n35713_ & new_n35716_;
  assign new_n35718_ = ~new_n35437_ & ~new_n35717_;
  assign new_n35719_ = \b[22]  & ~new_n35426_;
  assign new_n35720_ = ~new_n35420_ & new_n35719_;
  assign new_n35721_ = ~new_n35428_ & ~new_n35720_;
  assign new_n35722_ = ~new_n35718_ & new_n35721_;
  assign new_n35723_ = ~new_n35428_ & ~new_n35722_;
  assign new_n35724_ = \b[23]  & ~new_n35417_;
  assign new_n35725_ = ~new_n35411_ & new_n35724_;
  assign new_n35726_ = ~new_n35419_ & ~new_n35725_;
  assign new_n35727_ = ~new_n35723_ & new_n35726_;
  assign new_n35728_ = ~new_n35419_ & ~new_n35727_;
  assign new_n35729_ = \b[24]  & ~new_n35408_;
  assign new_n35730_ = ~new_n35402_ & new_n35729_;
  assign new_n35731_ = ~new_n35410_ & ~new_n35730_;
  assign new_n35732_ = ~new_n35728_ & new_n35731_;
  assign new_n35733_ = ~new_n35410_ & ~new_n35732_;
  assign new_n35734_ = \b[25]  & ~new_n35399_;
  assign new_n35735_ = ~new_n35393_ & new_n35734_;
  assign new_n35736_ = ~new_n35401_ & ~new_n35735_;
  assign new_n35737_ = ~new_n35733_ & new_n35736_;
  assign new_n35738_ = ~new_n35401_ & ~new_n35737_;
  assign new_n35739_ = \b[26]  & ~new_n35390_;
  assign new_n35740_ = ~new_n35384_ & new_n35739_;
  assign new_n35741_ = ~new_n35392_ & ~new_n35740_;
  assign new_n35742_ = ~new_n35738_ & new_n35741_;
  assign new_n35743_ = ~new_n35392_ & ~new_n35742_;
  assign new_n35744_ = \b[27]  & ~new_n35381_;
  assign new_n35745_ = ~new_n35375_ & new_n35744_;
  assign new_n35746_ = ~new_n35383_ & ~new_n35745_;
  assign new_n35747_ = ~new_n35743_ & new_n35746_;
  assign new_n35748_ = ~new_n35383_ & ~new_n35747_;
  assign new_n35749_ = \b[28]  & ~new_n35372_;
  assign new_n35750_ = ~new_n35366_ & new_n35749_;
  assign new_n35751_ = ~new_n35374_ & ~new_n35750_;
  assign new_n35752_ = ~new_n35748_ & new_n35751_;
  assign new_n35753_ = ~new_n35374_ & ~new_n35752_;
  assign new_n35754_ = \b[29]  & ~new_n35363_;
  assign new_n35755_ = ~new_n35357_ & new_n35754_;
  assign new_n35756_ = ~new_n35365_ & ~new_n35755_;
  assign new_n35757_ = ~new_n35753_ & new_n35756_;
  assign new_n35758_ = ~new_n35365_ & ~new_n35757_;
  assign new_n35759_ = \b[30]  & ~new_n35346_;
  assign new_n35760_ = ~new_n35340_ & new_n35759_;
  assign new_n35761_ = ~new_n35356_ & ~new_n35760_;
  assign new_n35762_ = ~new_n35758_ & new_n35761_;
  assign new_n35763_ = ~new_n35356_ & ~new_n35762_;
  assign new_n35764_ = \b[31]  & ~new_n35348_;
  assign new_n35765_ = ~new_n35353_ & new_n35764_;
  assign new_n35766_ = ~new_n35355_ & ~new_n35765_;
  assign new_n35767_ = ~new_n35763_ & new_n35766_;
  assign new_n35768_ = ~new_n35355_ & ~new_n35767_;
  assign new_n35769_ = new_n432_ & ~new_n35768_;
  assign new_n35770_ = ~new_n35347_ & ~new_n35769_;
  assign new_n35771_ = ~new_n35365_ & new_n35761_;
  assign new_n35772_ = ~new_n35757_ & new_n35771_;
  assign new_n35773_ = ~new_n35758_ & ~new_n35761_;
  assign new_n35774_ = ~new_n35772_ & ~new_n35773_;
  assign new_n35775_ = new_n432_ & ~new_n35774_;
  assign new_n35776_ = ~new_n35768_ & new_n35775_;
  assign new_n35777_ = ~new_n35770_ & ~new_n35776_;
  assign new_n35778_ = ~\b[31]  & ~new_n35777_;
  assign new_n35779_ = ~new_n35364_ & ~new_n35769_;
  assign new_n35780_ = ~new_n35374_ & new_n35756_;
  assign new_n35781_ = ~new_n35752_ & new_n35780_;
  assign new_n35782_ = ~new_n35753_ & ~new_n35756_;
  assign new_n35783_ = ~new_n35781_ & ~new_n35782_;
  assign new_n35784_ = new_n432_ & ~new_n35783_;
  assign new_n35785_ = ~new_n35768_ & new_n35784_;
  assign new_n35786_ = ~new_n35779_ & ~new_n35785_;
  assign new_n35787_ = ~\b[30]  & ~new_n35786_;
  assign new_n35788_ = ~new_n35373_ & ~new_n35769_;
  assign new_n35789_ = ~new_n35383_ & new_n35751_;
  assign new_n35790_ = ~new_n35747_ & new_n35789_;
  assign new_n35791_ = ~new_n35748_ & ~new_n35751_;
  assign new_n35792_ = ~new_n35790_ & ~new_n35791_;
  assign new_n35793_ = new_n432_ & ~new_n35792_;
  assign new_n35794_ = ~new_n35768_ & new_n35793_;
  assign new_n35795_ = ~new_n35788_ & ~new_n35794_;
  assign new_n35796_ = ~\b[29]  & ~new_n35795_;
  assign new_n35797_ = ~new_n35382_ & ~new_n35769_;
  assign new_n35798_ = ~new_n35392_ & new_n35746_;
  assign new_n35799_ = ~new_n35742_ & new_n35798_;
  assign new_n35800_ = ~new_n35743_ & ~new_n35746_;
  assign new_n35801_ = ~new_n35799_ & ~new_n35800_;
  assign new_n35802_ = new_n432_ & ~new_n35801_;
  assign new_n35803_ = ~new_n35768_ & new_n35802_;
  assign new_n35804_ = ~new_n35797_ & ~new_n35803_;
  assign new_n35805_ = ~\b[28]  & ~new_n35804_;
  assign new_n35806_ = ~new_n35391_ & ~new_n35769_;
  assign new_n35807_ = ~new_n35401_ & new_n35741_;
  assign new_n35808_ = ~new_n35737_ & new_n35807_;
  assign new_n35809_ = ~new_n35738_ & ~new_n35741_;
  assign new_n35810_ = ~new_n35808_ & ~new_n35809_;
  assign new_n35811_ = new_n432_ & ~new_n35810_;
  assign new_n35812_ = ~new_n35768_ & new_n35811_;
  assign new_n35813_ = ~new_n35806_ & ~new_n35812_;
  assign new_n35814_ = ~\b[27]  & ~new_n35813_;
  assign new_n35815_ = ~new_n35400_ & ~new_n35769_;
  assign new_n35816_ = ~new_n35410_ & new_n35736_;
  assign new_n35817_ = ~new_n35732_ & new_n35816_;
  assign new_n35818_ = ~new_n35733_ & ~new_n35736_;
  assign new_n35819_ = ~new_n35817_ & ~new_n35818_;
  assign new_n35820_ = new_n432_ & ~new_n35819_;
  assign new_n35821_ = ~new_n35768_ & new_n35820_;
  assign new_n35822_ = ~new_n35815_ & ~new_n35821_;
  assign new_n35823_ = ~\b[26]  & ~new_n35822_;
  assign new_n35824_ = ~new_n35409_ & ~new_n35769_;
  assign new_n35825_ = ~new_n35419_ & new_n35731_;
  assign new_n35826_ = ~new_n35727_ & new_n35825_;
  assign new_n35827_ = ~new_n35728_ & ~new_n35731_;
  assign new_n35828_ = ~new_n35826_ & ~new_n35827_;
  assign new_n35829_ = new_n432_ & ~new_n35828_;
  assign new_n35830_ = ~new_n35768_ & new_n35829_;
  assign new_n35831_ = ~new_n35824_ & ~new_n35830_;
  assign new_n35832_ = ~\b[25]  & ~new_n35831_;
  assign new_n35833_ = ~new_n35418_ & ~new_n35769_;
  assign new_n35834_ = ~new_n35428_ & new_n35726_;
  assign new_n35835_ = ~new_n35722_ & new_n35834_;
  assign new_n35836_ = ~new_n35723_ & ~new_n35726_;
  assign new_n35837_ = ~new_n35835_ & ~new_n35836_;
  assign new_n35838_ = new_n432_ & ~new_n35837_;
  assign new_n35839_ = ~new_n35768_ & new_n35838_;
  assign new_n35840_ = ~new_n35833_ & ~new_n35839_;
  assign new_n35841_ = ~\b[24]  & ~new_n35840_;
  assign new_n35842_ = ~new_n35427_ & ~new_n35769_;
  assign new_n35843_ = ~new_n35437_ & new_n35721_;
  assign new_n35844_ = ~new_n35717_ & new_n35843_;
  assign new_n35845_ = ~new_n35718_ & ~new_n35721_;
  assign new_n35846_ = ~new_n35844_ & ~new_n35845_;
  assign new_n35847_ = new_n432_ & ~new_n35846_;
  assign new_n35848_ = ~new_n35768_ & new_n35847_;
  assign new_n35849_ = ~new_n35842_ & ~new_n35848_;
  assign new_n35850_ = ~\b[23]  & ~new_n35849_;
  assign new_n35851_ = ~new_n35436_ & ~new_n35769_;
  assign new_n35852_ = ~new_n35446_ & new_n35716_;
  assign new_n35853_ = ~new_n35712_ & new_n35852_;
  assign new_n35854_ = ~new_n35713_ & ~new_n35716_;
  assign new_n35855_ = ~new_n35853_ & ~new_n35854_;
  assign new_n35856_ = new_n432_ & ~new_n35855_;
  assign new_n35857_ = ~new_n35768_ & new_n35856_;
  assign new_n35858_ = ~new_n35851_ & ~new_n35857_;
  assign new_n35859_ = ~\b[22]  & ~new_n35858_;
  assign new_n35860_ = ~new_n35445_ & ~new_n35769_;
  assign new_n35861_ = ~new_n35455_ & new_n35711_;
  assign new_n35862_ = ~new_n35707_ & new_n35861_;
  assign new_n35863_ = ~new_n35708_ & ~new_n35711_;
  assign new_n35864_ = ~new_n35862_ & ~new_n35863_;
  assign new_n35865_ = new_n432_ & ~new_n35864_;
  assign new_n35866_ = ~new_n35768_ & new_n35865_;
  assign new_n35867_ = ~new_n35860_ & ~new_n35866_;
  assign new_n35868_ = ~\b[21]  & ~new_n35867_;
  assign new_n35869_ = ~new_n35454_ & ~new_n35769_;
  assign new_n35870_ = ~new_n35464_ & new_n35706_;
  assign new_n35871_ = ~new_n35702_ & new_n35870_;
  assign new_n35872_ = ~new_n35703_ & ~new_n35706_;
  assign new_n35873_ = ~new_n35871_ & ~new_n35872_;
  assign new_n35874_ = new_n432_ & ~new_n35873_;
  assign new_n35875_ = ~new_n35768_ & new_n35874_;
  assign new_n35876_ = ~new_n35869_ & ~new_n35875_;
  assign new_n35877_ = ~\b[20]  & ~new_n35876_;
  assign new_n35878_ = ~new_n35463_ & ~new_n35769_;
  assign new_n35879_ = ~new_n35473_ & new_n35701_;
  assign new_n35880_ = ~new_n35697_ & new_n35879_;
  assign new_n35881_ = ~new_n35698_ & ~new_n35701_;
  assign new_n35882_ = ~new_n35880_ & ~new_n35881_;
  assign new_n35883_ = new_n432_ & ~new_n35882_;
  assign new_n35884_ = ~new_n35768_ & new_n35883_;
  assign new_n35885_ = ~new_n35878_ & ~new_n35884_;
  assign new_n35886_ = ~\b[19]  & ~new_n35885_;
  assign new_n35887_ = ~new_n35472_ & ~new_n35769_;
  assign new_n35888_ = ~new_n35482_ & new_n35696_;
  assign new_n35889_ = ~new_n35692_ & new_n35888_;
  assign new_n35890_ = ~new_n35693_ & ~new_n35696_;
  assign new_n35891_ = ~new_n35889_ & ~new_n35890_;
  assign new_n35892_ = new_n432_ & ~new_n35891_;
  assign new_n35893_ = ~new_n35768_ & new_n35892_;
  assign new_n35894_ = ~new_n35887_ & ~new_n35893_;
  assign new_n35895_ = ~\b[18]  & ~new_n35894_;
  assign new_n35896_ = ~new_n35481_ & ~new_n35769_;
  assign new_n35897_ = ~new_n35491_ & new_n35691_;
  assign new_n35898_ = ~new_n35687_ & new_n35897_;
  assign new_n35899_ = ~new_n35688_ & ~new_n35691_;
  assign new_n35900_ = ~new_n35898_ & ~new_n35899_;
  assign new_n35901_ = new_n432_ & ~new_n35900_;
  assign new_n35902_ = ~new_n35768_ & new_n35901_;
  assign new_n35903_ = ~new_n35896_ & ~new_n35902_;
  assign new_n35904_ = ~\b[17]  & ~new_n35903_;
  assign new_n35905_ = ~new_n35490_ & ~new_n35769_;
  assign new_n35906_ = ~new_n35500_ & new_n35686_;
  assign new_n35907_ = ~new_n35682_ & new_n35906_;
  assign new_n35908_ = ~new_n35683_ & ~new_n35686_;
  assign new_n35909_ = ~new_n35907_ & ~new_n35908_;
  assign new_n35910_ = new_n432_ & ~new_n35909_;
  assign new_n35911_ = ~new_n35768_ & new_n35910_;
  assign new_n35912_ = ~new_n35905_ & ~new_n35911_;
  assign new_n35913_ = ~\b[16]  & ~new_n35912_;
  assign new_n35914_ = ~new_n35499_ & ~new_n35769_;
  assign new_n35915_ = ~new_n35509_ & new_n35681_;
  assign new_n35916_ = ~new_n35677_ & new_n35915_;
  assign new_n35917_ = ~new_n35678_ & ~new_n35681_;
  assign new_n35918_ = ~new_n35916_ & ~new_n35917_;
  assign new_n35919_ = new_n432_ & ~new_n35918_;
  assign new_n35920_ = ~new_n35768_ & new_n35919_;
  assign new_n35921_ = ~new_n35914_ & ~new_n35920_;
  assign new_n35922_ = ~\b[15]  & ~new_n35921_;
  assign new_n35923_ = ~new_n35508_ & ~new_n35769_;
  assign new_n35924_ = ~new_n35518_ & new_n35676_;
  assign new_n35925_ = ~new_n35672_ & new_n35924_;
  assign new_n35926_ = ~new_n35673_ & ~new_n35676_;
  assign new_n35927_ = ~new_n35925_ & ~new_n35926_;
  assign new_n35928_ = new_n432_ & ~new_n35927_;
  assign new_n35929_ = ~new_n35768_ & new_n35928_;
  assign new_n35930_ = ~new_n35923_ & ~new_n35929_;
  assign new_n35931_ = ~\b[14]  & ~new_n35930_;
  assign new_n35932_ = ~new_n35517_ & ~new_n35769_;
  assign new_n35933_ = ~new_n35527_ & new_n35671_;
  assign new_n35934_ = ~new_n35667_ & new_n35933_;
  assign new_n35935_ = ~new_n35668_ & ~new_n35671_;
  assign new_n35936_ = ~new_n35934_ & ~new_n35935_;
  assign new_n35937_ = new_n432_ & ~new_n35936_;
  assign new_n35938_ = ~new_n35768_ & new_n35937_;
  assign new_n35939_ = ~new_n35932_ & ~new_n35938_;
  assign new_n35940_ = ~\b[13]  & ~new_n35939_;
  assign new_n35941_ = ~new_n35526_ & ~new_n35769_;
  assign new_n35942_ = ~new_n35536_ & new_n35666_;
  assign new_n35943_ = ~new_n35662_ & new_n35942_;
  assign new_n35944_ = ~new_n35663_ & ~new_n35666_;
  assign new_n35945_ = ~new_n35943_ & ~new_n35944_;
  assign new_n35946_ = new_n432_ & ~new_n35945_;
  assign new_n35947_ = ~new_n35768_ & new_n35946_;
  assign new_n35948_ = ~new_n35941_ & ~new_n35947_;
  assign new_n35949_ = ~\b[12]  & ~new_n35948_;
  assign new_n35950_ = ~new_n35535_ & ~new_n35769_;
  assign new_n35951_ = ~new_n35545_ & new_n35661_;
  assign new_n35952_ = ~new_n35657_ & new_n35951_;
  assign new_n35953_ = ~new_n35658_ & ~new_n35661_;
  assign new_n35954_ = ~new_n35952_ & ~new_n35953_;
  assign new_n35955_ = new_n432_ & ~new_n35954_;
  assign new_n35956_ = ~new_n35768_ & new_n35955_;
  assign new_n35957_ = ~new_n35950_ & ~new_n35956_;
  assign new_n35958_ = ~\b[11]  & ~new_n35957_;
  assign new_n35959_ = ~new_n35544_ & ~new_n35769_;
  assign new_n35960_ = ~new_n35554_ & new_n35656_;
  assign new_n35961_ = ~new_n35652_ & new_n35960_;
  assign new_n35962_ = ~new_n35653_ & ~new_n35656_;
  assign new_n35963_ = ~new_n35961_ & ~new_n35962_;
  assign new_n35964_ = new_n432_ & ~new_n35963_;
  assign new_n35965_ = ~new_n35768_ & new_n35964_;
  assign new_n35966_ = ~new_n35959_ & ~new_n35965_;
  assign new_n35967_ = ~\b[10]  & ~new_n35966_;
  assign new_n35968_ = ~new_n35553_ & ~new_n35769_;
  assign new_n35969_ = ~new_n35563_ & new_n35651_;
  assign new_n35970_ = ~new_n35647_ & new_n35969_;
  assign new_n35971_ = ~new_n35648_ & ~new_n35651_;
  assign new_n35972_ = ~new_n35970_ & ~new_n35971_;
  assign new_n35973_ = new_n432_ & ~new_n35972_;
  assign new_n35974_ = ~new_n35768_ & new_n35973_;
  assign new_n35975_ = ~new_n35968_ & ~new_n35974_;
  assign new_n35976_ = ~\b[9]  & ~new_n35975_;
  assign new_n35977_ = ~new_n35562_ & ~new_n35769_;
  assign new_n35978_ = ~new_n35572_ & new_n35646_;
  assign new_n35979_ = ~new_n35642_ & new_n35978_;
  assign new_n35980_ = ~new_n35643_ & ~new_n35646_;
  assign new_n35981_ = ~new_n35979_ & ~new_n35980_;
  assign new_n35982_ = new_n432_ & ~new_n35981_;
  assign new_n35983_ = ~new_n35768_ & new_n35982_;
  assign new_n35984_ = ~new_n35977_ & ~new_n35983_;
  assign new_n35985_ = ~\b[8]  & ~new_n35984_;
  assign new_n35986_ = ~new_n35571_ & ~new_n35769_;
  assign new_n35987_ = ~new_n35581_ & new_n35641_;
  assign new_n35988_ = ~new_n35637_ & new_n35987_;
  assign new_n35989_ = ~new_n35638_ & ~new_n35641_;
  assign new_n35990_ = ~new_n35988_ & ~new_n35989_;
  assign new_n35991_ = new_n432_ & ~new_n35990_;
  assign new_n35992_ = ~new_n35768_ & new_n35991_;
  assign new_n35993_ = ~new_n35986_ & ~new_n35992_;
  assign new_n35994_ = ~\b[7]  & ~new_n35993_;
  assign new_n35995_ = ~new_n35580_ & ~new_n35769_;
  assign new_n35996_ = ~new_n35590_ & new_n35636_;
  assign new_n35997_ = ~new_n35632_ & new_n35996_;
  assign new_n35998_ = ~new_n35633_ & ~new_n35636_;
  assign new_n35999_ = ~new_n35997_ & ~new_n35998_;
  assign new_n36000_ = new_n432_ & ~new_n35999_;
  assign new_n36001_ = ~new_n35768_ & new_n36000_;
  assign new_n36002_ = ~new_n35995_ & ~new_n36001_;
  assign new_n36003_ = ~\b[6]  & ~new_n36002_;
  assign new_n36004_ = ~new_n35589_ & ~new_n35769_;
  assign new_n36005_ = ~new_n35599_ & new_n35631_;
  assign new_n36006_ = ~new_n35627_ & new_n36005_;
  assign new_n36007_ = ~new_n35628_ & ~new_n35631_;
  assign new_n36008_ = ~new_n36006_ & ~new_n36007_;
  assign new_n36009_ = new_n432_ & ~new_n36008_;
  assign new_n36010_ = ~new_n35768_ & new_n36009_;
  assign new_n36011_ = ~new_n36004_ & ~new_n36010_;
  assign new_n36012_ = ~\b[5]  & ~new_n36011_;
  assign new_n36013_ = ~new_n35598_ & ~new_n35769_;
  assign new_n36014_ = ~new_n35607_ & new_n35626_;
  assign new_n36015_ = ~new_n35622_ & new_n36014_;
  assign new_n36016_ = ~new_n35623_ & ~new_n35626_;
  assign new_n36017_ = ~new_n36015_ & ~new_n36016_;
  assign new_n36018_ = new_n432_ & ~new_n36017_;
  assign new_n36019_ = ~new_n35768_ & new_n36018_;
  assign new_n36020_ = ~new_n36013_ & ~new_n36019_;
  assign new_n36021_ = ~\b[4]  & ~new_n36020_;
  assign new_n36022_ = ~new_n35606_ & ~new_n35769_;
  assign new_n36023_ = ~new_n35617_ & new_n35621_;
  assign new_n36024_ = ~new_n35616_ & new_n36023_;
  assign new_n36025_ = ~new_n35618_ & ~new_n35621_;
  assign new_n36026_ = ~new_n36024_ & ~new_n36025_;
  assign new_n36027_ = new_n432_ & ~new_n36026_;
  assign new_n36028_ = ~new_n35768_ & new_n36027_;
  assign new_n36029_ = ~new_n36022_ & ~new_n36028_;
  assign new_n36030_ = ~\b[3]  & ~new_n36029_;
  assign new_n36031_ = ~new_n35611_ & ~new_n35769_;
  assign new_n36032_ = new_n7448_ & ~new_n35614_;
  assign new_n36033_ = ~new_n35612_ & new_n36032_;
  assign new_n36034_ = new_n432_ & ~new_n36033_;
  assign new_n36035_ = ~new_n35616_ & new_n36034_;
  assign new_n36036_ = ~new_n35768_ & new_n36035_;
  assign new_n36037_ = ~new_n36031_ & ~new_n36036_;
  assign new_n36038_ = ~\b[2]  & ~new_n36037_;
  assign new_n36039_ = new_n7875_ & ~new_n35768_;
  assign new_n36040_ = \a[32]  & ~new_n36039_;
  assign new_n36041_ = new_n7880_ & ~new_n35768_;
  assign new_n36042_ = ~new_n36040_ & ~new_n36041_;
  assign new_n36043_ = \b[1]  & ~new_n36042_;
  assign new_n36044_ = ~\b[1]  & ~new_n36041_;
  assign new_n36045_ = ~new_n36040_ & new_n36044_;
  assign new_n36046_ = ~new_n36043_ & ~new_n36045_;
  assign new_n36047_ = ~new_n7887_ & ~new_n36046_;
  assign new_n36048_ = ~\b[1]  & ~new_n36042_;
  assign new_n36049_ = ~new_n36047_ & ~new_n36048_;
  assign new_n36050_ = \b[2]  & ~new_n36036_;
  assign new_n36051_ = ~new_n36031_ & new_n36050_;
  assign new_n36052_ = ~new_n36038_ & ~new_n36051_;
  assign new_n36053_ = ~new_n36049_ & new_n36052_;
  assign new_n36054_ = ~new_n36038_ & ~new_n36053_;
  assign new_n36055_ = \b[3]  & ~new_n36028_;
  assign new_n36056_ = ~new_n36022_ & new_n36055_;
  assign new_n36057_ = ~new_n36030_ & ~new_n36056_;
  assign new_n36058_ = ~new_n36054_ & new_n36057_;
  assign new_n36059_ = ~new_n36030_ & ~new_n36058_;
  assign new_n36060_ = \b[4]  & ~new_n36019_;
  assign new_n36061_ = ~new_n36013_ & new_n36060_;
  assign new_n36062_ = ~new_n36021_ & ~new_n36061_;
  assign new_n36063_ = ~new_n36059_ & new_n36062_;
  assign new_n36064_ = ~new_n36021_ & ~new_n36063_;
  assign new_n36065_ = \b[5]  & ~new_n36010_;
  assign new_n36066_ = ~new_n36004_ & new_n36065_;
  assign new_n36067_ = ~new_n36012_ & ~new_n36066_;
  assign new_n36068_ = ~new_n36064_ & new_n36067_;
  assign new_n36069_ = ~new_n36012_ & ~new_n36068_;
  assign new_n36070_ = \b[6]  & ~new_n36001_;
  assign new_n36071_ = ~new_n35995_ & new_n36070_;
  assign new_n36072_ = ~new_n36003_ & ~new_n36071_;
  assign new_n36073_ = ~new_n36069_ & new_n36072_;
  assign new_n36074_ = ~new_n36003_ & ~new_n36073_;
  assign new_n36075_ = \b[7]  & ~new_n35992_;
  assign new_n36076_ = ~new_n35986_ & new_n36075_;
  assign new_n36077_ = ~new_n35994_ & ~new_n36076_;
  assign new_n36078_ = ~new_n36074_ & new_n36077_;
  assign new_n36079_ = ~new_n35994_ & ~new_n36078_;
  assign new_n36080_ = \b[8]  & ~new_n35983_;
  assign new_n36081_ = ~new_n35977_ & new_n36080_;
  assign new_n36082_ = ~new_n35985_ & ~new_n36081_;
  assign new_n36083_ = ~new_n36079_ & new_n36082_;
  assign new_n36084_ = ~new_n35985_ & ~new_n36083_;
  assign new_n36085_ = \b[9]  & ~new_n35974_;
  assign new_n36086_ = ~new_n35968_ & new_n36085_;
  assign new_n36087_ = ~new_n35976_ & ~new_n36086_;
  assign new_n36088_ = ~new_n36084_ & new_n36087_;
  assign new_n36089_ = ~new_n35976_ & ~new_n36088_;
  assign new_n36090_ = \b[10]  & ~new_n35965_;
  assign new_n36091_ = ~new_n35959_ & new_n36090_;
  assign new_n36092_ = ~new_n35967_ & ~new_n36091_;
  assign new_n36093_ = ~new_n36089_ & new_n36092_;
  assign new_n36094_ = ~new_n35967_ & ~new_n36093_;
  assign new_n36095_ = \b[11]  & ~new_n35956_;
  assign new_n36096_ = ~new_n35950_ & new_n36095_;
  assign new_n36097_ = ~new_n35958_ & ~new_n36096_;
  assign new_n36098_ = ~new_n36094_ & new_n36097_;
  assign new_n36099_ = ~new_n35958_ & ~new_n36098_;
  assign new_n36100_ = \b[12]  & ~new_n35947_;
  assign new_n36101_ = ~new_n35941_ & new_n36100_;
  assign new_n36102_ = ~new_n35949_ & ~new_n36101_;
  assign new_n36103_ = ~new_n36099_ & new_n36102_;
  assign new_n36104_ = ~new_n35949_ & ~new_n36103_;
  assign new_n36105_ = \b[13]  & ~new_n35938_;
  assign new_n36106_ = ~new_n35932_ & new_n36105_;
  assign new_n36107_ = ~new_n35940_ & ~new_n36106_;
  assign new_n36108_ = ~new_n36104_ & new_n36107_;
  assign new_n36109_ = ~new_n35940_ & ~new_n36108_;
  assign new_n36110_ = \b[14]  & ~new_n35929_;
  assign new_n36111_ = ~new_n35923_ & new_n36110_;
  assign new_n36112_ = ~new_n35931_ & ~new_n36111_;
  assign new_n36113_ = ~new_n36109_ & new_n36112_;
  assign new_n36114_ = ~new_n35931_ & ~new_n36113_;
  assign new_n36115_ = \b[15]  & ~new_n35920_;
  assign new_n36116_ = ~new_n35914_ & new_n36115_;
  assign new_n36117_ = ~new_n35922_ & ~new_n36116_;
  assign new_n36118_ = ~new_n36114_ & new_n36117_;
  assign new_n36119_ = ~new_n35922_ & ~new_n36118_;
  assign new_n36120_ = \b[16]  & ~new_n35911_;
  assign new_n36121_ = ~new_n35905_ & new_n36120_;
  assign new_n36122_ = ~new_n35913_ & ~new_n36121_;
  assign new_n36123_ = ~new_n36119_ & new_n36122_;
  assign new_n36124_ = ~new_n35913_ & ~new_n36123_;
  assign new_n36125_ = \b[17]  & ~new_n35902_;
  assign new_n36126_ = ~new_n35896_ & new_n36125_;
  assign new_n36127_ = ~new_n35904_ & ~new_n36126_;
  assign new_n36128_ = ~new_n36124_ & new_n36127_;
  assign new_n36129_ = ~new_n35904_ & ~new_n36128_;
  assign new_n36130_ = \b[18]  & ~new_n35893_;
  assign new_n36131_ = ~new_n35887_ & new_n36130_;
  assign new_n36132_ = ~new_n35895_ & ~new_n36131_;
  assign new_n36133_ = ~new_n36129_ & new_n36132_;
  assign new_n36134_ = ~new_n35895_ & ~new_n36133_;
  assign new_n36135_ = \b[19]  & ~new_n35884_;
  assign new_n36136_ = ~new_n35878_ & new_n36135_;
  assign new_n36137_ = ~new_n35886_ & ~new_n36136_;
  assign new_n36138_ = ~new_n36134_ & new_n36137_;
  assign new_n36139_ = ~new_n35886_ & ~new_n36138_;
  assign new_n36140_ = \b[20]  & ~new_n35875_;
  assign new_n36141_ = ~new_n35869_ & new_n36140_;
  assign new_n36142_ = ~new_n35877_ & ~new_n36141_;
  assign new_n36143_ = ~new_n36139_ & new_n36142_;
  assign new_n36144_ = ~new_n35877_ & ~new_n36143_;
  assign new_n36145_ = \b[21]  & ~new_n35866_;
  assign new_n36146_ = ~new_n35860_ & new_n36145_;
  assign new_n36147_ = ~new_n35868_ & ~new_n36146_;
  assign new_n36148_ = ~new_n36144_ & new_n36147_;
  assign new_n36149_ = ~new_n35868_ & ~new_n36148_;
  assign new_n36150_ = \b[22]  & ~new_n35857_;
  assign new_n36151_ = ~new_n35851_ & new_n36150_;
  assign new_n36152_ = ~new_n35859_ & ~new_n36151_;
  assign new_n36153_ = ~new_n36149_ & new_n36152_;
  assign new_n36154_ = ~new_n35859_ & ~new_n36153_;
  assign new_n36155_ = \b[23]  & ~new_n35848_;
  assign new_n36156_ = ~new_n35842_ & new_n36155_;
  assign new_n36157_ = ~new_n35850_ & ~new_n36156_;
  assign new_n36158_ = ~new_n36154_ & new_n36157_;
  assign new_n36159_ = ~new_n35850_ & ~new_n36158_;
  assign new_n36160_ = \b[24]  & ~new_n35839_;
  assign new_n36161_ = ~new_n35833_ & new_n36160_;
  assign new_n36162_ = ~new_n35841_ & ~new_n36161_;
  assign new_n36163_ = ~new_n36159_ & new_n36162_;
  assign new_n36164_ = ~new_n35841_ & ~new_n36163_;
  assign new_n36165_ = \b[25]  & ~new_n35830_;
  assign new_n36166_ = ~new_n35824_ & new_n36165_;
  assign new_n36167_ = ~new_n35832_ & ~new_n36166_;
  assign new_n36168_ = ~new_n36164_ & new_n36167_;
  assign new_n36169_ = ~new_n35832_ & ~new_n36168_;
  assign new_n36170_ = \b[26]  & ~new_n35821_;
  assign new_n36171_ = ~new_n35815_ & new_n36170_;
  assign new_n36172_ = ~new_n35823_ & ~new_n36171_;
  assign new_n36173_ = ~new_n36169_ & new_n36172_;
  assign new_n36174_ = ~new_n35823_ & ~new_n36173_;
  assign new_n36175_ = \b[27]  & ~new_n35812_;
  assign new_n36176_ = ~new_n35806_ & new_n36175_;
  assign new_n36177_ = ~new_n35814_ & ~new_n36176_;
  assign new_n36178_ = ~new_n36174_ & new_n36177_;
  assign new_n36179_ = ~new_n35814_ & ~new_n36178_;
  assign new_n36180_ = \b[28]  & ~new_n35803_;
  assign new_n36181_ = ~new_n35797_ & new_n36180_;
  assign new_n36182_ = ~new_n35805_ & ~new_n36181_;
  assign new_n36183_ = ~new_n36179_ & new_n36182_;
  assign new_n36184_ = ~new_n35805_ & ~new_n36183_;
  assign new_n36185_ = \b[29]  & ~new_n35794_;
  assign new_n36186_ = ~new_n35788_ & new_n36185_;
  assign new_n36187_ = ~new_n35796_ & ~new_n36186_;
  assign new_n36188_ = ~new_n36184_ & new_n36187_;
  assign new_n36189_ = ~new_n35796_ & ~new_n36188_;
  assign new_n36190_ = \b[30]  & ~new_n35785_;
  assign new_n36191_ = ~new_n35779_ & new_n36190_;
  assign new_n36192_ = ~new_n35787_ & ~new_n36191_;
  assign new_n36193_ = ~new_n36189_ & new_n36192_;
  assign new_n36194_ = ~new_n35787_ & ~new_n36193_;
  assign new_n36195_ = \b[31]  & ~new_n35776_;
  assign new_n36196_ = ~new_n35770_ & new_n36195_;
  assign new_n36197_ = ~new_n35778_ & ~new_n36196_;
  assign new_n36198_ = ~new_n36194_ & new_n36197_;
  assign new_n36199_ = ~new_n35778_ & ~new_n36198_;
  assign new_n36200_ = ~new_n35354_ & ~new_n35769_;
  assign new_n36201_ = ~new_n35356_ & new_n35766_;
  assign new_n36202_ = ~new_n35762_ & new_n36201_;
  assign new_n36203_ = ~new_n35763_ & ~new_n35766_;
  assign new_n36204_ = ~new_n36202_ & ~new_n36203_;
  assign new_n36205_ = new_n35769_ & ~new_n36204_;
  assign new_n36206_ = ~new_n36200_ & ~new_n36205_;
  assign new_n36207_ = ~\b[32]  & ~new_n36206_;
  assign new_n36208_ = \b[32]  & ~new_n36200_;
  assign new_n36209_ = ~new_n36205_ & new_n36208_;
  assign new_n36210_ = new_n424_ & ~new_n36209_;
  assign new_n36211_ = ~new_n36207_ & new_n36210_;
  assign new_n36212_ = ~new_n36199_ & new_n36211_;
  assign new_n36213_ = new_n432_ & ~new_n36206_;
  assign new_n36214_ = ~new_n36212_ & ~new_n36213_;
  assign new_n36215_ = ~new_n35787_ & new_n36197_;
  assign new_n36216_ = ~new_n36193_ & new_n36215_;
  assign new_n36217_ = ~new_n36194_ & ~new_n36197_;
  assign new_n36218_ = ~new_n36216_ & ~new_n36217_;
  assign new_n36219_ = ~new_n36214_ & ~new_n36218_;
  assign new_n36220_ = ~new_n35777_ & ~new_n36213_;
  assign new_n36221_ = ~new_n36212_ & new_n36220_;
  assign new_n36222_ = ~new_n36219_ & ~new_n36221_;
  assign new_n36223_ = ~new_n35778_ & ~new_n36209_;
  assign new_n36224_ = ~new_n36207_ & new_n36223_;
  assign new_n36225_ = ~new_n36198_ & new_n36224_;
  assign new_n36226_ = ~new_n36207_ & ~new_n36209_;
  assign new_n36227_ = ~new_n36199_ & ~new_n36226_;
  assign new_n36228_ = ~new_n36225_ & ~new_n36227_;
  assign new_n36229_ = ~new_n36214_ & ~new_n36228_;
  assign new_n36230_ = ~new_n36206_ & ~new_n36213_;
  assign new_n36231_ = ~new_n36212_ & new_n36230_;
  assign new_n36232_ = ~new_n36229_ & ~new_n36231_;
  assign new_n36233_ = ~\b[33]  & ~new_n36232_;
  assign new_n36234_ = ~\b[32]  & ~new_n36222_;
  assign new_n36235_ = ~new_n35796_ & new_n36192_;
  assign new_n36236_ = ~new_n36188_ & new_n36235_;
  assign new_n36237_ = ~new_n36189_ & ~new_n36192_;
  assign new_n36238_ = ~new_n36236_ & ~new_n36237_;
  assign new_n36239_ = ~new_n36214_ & ~new_n36238_;
  assign new_n36240_ = ~new_n35786_ & ~new_n36213_;
  assign new_n36241_ = ~new_n36212_ & new_n36240_;
  assign new_n36242_ = ~new_n36239_ & ~new_n36241_;
  assign new_n36243_ = ~\b[31]  & ~new_n36242_;
  assign new_n36244_ = ~new_n35805_ & new_n36187_;
  assign new_n36245_ = ~new_n36183_ & new_n36244_;
  assign new_n36246_ = ~new_n36184_ & ~new_n36187_;
  assign new_n36247_ = ~new_n36245_ & ~new_n36246_;
  assign new_n36248_ = ~new_n36214_ & ~new_n36247_;
  assign new_n36249_ = ~new_n35795_ & ~new_n36213_;
  assign new_n36250_ = ~new_n36212_ & new_n36249_;
  assign new_n36251_ = ~new_n36248_ & ~new_n36250_;
  assign new_n36252_ = ~\b[30]  & ~new_n36251_;
  assign new_n36253_ = ~new_n35814_ & new_n36182_;
  assign new_n36254_ = ~new_n36178_ & new_n36253_;
  assign new_n36255_ = ~new_n36179_ & ~new_n36182_;
  assign new_n36256_ = ~new_n36254_ & ~new_n36255_;
  assign new_n36257_ = ~new_n36214_ & ~new_n36256_;
  assign new_n36258_ = ~new_n35804_ & ~new_n36213_;
  assign new_n36259_ = ~new_n36212_ & new_n36258_;
  assign new_n36260_ = ~new_n36257_ & ~new_n36259_;
  assign new_n36261_ = ~\b[29]  & ~new_n36260_;
  assign new_n36262_ = ~new_n35823_ & new_n36177_;
  assign new_n36263_ = ~new_n36173_ & new_n36262_;
  assign new_n36264_ = ~new_n36174_ & ~new_n36177_;
  assign new_n36265_ = ~new_n36263_ & ~new_n36264_;
  assign new_n36266_ = ~new_n36214_ & ~new_n36265_;
  assign new_n36267_ = ~new_n35813_ & ~new_n36213_;
  assign new_n36268_ = ~new_n36212_ & new_n36267_;
  assign new_n36269_ = ~new_n36266_ & ~new_n36268_;
  assign new_n36270_ = ~\b[28]  & ~new_n36269_;
  assign new_n36271_ = ~new_n35832_ & new_n36172_;
  assign new_n36272_ = ~new_n36168_ & new_n36271_;
  assign new_n36273_ = ~new_n36169_ & ~new_n36172_;
  assign new_n36274_ = ~new_n36272_ & ~new_n36273_;
  assign new_n36275_ = ~new_n36214_ & ~new_n36274_;
  assign new_n36276_ = ~new_n35822_ & ~new_n36213_;
  assign new_n36277_ = ~new_n36212_ & new_n36276_;
  assign new_n36278_ = ~new_n36275_ & ~new_n36277_;
  assign new_n36279_ = ~\b[27]  & ~new_n36278_;
  assign new_n36280_ = ~new_n35841_ & new_n36167_;
  assign new_n36281_ = ~new_n36163_ & new_n36280_;
  assign new_n36282_ = ~new_n36164_ & ~new_n36167_;
  assign new_n36283_ = ~new_n36281_ & ~new_n36282_;
  assign new_n36284_ = ~new_n36214_ & ~new_n36283_;
  assign new_n36285_ = ~new_n35831_ & ~new_n36213_;
  assign new_n36286_ = ~new_n36212_ & new_n36285_;
  assign new_n36287_ = ~new_n36284_ & ~new_n36286_;
  assign new_n36288_ = ~\b[26]  & ~new_n36287_;
  assign new_n36289_ = ~new_n35850_ & new_n36162_;
  assign new_n36290_ = ~new_n36158_ & new_n36289_;
  assign new_n36291_ = ~new_n36159_ & ~new_n36162_;
  assign new_n36292_ = ~new_n36290_ & ~new_n36291_;
  assign new_n36293_ = ~new_n36214_ & ~new_n36292_;
  assign new_n36294_ = ~new_n35840_ & ~new_n36213_;
  assign new_n36295_ = ~new_n36212_ & new_n36294_;
  assign new_n36296_ = ~new_n36293_ & ~new_n36295_;
  assign new_n36297_ = ~\b[25]  & ~new_n36296_;
  assign new_n36298_ = ~new_n35859_ & new_n36157_;
  assign new_n36299_ = ~new_n36153_ & new_n36298_;
  assign new_n36300_ = ~new_n36154_ & ~new_n36157_;
  assign new_n36301_ = ~new_n36299_ & ~new_n36300_;
  assign new_n36302_ = ~new_n36214_ & ~new_n36301_;
  assign new_n36303_ = ~new_n35849_ & ~new_n36213_;
  assign new_n36304_ = ~new_n36212_ & new_n36303_;
  assign new_n36305_ = ~new_n36302_ & ~new_n36304_;
  assign new_n36306_ = ~\b[24]  & ~new_n36305_;
  assign new_n36307_ = ~new_n35868_ & new_n36152_;
  assign new_n36308_ = ~new_n36148_ & new_n36307_;
  assign new_n36309_ = ~new_n36149_ & ~new_n36152_;
  assign new_n36310_ = ~new_n36308_ & ~new_n36309_;
  assign new_n36311_ = ~new_n36214_ & ~new_n36310_;
  assign new_n36312_ = ~new_n35858_ & ~new_n36213_;
  assign new_n36313_ = ~new_n36212_ & new_n36312_;
  assign new_n36314_ = ~new_n36311_ & ~new_n36313_;
  assign new_n36315_ = ~\b[23]  & ~new_n36314_;
  assign new_n36316_ = ~new_n35877_ & new_n36147_;
  assign new_n36317_ = ~new_n36143_ & new_n36316_;
  assign new_n36318_ = ~new_n36144_ & ~new_n36147_;
  assign new_n36319_ = ~new_n36317_ & ~new_n36318_;
  assign new_n36320_ = ~new_n36214_ & ~new_n36319_;
  assign new_n36321_ = ~new_n35867_ & ~new_n36213_;
  assign new_n36322_ = ~new_n36212_ & new_n36321_;
  assign new_n36323_ = ~new_n36320_ & ~new_n36322_;
  assign new_n36324_ = ~\b[22]  & ~new_n36323_;
  assign new_n36325_ = ~new_n35886_ & new_n36142_;
  assign new_n36326_ = ~new_n36138_ & new_n36325_;
  assign new_n36327_ = ~new_n36139_ & ~new_n36142_;
  assign new_n36328_ = ~new_n36326_ & ~new_n36327_;
  assign new_n36329_ = ~new_n36214_ & ~new_n36328_;
  assign new_n36330_ = ~new_n35876_ & ~new_n36213_;
  assign new_n36331_ = ~new_n36212_ & new_n36330_;
  assign new_n36332_ = ~new_n36329_ & ~new_n36331_;
  assign new_n36333_ = ~\b[21]  & ~new_n36332_;
  assign new_n36334_ = ~new_n35895_ & new_n36137_;
  assign new_n36335_ = ~new_n36133_ & new_n36334_;
  assign new_n36336_ = ~new_n36134_ & ~new_n36137_;
  assign new_n36337_ = ~new_n36335_ & ~new_n36336_;
  assign new_n36338_ = ~new_n36214_ & ~new_n36337_;
  assign new_n36339_ = ~new_n35885_ & ~new_n36213_;
  assign new_n36340_ = ~new_n36212_ & new_n36339_;
  assign new_n36341_ = ~new_n36338_ & ~new_n36340_;
  assign new_n36342_ = ~\b[20]  & ~new_n36341_;
  assign new_n36343_ = ~new_n35904_ & new_n36132_;
  assign new_n36344_ = ~new_n36128_ & new_n36343_;
  assign new_n36345_ = ~new_n36129_ & ~new_n36132_;
  assign new_n36346_ = ~new_n36344_ & ~new_n36345_;
  assign new_n36347_ = ~new_n36214_ & ~new_n36346_;
  assign new_n36348_ = ~new_n35894_ & ~new_n36213_;
  assign new_n36349_ = ~new_n36212_ & new_n36348_;
  assign new_n36350_ = ~new_n36347_ & ~new_n36349_;
  assign new_n36351_ = ~\b[19]  & ~new_n36350_;
  assign new_n36352_ = ~new_n35913_ & new_n36127_;
  assign new_n36353_ = ~new_n36123_ & new_n36352_;
  assign new_n36354_ = ~new_n36124_ & ~new_n36127_;
  assign new_n36355_ = ~new_n36353_ & ~new_n36354_;
  assign new_n36356_ = ~new_n36214_ & ~new_n36355_;
  assign new_n36357_ = ~new_n35903_ & ~new_n36213_;
  assign new_n36358_ = ~new_n36212_ & new_n36357_;
  assign new_n36359_ = ~new_n36356_ & ~new_n36358_;
  assign new_n36360_ = ~\b[18]  & ~new_n36359_;
  assign new_n36361_ = ~new_n35922_ & new_n36122_;
  assign new_n36362_ = ~new_n36118_ & new_n36361_;
  assign new_n36363_ = ~new_n36119_ & ~new_n36122_;
  assign new_n36364_ = ~new_n36362_ & ~new_n36363_;
  assign new_n36365_ = ~new_n36214_ & ~new_n36364_;
  assign new_n36366_ = ~new_n35912_ & ~new_n36213_;
  assign new_n36367_ = ~new_n36212_ & new_n36366_;
  assign new_n36368_ = ~new_n36365_ & ~new_n36367_;
  assign new_n36369_ = ~\b[17]  & ~new_n36368_;
  assign new_n36370_ = ~new_n35931_ & new_n36117_;
  assign new_n36371_ = ~new_n36113_ & new_n36370_;
  assign new_n36372_ = ~new_n36114_ & ~new_n36117_;
  assign new_n36373_ = ~new_n36371_ & ~new_n36372_;
  assign new_n36374_ = ~new_n36214_ & ~new_n36373_;
  assign new_n36375_ = ~new_n35921_ & ~new_n36213_;
  assign new_n36376_ = ~new_n36212_ & new_n36375_;
  assign new_n36377_ = ~new_n36374_ & ~new_n36376_;
  assign new_n36378_ = ~\b[16]  & ~new_n36377_;
  assign new_n36379_ = ~new_n35940_ & new_n36112_;
  assign new_n36380_ = ~new_n36108_ & new_n36379_;
  assign new_n36381_ = ~new_n36109_ & ~new_n36112_;
  assign new_n36382_ = ~new_n36380_ & ~new_n36381_;
  assign new_n36383_ = ~new_n36214_ & ~new_n36382_;
  assign new_n36384_ = ~new_n35930_ & ~new_n36213_;
  assign new_n36385_ = ~new_n36212_ & new_n36384_;
  assign new_n36386_ = ~new_n36383_ & ~new_n36385_;
  assign new_n36387_ = ~\b[15]  & ~new_n36386_;
  assign new_n36388_ = ~new_n35949_ & new_n36107_;
  assign new_n36389_ = ~new_n36103_ & new_n36388_;
  assign new_n36390_ = ~new_n36104_ & ~new_n36107_;
  assign new_n36391_ = ~new_n36389_ & ~new_n36390_;
  assign new_n36392_ = ~new_n36214_ & ~new_n36391_;
  assign new_n36393_ = ~new_n35939_ & ~new_n36213_;
  assign new_n36394_ = ~new_n36212_ & new_n36393_;
  assign new_n36395_ = ~new_n36392_ & ~new_n36394_;
  assign new_n36396_ = ~\b[14]  & ~new_n36395_;
  assign new_n36397_ = ~new_n35958_ & new_n36102_;
  assign new_n36398_ = ~new_n36098_ & new_n36397_;
  assign new_n36399_ = ~new_n36099_ & ~new_n36102_;
  assign new_n36400_ = ~new_n36398_ & ~new_n36399_;
  assign new_n36401_ = ~new_n36214_ & ~new_n36400_;
  assign new_n36402_ = ~new_n35948_ & ~new_n36213_;
  assign new_n36403_ = ~new_n36212_ & new_n36402_;
  assign new_n36404_ = ~new_n36401_ & ~new_n36403_;
  assign new_n36405_ = ~\b[13]  & ~new_n36404_;
  assign new_n36406_ = ~new_n35967_ & new_n36097_;
  assign new_n36407_ = ~new_n36093_ & new_n36406_;
  assign new_n36408_ = ~new_n36094_ & ~new_n36097_;
  assign new_n36409_ = ~new_n36407_ & ~new_n36408_;
  assign new_n36410_ = ~new_n36214_ & ~new_n36409_;
  assign new_n36411_ = ~new_n35957_ & ~new_n36213_;
  assign new_n36412_ = ~new_n36212_ & new_n36411_;
  assign new_n36413_ = ~new_n36410_ & ~new_n36412_;
  assign new_n36414_ = ~\b[12]  & ~new_n36413_;
  assign new_n36415_ = ~new_n35976_ & new_n36092_;
  assign new_n36416_ = ~new_n36088_ & new_n36415_;
  assign new_n36417_ = ~new_n36089_ & ~new_n36092_;
  assign new_n36418_ = ~new_n36416_ & ~new_n36417_;
  assign new_n36419_ = ~new_n36214_ & ~new_n36418_;
  assign new_n36420_ = ~new_n35966_ & ~new_n36213_;
  assign new_n36421_ = ~new_n36212_ & new_n36420_;
  assign new_n36422_ = ~new_n36419_ & ~new_n36421_;
  assign new_n36423_ = ~\b[11]  & ~new_n36422_;
  assign new_n36424_ = ~new_n35985_ & new_n36087_;
  assign new_n36425_ = ~new_n36083_ & new_n36424_;
  assign new_n36426_ = ~new_n36084_ & ~new_n36087_;
  assign new_n36427_ = ~new_n36425_ & ~new_n36426_;
  assign new_n36428_ = ~new_n36214_ & ~new_n36427_;
  assign new_n36429_ = ~new_n35975_ & ~new_n36213_;
  assign new_n36430_ = ~new_n36212_ & new_n36429_;
  assign new_n36431_ = ~new_n36428_ & ~new_n36430_;
  assign new_n36432_ = ~\b[10]  & ~new_n36431_;
  assign new_n36433_ = ~new_n35994_ & new_n36082_;
  assign new_n36434_ = ~new_n36078_ & new_n36433_;
  assign new_n36435_ = ~new_n36079_ & ~new_n36082_;
  assign new_n36436_ = ~new_n36434_ & ~new_n36435_;
  assign new_n36437_ = ~new_n36214_ & ~new_n36436_;
  assign new_n36438_ = ~new_n35984_ & ~new_n36213_;
  assign new_n36439_ = ~new_n36212_ & new_n36438_;
  assign new_n36440_ = ~new_n36437_ & ~new_n36439_;
  assign new_n36441_ = ~\b[9]  & ~new_n36440_;
  assign new_n36442_ = ~new_n36003_ & new_n36077_;
  assign new_n36443_ = ~new_n36073_ & new_n36442_;
  assign new_n36444_ = ~new_n36074_ & ~new_n36077_;
  assign new_n36445_ = ~new_n36443_ & ~new_n36444_;
  assign new_n36446_ = ~new_n36214_ & ~new_n36445_;
  assign new_n36447_ = ~new_n35993_ & ~new_n36213_;
  assign new_n36448_ = ~new_n36212_ & new_n36447_;
  assign new_n36449_ = ~new_n36446_ & ~new_n36448_;
  assign new_n36450_ = ~\b[8]  & ~new_n36449_;
  assign new_n36451_ = ~new_n36012_ & new_n36072_;
  assign new_n36452_ = ~new_n36068_ & new_n36451_;
  assign new_n36453_ = ~new_n36069_ & ~new_n36072_;
  assign new_n36454_ = ~new_n36452_ & ~new_n36453_;
  assign new_n36455_ = ~new_n36214_ & ~new_n36454_;
  assign new_n36456_ = ~new_n36002_ & ~new_n36213_;
  assign new_n36457_ = ~new_n36212_ & new_n36456_;
  assign new_n36458_ = ~new_n36455_ & ~new_n36457_;
  assign new_n36459_ = ~\b[7]  & ~new_n36458_;
  assign new_n36460_ = ~new_n36021_ & new_n36067_;
  assign new_n36461_ = ~new_n36063_ & new_n36460_;
  assign new_n36462_ = ~new_n36064_ & ~new_n36067_;
  assign new_n36463_ = ~new_n36461_ & ~new_n36462_;
  assign new_n36464_ = ~new_n36214_ & ~new_n36463_;
  assign new_n36465_ = ~new_n36011_ & ~new_n36213_;
  assign new_n36466_ = ~new_n36212_ & new_n36465_;
  assign new_n36467_ = ~new_n36464_ & ~new_n36466_;
  assign new_n36468_ = ~\b[6]  & ~new_n36467_;
  assign new_n36469_ = ~new_n36030_ & new_n36062_;
  assign new_n36470_ = ~new_n36058_ & new_n36469_;
  assign new_n36471_ = ~new_n36059_ & ~new_n36062_;
  assign new_n36472_ = ~new_n36470_ & ~new_n36471_;
  assign new_n36473_ = ~new_n36214_ & ~new_n36472_;
  assign new_n36474_ = ~new_n36020_ & ~new_n36213_;
  assign new_n36475_ = ~new_n36212_ & new_n36474_;
  assign new_n36476_ = ~new_n36473_ & ~new_n36475_;
  assign new_n36477_ = ~\b[5]  & ~new_n36476_;
  assign new_n36478_ = ~new_n36038_ & new_n36057_;
  assign new_n36479_ = ~new_n36053_ & new_n36478_;
  assign new_n36480_ = ~new_n36054_ & ~new_n36057_;
  assign new_n36481_ = ~new_n36479_ & ~new_n36480_;
  assign new_n36482_ = ~new_n36214_ & ~new_n36481_;
  assign new_n36483_ = ~new_n36029_ & ~new_n36213_;
  assign new_n36484_ = ~new_n36212_ & new_n36483_;
  assign new_n36485_ = ~new_n36482_ & ~new_n36484_;
  assign new_n36486_ = ~\b[4]  & ~new_n36485_;
  assign new_n36487_ = ~new_n36048_ & new_n36052_;
  assign new_n36488_ = ~new_n36047_ & new_n36487_;
  assign new_n36489_ = ~new_n36049_ & ~new_n36052_;
  assign new_n36490_ = ~new_n36488_ & ~new_n36489_;
  assign new_n36491_ = ~new_n36214_ & ~new_n36490_;
  assign new_n36492_ = ~new_n36037_ & ~new_n36213_;
  assign new_n36493_ = ~new_n36212_ & new_n36492_;
  assign new_n36494_ = ~new_n36491_ & ~new_n36493_;
  assign new_n36495_ = ~\b[3]  & ~new_n36494_;
  assign new_n36496_ = new_n7887_ & ~new_n36045_;
  assign new_n36497_ = ~new_n36043_ & new_n36496_;
  assign new_n36498_ = ~new_n36047_ & ~new_n36497_;
  assign new_n36499_ = ~new_n36214_ & new_n36498_;
  assign new_n36500_ = ~new_n36042_ & ~new_n36213_;
  assign new_n36501_ = ~new_n36212_ & new_n36500_;
  assign new_n36502_ = ~new_n36499_ & ~new_n36501_;
  assign new_n36503_ = ~\b[2]  & ~new_n36502_;
  assign new_n36504_ = \b[0]  & ~new_n36214_;
  assign new_n36505_ = \a[31]  & ~new_n36504_;
  assign new_n36506_ = new_n7887_ & ~new_n36214_;
  assign new_n36507_ = ~new_n36505_ & ~new_n36506_;
  assign new_n36508_ = \b[1]  & ~new_n36507_;
  assign new_n36509_ = ~\b[1]  & ~new_n36506_;
  assign new_n36510_ = ~new_n36505_ & new_n36509_;
  assign new_n36511_ = ~new_n36508_ & ~new_n36510_;
  assign new_n36512_ = ~new_n8353_ & ~new_n36511_;
  assign new_n36513_ = ~\b[1]  & ~new_n36507_;
  assign new_n36514_ = ~new_n36512_ & ~new_n36513_;
  assign new_n36515_ = \b[2]  & ~new_n36501_;
  assign new_n36516_ = ~new_n36499_ & new_n36515_;
  assign new_n36517_ = ~new_n36503_ & ~new_n36516_;
  assign new_n36518_ = ~new_n36514_ & new_n36517_;
  assign new_n36519_ = ~new_n36503_ & ~new_n36518_;
  assign new_n36520_ = \b[3]  & ~new_n36493_;
  assign new_n36521_ = ~new_n36491_ & new_n36520_;
  assign new_n36522_ = ~new_n36495_ & ~new_n36521_;
  assign new_n36523_ = ~new_n36519_ & new_n36522_;
  assign new_n36524_ = ~new_n36495_ & ~new_n36523_;
  assign new_n36525_ = \b[4]  & ~new_n36484_;
  assign new_n36526_ = ~new_n36482_ & new_n36525_;
  assign new_n36527_ = ~new_n36486_ & ~new_n36526_;
  assign new_n36528_ = ~new_n36524_ & new_n36527_;
  assign new_n36529_ = ~new_n36486_ & ~new_n36528_;
  assign new_n36530_ = \b[5]  & ~new_n36475_;
  assign new_n36531_ = ~new_n36473_ & new_n36530_;
  assign new_n36532_ = ~new_n36477_ & ~new_n36531_;
  assign new_n36533_ = ~new_n36529_ & new_n36532_;
  assign new_n36534_ = ~new_n36477_ & ~new_n36533_;
  assign new_n36535_ = \b[6]  & ~new_n36466_;
  assign new_n36536_ = ~new_n36464_ & new_n36535_;
  assign new_n36537_ = ~new_n36468_ & ~new_n36536_;
  assign new_n36538_ = ~new_n36534_ & new_n36537_;
  assign new_n36539_ = ~new_n36468_ & ~new_n36538_;
  assign new_n36540_ = \b[7]  & ~new_n36457_;
  assign new_n36541_ = ~new_n36455_ & new_n36540_;
  assign new_n36542_ = ~new_n36459_ & ~new_n36541_;
  assign new_n36543_ = ~new_n36539_ & new_n36542_;
  assign new_n36544_ = ~new_n36459_ & ~new_n36543_;
  assign new_n36545_ = \b[8]  & ~new_n36448_;
  assign new_n36546_ = ~new_n36446_ & new_n36545_;
  assign new_n36547_ = ~new_n36450_ & ~new_n36546_;
  assign new_n36548_ = ~new_n36544_ & new_n36547_;
  assign new_n36549_ = ~new_n36450_ & ~new_n36548_;
  assign new_n36550_ = \b[9]  & ~new_n36439_;
  assign new_n36551_ = ~new_n36437_ & new_n36550_;
  assign new_n36552_ = ~new_n36441_ & ~new_n36551_;
  assign new_n36553_ = ~new_n36549_ & new_n36552_;
  assign new_n36554_ = ~new_n36441_ & ~new_n36553_;
  assign new_n36555_ = \b[10]  & ~new_n36430_;
  assign new_n36556_ = ~new_n36428_ & new_n36555_;
  assign new_n36557_ = ~new_n36432_ & ~new_n36556_;
  assign new_n36558_ = ~new_n36554_ & new_n36557_;
  assign new_n36559_ = ~new_n36432_ & ~new_n36558_;
  assign new_n36560_ = \b[11]  & ~new_n36421_;
  assign new_n36561_ = ~new_n36419_ & new_n36560_;
  assign new_n36562_ = ~new_n36423_ & ~new_n36561_;
  assign new_n36563_ = ~new_n36559_ & new_n36562_;
  assign new_n36564_ = ~new_n36423_ & ~new_n36563_;
  assign new_n36565_ = \b[12]  & ~new_n36412_;
  assign new_n36566_ = ~new_n36410_ & new_n36565_;
  assign new_n36567_ = ~new_n36414_ & ~new_n36566_;
  assign new_n36568_ = ~new_n36564_ & new_n36567_;
  assign new_n36569_ = ~new_n36414_ & ~new_n36568_;
  assign new_n36570_ = \b[13]  & ~new_n36403_;
  assign new_n36571_ = ~new_n36401_ & new_n36570_;
  assign new_n36572_ = ~new_n36405_ & ~new_n36571_;
  assign new_n36573_ = ~new_n36569_ & new_n36572_;
  assign new_n36574_ = ~new_n36405_ & ~new_n36573_;
  assign new_n36575_ = \b[14]  & ~new_n36394_;
  assign new_n36576_ = ~new_n36392_ & new_n36575_;
  assign new_n36577_ = ~new_n36396_ & ~new_n36576_;
  assign new_n36578_ = ~new_n36574_ & new_n36577_;
  assign new_n36579_ = ~new_n36396_ & ~new_n36578_;
  assign new_n36580_ = \b[15]  & ~new_n36385_;
  assign new_n36581_ = ~new_n36383_ & new_n36580_;
  assign new_n36582_ = ~new_n36387_ & ~new_n36581_;
  assign new_n36583_ = ~new_n36579_ & new_n36582_;
  assign new_n36584_ = ~new_n36387_ & ~new_n36583_;
  assign new_n36585_ = \b[16]  & ~new_n36376_;
  assign new_n36586_ = ~new_n36374_ & new_n36585_;
  assign new_n36587_ = ~new_n36378_ & ~new_n36586_;
  assign new_n36588_ = ~new_n36584_ & new_n36587_;
  assign new_n36589_ = ~new_n36378_ & ~new_n36588_;
  assign new_n36590_ = \b[17]  & ~new_n36367_;
  assign new_n36591_ = ~new_n36365_ & new_n36590_;
  assign new_n36592_ = ~new_n36369_ & ~new_n36591_;
  assign new_n36593_ = ~new_n36589_ & new_n36592_;
  assign new_n36594_ = ~new_n36369_ & ~new_n36593_;
  assign new_n36595_ = \b[18]  & ~new_n36358_;
  assign new_n36596_ = ~new_n36356_ & new_n36595_;
  assign new_n36597_ = ~new_n36360_ & ~new_n36596_;
  assign new_n36598_ = ~new_n36594_ & new_n36597_;
  assign new_n36599_ = ~new_n36360_ & ~new_n36598_;
  assign new_n36600_ = \b[19]  & ~new_n36349_;
  assign new_n36601_ = ~new_n36347_ & new_n36600_;
  assign new_n36602_ = ~new_n36351_ & ~new_n36601_;
  assign new_n36603_ = ~new_n36599_ & new_n36602_;
  assign new_n36604_ = ~new_n36351_ & ~new_n36603_;
  assign new_n36605_ = \b[20]  & ~new_n36340_;
  assign new_n36606_ = ~new_n36338_ & new_n36605_;
  assign new_n36607_ = ~new_n36342_ & ~new_n36606_;
  assign new_n36608_ = ~new_n36604_ & new_n36607_;
  assign new_n36609_ = ~new_n36342_ & ~new_n36608_;
  assign new_n36610_ = \b[21]  & ~new_n36331_;
  assign new_n36611_ = ~new_n36329_ & new_n36610_;
  assign new_n36612_ = ~new_n36333_ & ~new_n36611_;
  assign new_n36613_ = ~new_n36609_ & new_n36612_;
  assign new_n36614_ = ~new_n36333_ & ~new_n36613_;
  assign new_n36615_ = \b[22]  & ~new_n36322_;
  assign new_n36616_ = ~new_n36320_ & new_n36615_;
  assign new_n36617_ = ~new_n36324_ & ~new_n36616_;
  assign new_n36618_ = ~new_n36614_ & new_n36617_;
  assign new_n36619_ = ~new_n36324_ & ~new_n36618_;
  assign new_n36620_ = \b[23]  & ~new_n36313_;
  assign new_n36621_ = ~new_n36311_ & new_n36620_;
  assign new_n36622_ = ~new_n36315_ & ~new_n36621_;
  assign new_n36623_ = ~new_n36619_ & new_n36622_;
  assign new_n36624_ = ~new_n36315_ & ~new_n36623_;
  assign new_n36625_ = \b[24]  & ~new_n36304_;
  assign new_n36626_ = ~new_n36302_ & new_n36625_;
  assign new_n36627_ = ~new_n36306_ & ~new_n36626_;
  assign new_n36628_ = ~new_n36624_ & new_n36627_;
  assign new_n36629_ = ~new_n36306_ & ~new_n36628_;
  assign new_n36630_ = \b[25]  & ~new_n36295_;
  assign new_n36631_ = ~new_n36293_ & new_n36630_;
  assign new_n36632_ = ~new_n36297_ & ~new_n36631_;
  assign new_n36633_ = ~new_n36629_ & new_n36632_;
  assign new_n36634_ = ~new_n36297_ & ~new_n36633_;
  assign new_n36635_ = \b[26]  & ~new_n36286_;
  assign new_n36636_ = ~new_n36284_ & new_n36635_;
  assign new_n36637_ = ~new_n36288_ & ~new_n36636_;
  assign new_n36638_ = ~new_n36634_ & new_n36637_;
  assign new_n36639_ = ~new_n36288_ & ~new_n36638_;
  assign new_n36640_ = \b[27]  & ~new_n36277_;
  assign new_n36641_ = ~new_n36275_ & new_n36640_;
  assign new_n36642_ = ~new_n36279_ & ~new_n36641_;
  assign new_n36643_ = ~new_n36639_ & new_n36642_;
  assign new_n36644_ = ~new_n36279_ & ~new_n36643_;
  assign new_n36645_ = \b[28]  & ~new_n36268_;
  assign new_n36646_ = ~new_n36266_ & new_n36645_;
  assign new_n36647_ = ~new_n36270_ & ~new_n36646_;
  assign new_n36648_ = ~new_n36644_ & new_n36647_;
  assign new_n36649_ = ~new_n36270_ & ~new_n36648_;
  assign new_n36650_ = \b[29]  & ~new_n36259_;
  assign new_n36651_ = ~new_n36257_ & new_n36650_;
  assign new_n36652_ = ~new_n36261_ & ~new_n36651_;
  assign new_n36653_ = ~new_n36649_ & new_n36652_;
  assign new_n36654_ = ~new_n36261_ & ~new_n36653_;
  assign new_n36655_ = \b[30]  & ~new_n36250_;
  assign new_n36656_ = ~new_n36248_ & new_n36655_;
  assign new_n36657_ = ~new_n36252_ & ~new_n36656_;
  assign new_n36658_ = ~new_n36654_ & new_n36657_;
  assign new_n36659_ = ~new_n36252_ & ~new_n36658_;
  assign new_n36660_ = \b[31]  & ~new_n36241_;
  assign new_n36661_ = ~new_n36239_ & new_n36660_;
  assign new_n36662_ = ~new_n36243_ & ~new_n36661_;
  assign new_n36663_ = ~new_n36659_ & new_n36662_;
  assign new_n36664_ = ~new_n36243_ & ~new_n36663_;
  assign new_n36665_ = \b[32]  & ~new_n36221_;
  assign new_n36666_ = ~new_n36219_ & new_n36665_;
  assign new_n36667_ = ~new_n36234_ & ~new_n36666_;
  assign new_n36668_ = ~new_n36664_ & new_n36667_;
  assign new_n36669_ = ~new_n36234_ & ~new_n36668_;
  assign new_n36670_ = \b[33]  & ~new_n36231_;
  assign new_n36671_ = ~new_n36229_ & new_n36670_;
  assign new_n36672_ = ~new_n36233_ & ~new_n36671_;
  assign new_n36673_ = ~new_n36669_ & new_n36672_;
  assign new_n36674_ = ~new_n36233_ & ~new_n36673_;
  assign new_n36675_ = new_n8519_ & ~new_n36674_;
  assign new_n36676_ = ~new_n36222_ & ~new_n36675_;
  assign new_n36677_ = ~new_n36243_ & new_n36667_;
  assign new_n36678_ = ~new_n36663_ & new_n36677_;
  assign new_n36679_ = ~new_n36664_ & ~new_n36667_;
  assign new_n36680_ = ~new_n36678_ & ~new_n36679_;
  assign new_n36681_ = new_n8519_ & ~new_n36680_;
  assign new_n36682_ = ~new_n36674_ & new_n36681_;
  assign new_n36683_ = ~new_n36676_ & ~new_n36682_;
  assign new_n36684_ = ~new_n36232_ & ~new_n36675_;
  assign new_n36685_ = ~new_n36234_ & new_n36672_;
  assign new_n36686_ = ~new_n36668_ & new_n36685_;
  assign new_n36687_ = ~new_n36669_ & ~new_n36672_;
  assign new_n36688_ = ~new_n36686_ & ~new_n36687_;
  assign new_n36689_ = new_n36675_ & ~new_n36688_;
  assign new_n36690_ = ~new_n36684_ & ~new_n36689_;
  assign new_n36691_ = ~\b[34]  & ~new_n36690_;
  assign new_n36692_ = ~\b[33]  & ~new_n36683_;
  assign new_n36693_ = ~new_n36242_ & ~new_n36675_;
  assign new_n36694_ = ~new_n36252_ & new_n36662_;
  assign new_n36695_ = ~new_n36658_ & new_n36694_;
  assign new_n36696_ = ~new_n36659_ & ~new_n36662_;
  assign new_n36697_ = ~new_n36695_ & ~new_n36696_;
  assign new_n36698_ = new_n8519_ & ~new_n36697_;
  assign new_n36699_ = ~new_n36674_ & new_n36698_;
  assign new_n36700_ = ~new_n36693_ & ~new_n36699_;
  assign new_n36701_ = ~\b[32]  & ~new_n36700_;
  assign new_n36702_ = ~new_n36251_ & ~new_n36675_;
  assign new_n36703_ = ~new_n36261_ & new_n36657_;
  assign new_n36704_ = ~new_n36653_ & new_n36703_;
  assign new_n36705_ = ~new_n36654_ & ~new_n36657_;
  assign new_n36706_ = ~new_n36704_ & ~new_n36705_;
  assign new_n36707_ = new_n8519_ & ~new_n36706_;
  assign new_n36708_ = ~new_n36674_ & new_n36707_;
  assign new_n36709_ = ~new_n36702_ & ~new_n36708_;
  assign new_n36710_ = ~\b[31]  & ~new_n36709_;
  assign new_n36711_ = ~new_n36260_ & ~new_n36675_;
  assign new_n36712_ = ~new_n36270_ & new_n36652_;
  assign new_n36713_ = ~new_n36648_ & new_n36712_;
  assign new_n36714_ = ~new_n36649_ & ~new_n36652_;
  assign new_n36715_ = ~new_n36713_ & ~new_n36714_;
  assign new_n36716_ = new_n8519_ & ~new_n36715_;
  assign new_n36717_ = ~new_n36674_ & new_n36716_;
  assign new_n36718_ = ~new_n36711_ & ~new_n36717_;
  assign new_n36719_ = ~\b[30]  & ~new_n36718_;
  assign new_n36720_ = ~new_n36269_ & ~new_n36675_;
  assign new_n36721_ = ~new_n36279_ & new_n36647_;
  assign new_n36722_ = ~new_n36643_ & new_n36721_;
  assign new_n36723_ = ~new_n36644_ & ~new_n36647_;
  assign new_n36724_ = ~new_n36722_ & ~new_n36723_;
  assign new_n36725_ = new_n8519_ & ~new_n36724_;
  assign new_n36726_ = ~new_n36674_ & new_n36725_;
  assign new_n36727_ = ~new_n36720_ & ~new_n36726_;
  assign new_n36728_ = ~\b[29]  & ~new_n36727_;
  assign new_n36729_ = ~new_n36278_ & ~new_n36675_;
  assign new_n36730_ = ~new_n36288_ & new_n36642_;
  assign new_n36731_ = ~new_n36638_ & new_n36730_;
  assign new_n36732_ = ~new_n36639_ & ~new_n36642_;
  assign new_n36733_ = ~new_n36731_ & ~new_n36732_;
  assign new_n36734_ = new_n8519_ & ~new_n36733_;
  assign new_n36735_ = ~new_n36674_ & new_n36734_;
  assign new_n36736_ = ~new_n36729_ & ~new_n36735_;
  assign new_n36737_ = ~\b[28]  & ~new_n36736_;
  assign new_n36738_ = ~new_n36287_ & ~new_n36675_;
  assign new_n36739_ = ~new_n36297_ & new_n36637_;
  assign new_n36740_ = ~new_n36633_ & new_n36739_;
  assign new_n36741_ = ~new_n36634_ & ~new_n36637_;
  assign new_n36742_ = ~new_n36740_ & ~new_n36741_;
  assign new_n36743_ = new_n8519_ & ~new_n36742_;
  assign new_n36744_ = ~new_n36674_ & new_n36743_;
  assign new_n36745_ = ~new_n36738_ & ~new_n36744_;
  assign new_n36746_ = ~\b[27]  & ~new_n36745_;
  assign new_n36747_ = ~new_n36296_ & ~new_n36675_;
  assign new_n36748_ = ~new_n36306_ & new_n36632_;
  assign new_n36749_ = ~new_n36628_ & new_n36748_;
  assign new_n36750_ = ~new_n36629_ & ~new_n36632_;
  assign new_n36751_ = ~new_n36749_ & ~new_n36750_;
  assign new_n36752_ = new_n8519_ & ~new_n36751_;
  assign new_n36753_ = ~new_n36674_ & new_n36752_;
  assign new_n36754_ = ~new_n36747_ & ~new_n36753_;
  assign new_n36755_ = ~\b[26]  & ~new_n36754_;
  assign new_n36756_ = ~new_n36305_ & ~new_n36675_;
  assign new_n36757_ = ~new_n36315_ & new_n36627_;
  assign new_n36758_ = ~new_n36623_ & new_n36757_;
  assign new_n36759_ = ~new_n36624_ & ~new_n36627_;
  assign new_n36760_ = ~new_n36758_ & ~new_n36759_;
  assign new_n36761_ = new_n8519_ & ~new_n36760_;
  assign new_n36762_ = ~new_n36674_ & new_n36761_;
  assign new_n36763_ = ~new_n36756_ & ~new_n36762_;
  assign new_n36764_ = ~\b[25]  & ~new_n36763_;
  assign new_n36765_ = ~new_n36314_ & ~new_n36675_;
  assign new_n36766_ = ~new_n36324_ & new_n36622_;
  assign new_n36767_ = ~new_n36618_ & new_n36766_;
  assign new_n36768_ = ~new_n36619_ & ~new_n36622_;
  assign new_n36769_ = ~new_n36767_ & ~new_n36768_;
  assign new_n36770_ = new_n8519_ & ~new_n36769_;
  assign new_n36771_ = ~new_n36674_ & new_n36770_;
  assign new_n36772_ = ~new_n36765_ & ~new_n36771_;
  assign new_n36773_ = ~\b[24]  & ~new_n36772_;
  assign new_n36774_ = ~new_n36323_ & ~new_n36675_;
  assign new_n36775_ = ~new_n36333_ & new_n36617_;
  assign new_n36776_ = ~new_n36613_ & new_n36775_;
  assign new_n36777_ = ~new_n36614_ & ~new_n36617_;
  assign new_n36778_ = ~new_n36776_ & ~new_n36777_;
  assign new_n36779_ = new_n8519_ & ~new_n36778_;
  assign new_n36780_ = ~new_n36674_ & new_n36779_;
  assign new_n36781_ = ~new_n36774_ & ~new_n36780_;
  assign new_n36782_ = ~\b[23]  & ~new_n36781_;
  assign new_n36783_ = ~new_n36332_ & ~new_n36675_;
  assign new_n36784_ = ~new_n36342_ & new_n36612_;
  assign new_n36785_ = ~new_n36608_ & new_n36784_;
  assign new_n36786_ = ~new_n36609_ & ~new_n36612_;
  assign new_n36787_ = ~new_n36785_ & ~new_n36786_;
  assign new_n36788_ = new_n8519_ & ~new_n36787_;
  assign new_n36789_ = ~new_n36674_ & new_n36788_;
  assign new_n36790_ = ~new_n36783_ & ~new_n36789_;
  assign new_n36791_ = ~\b[22]  & ~new_n36790_;
  assign new_n36792_ = ~new_n36341_ & ~new_n36675_;
  assign new_n36793_ = ~new_n36351_ & new_n36607_;
  assign new_n36794_ = ~new_n36603_ & new_n36793_;
  assign new_n36795_ = ~new_n36604_ & ~new_n36607_;
  assign new_n36796_ = ~new_n36794_ & ~new_n36795_;
  assign new_n36797_ = new_n8519_ & ~new_n36796_;
  assign new_n36798_ = ~new_n36674_ & new_n36797_;
  assign new_n36799_ = ~new_n36792_ & ~new_n36798_;
  assign new_n36800_ = ~\b[21]  & ~new_n36799_;
  assign new_n36801_ = ~new_n36350_ & ~new_n36675_;
  assign new_n36802_ = ~new_n36360_ & new_n36602_;
  assign new_n36803_ = ~new_n36598_ & new_n36802_;
  assign new_n36804_ = ~new_n36599_ & ~new_n36602_;
  assign new_n36805_ = ~new_n36803_ & ~new_n36804_;
  assign new_n36806_ = new_n8519_ & ~new_n36805_;
  assign new_n36807_ = ~new_n36674_ & new_n36806_;
  assign new_n36808_ = ~new_n36801_ & ~new_n36807_;
  assign new_n36809_ = ~\b[20]  & ~new_n36808_;
  assign new_n36810_ = ~new_n36359_ & ~new_n36675_;
  assign new_n36811_ = ~new_n36369_ & new_n36597_;
  assign new_n36812_ = ~new_n36593_ & new_n36811_;
  assign new_n36813_ = ~new_n36594_ & ~new_n36597_;
  assign new_n36814_ = ~new_n36812_ & ~new_n36813_;
  assign new_n36815_ = new_n8519_ & ~new_n36814_;
  assign new_n36816_ = ~new_n36674_ & new_n36815_;
  assign new_n36817_ = ~new_n36810_ & ~new_n36816_;
  assign new_n36818_ = ~\b[19]  & ~new_n36817_;
  assign new_n36819_ = ~new_n36368_ & ~new_n36675_;
  assign new_n36820_ = ~new_n36378_ & new_n36592_;
  assign new_n36821_ = ~new_n36588_ & new_n36820_;
  assign new_n36822_ = ~new_n36589_ & ~new_n36592_;
  assign new_n36823_ = ~new_n36821_ & ~new_n36822_;
  assign new_n36824_ = new_n8519_ & ~new_n36823_;
  assign new_n36825_ = ~new_n36674_ & new_n36824_;
  assign new_n36826_ = ~new_n36819_ & ~new_n36825_;
  assign new_n36827_ = ~\b[18]  & ~new_n36826_;
  assign new_n36828_ = ~new_n36377_ & ~new_n36675_;
  assign new_n36829_ = ~new_n36387_ & new_n36587_;
  assign new_n36830_ = ~new_n36583_ & new_n36829_;
  assign new_n36831_ = ~new_n36584_ & ~new_n36587_;
  assign new_n36832_ = ~new_n36830_ & ~new_n36831_;
  assign new_n36833_ = new_n8519_ & ~new_n36832_;
  assign new_n36834_ = ~new_n36674_ & new_n36833_;
  assign new_n36835_ = ~new_n36828_ & ~new_n36834_;
  assign new_n36836_ = ~\b[17]  & ~new_n36835_;
  assign new_n36837_ = ~new_n36386_ & ~new_n36675_;
  assign new_n36838_ = ~new_n36396_ & new_n36582_;
  assign new_n36839_ = ~new_n36578_ & new_n36838_;
  assign new_n36840_ = ~new_n36579_ & ~new_n36582_;
  assign new_n36841_ = ~new_n36839_ & ~new_n36840_;
  assign new_n36842_ = new_n8519_ & ~new_n36841_;
  assign new_n36843_ = ~new_n36674_ & new_n36842_;
  assign new_n36844_ = ~new_n36837_ & ~new_n36843_;
  assign new_n36845_ = ~\b[16]  & ~new_n36844_;
  assign new_n36846_ = ~new_n36395_ & ~new_n36675_;
  assign new_n36847_ = ~new_n36405_ & new_n36577_;
  assign new_n36848_ = ~new_n36573_ & new_n36847_;
  assign new_n36849_ = ~new_n36574_ & ~new_n36577_;
  assign new_n36850_ = ~new_n36848_ & ~new_n36849_;
  assign new_n36851_ = new_n8519_ & ~new_n36850_;
  assign new_n36852_ = ~new_n36674_ & new_n36851_;
  assign new_n36853_ = ~new_n36846_ & ~new_n36852_;
  assign new_n36854_ = ~\b[15]  & ~new_n36853_;
  assign new_n36855_ = ~new_n36404_ & ~new_n36675_;
  assign new_n36856_ = ~new_n36414_ & new_n36572_;
  assign new_n36857_ = ~new_n36568_ & new_n36856_;
  assign new_n36858_ = ~new_n36569_ & ~new_n36572_;
  assign new_n36859_ = ~new_n36857_ & ~new_n36858_;
  assign new_n36860_ = new_n8519_ & ~new_n36859_;
  assign new_n36861_ = ~new_n36674_ & new_n36860_;
  assign new_n36862_ = ~new_n36855_ & ~new_n36861_;
  assign new_n36863_ = ~\b[14]  & ~new_n36862_;
  assign new_n36864_ = ~new_n36413_ & ~new_n36675_;
  assign new_n36865_ = ~new_n36423_ & new_n36567_;
  assign new_n36866_ = ~new_n36563_ & new_n36865_;
  assign new_n36867_ = ~new_n36564_ & ~new_n36567_;
  assign new_n36868_ = ~new_n36866_ & ~new_n36867_;
  assign new_n36869_ = new_n8519_ & ~new_n36868_;
  assign new_n36870_ = ~new_n36674_ & new_n36869_;
  assign new_n36871_ = ~new_n36864_ & ~new_n36870_;
  assign new_n36872_ = ~\b[13]  & ~new_n36871_;
  assign new_n36873_ = ~new_n36422_ & ~new_n36675_;
  assign new_n36874_ = ~new_n36432_ & new_n36562_;
  assign new_n36875_ = ~new_n36558_ & new_n36874_;
  assign new_n36876_ = ~new_n36559_ & ~new_n36562_;
  assign new_n36877_ = ~new_n36875_ & ~new_n36876_;
  assign new_n36878_ = new_n8519_ & ~new_n36877_;
  assign new_n36879_ = ~new_n36674_ & new_n36878_;
  assign new_n36880_ = ~new_n36873_ & ~new_n36879_;
  assign new_n36881_ = ~\b[12]  & ~new_n36880_;
  assign new_n36882_ = ~new_n36431_ & ~new_n36675_;
  assign new_n36883_ = ~new_n36441_ & new_n36557_;
  assign new_n36884_ = ~new_n36553_ & new_n36883_;
  assign new_n36885_ = ~new_n36554_ & ~new_n36557_;
  assign new_n36886_ = ~new_n36884_ & ~new_n36885_;
  assign new_n36887_ = new_n8519_ & ~new_n36886_;
  assign new_n36888_ = ~new_n36674_ & new_n36887_;
  assign new_n36889_ = ~new_n36882_ & ~new_n36888_;
  assign new_n36890_ = ~\b[11]  & ~new_n36889_;
  assign new_n36891_ = ~new_n36440_ & ~new_n36675_;
  assign new_n36892_ = ~new_n36450_ & new_n36552_;
  assign new_n36893_ = ~new_n36548_ & new_n36892_;
  assign new_n36894_ = ~new_n36549_ & ~new_n36552_;
  assign new_n36895_ = ~new_n36893_ & ~new_n36894_;
  assign new_n36896_ = new_n8519_ & ~new_n36895_;
  assign new_n36897_ = ~new_n36674_ & new_n36896_;
  assign new_n36898_ = ~new_n36891_ & ~new_n36897_;
  assign new_n36899_ = ~\b[10]  & ~new_n36898_;
  assign new_n36900_ = ~new_n36449_ & ~new_n36675_;
  assign new_n36901_ = ~new_n36459_ & new_n36547_;
  assign new_n36902_ = ~new_n36543_ & new_n36901_;
  assign new_n36903_ = ~new_n36544_ & ~new_n36547_;
  assign new_n36904_ = ~new_n36902_ & ~new_n36903_;
  assign new_n36905_ = new_n8519_ & ~new_n36904_;
  assign new_n36906_ = ~new_n36674_ & new_n36905_;
  assign new_n36907_ = ~new_n36900_ & ~new_n36906_;
  assign new_n36908_ = ~\b[9]  & ~new_n36907_;
  assign new_n36909_ = ~new_n36458_ & ~new_n36675_;
  assign new_n36910_ = ~new_n36468_ & new_n36542_;
  assign new_n36911_ = ~new_n36538_ & new_n36910_;
  assign new_n36912_ = ~new_n36539_ & ~new_n36542_;
  assign new_n36913_ = ~new_n36911_ & ~new_n36912_;
  assign new_n36914_ = new_n8519_ & ~new_n36913_;
  assign new_n36915_ = ~new_n36674_ & new_n36914_;
  assign new_n36916_ = ~new_n36909_ & ~new_n36915_;
  assign new_n36917_ = ~\b[8]  & ~new_n36916_;
  assign new_n36918_ = ~new_n36467_ & ~new_n36675_;
  assign new_n36919_ = ~new_n36477_ & new_n36537_;
  assign new_n36920_ = ~new_n36533_ & new_n36919_;
  assign new_n36921_ = ~new_n36534_ & ~new_n36537_;
  assign new_n36922_ = ~new_n36920_ & ~new_n36921_;
  assign new_n36923_ = new_n8519_ & ~new_n36922_;
  assign new_n36924_ = ~new_n36674_ & new_n36923_;
  assign new_n36925_ = ~new_n36918_ & ~new_n36924_;
  assign new_n36926_ = ~\b[7]  & ~new_n36925_;
  assign new_n36927_ = ~new_n36476_ & ~new_n36675_;
  assign new_n36928_ = ~new_n36486_ & new_n36532_;
  assign new_n36929_ = ~new_n36528_ & new_n36928_;
  assign new_n36930_ = ~new_n36529_ & ~new_n36532_;
  assign new_n36931_ = ~new_n36929_ & ~new_n36930_;
  assign new_n36932_ = new_n8519_ & ~new_n36931_;
  assign new_n36933_ = ~new_n36674_ & new_n36932_;
  assign new_n36934_ = ~new_n36927_ & ~new_n36933_;
  assign new_n36935_ = ~\b[6]  & ~new_n36934_;
  assign new_n36936_ = ~new_n36485_ & ~new_n36675_;
  assign new_n36937_ = ~new_n36495_ & new_n36527_;
  assign new_n36938_ = ~new_n36523_ & new_n36937_;
  assign new_n36939_ = ~new_n36524_ & ~new_n36527_;
  assign new_n36940_ = ~new_n36938_ & ~new_n36939_;
  assign new_n36941_ = new_n8519_ & ~new_n36940_;
  assign new_n36942_ = ~new_n36674_ & new_n36941_;
  assign new_n36943_ = ~new_n36936_ & ~new_n36942_;
  assign new_n36944_ = ~\b[5]  & ~new_n36943_;
  assign new_n36945_ = ~new_n36494_ & ~new_n36675_;
  assign new_n36946_ = ~new_n36503_ & new_n36522_;
  assign new_n36947_ = ~new_n36518_ & new_n36946_;
  assign new_n36948_ = ~new_n36519_ & ~new_n36522_;
  assign new_n36949_ = ~new_n36947_ & ~new_n36948_;
  assign new_n36950_ = new_n8519_ & ~new_n36949_;
  assign new_n36951_ = ~new_n36674_ & new_n36950_;
  assign new_n36952_ = ~new_n36945_ & ~new_n36951_;
  assign new_n36953_ = ~\b[4]  & ~new_n36952_;
  assign new_n36954_ = ~new_n36502_ & ~new_n36675_;
  assign new_n36955_ = ~new_n36513_ & new_n36517_;
  assign new_n36956_ = ~new_n36512_ & new_n36955_;
  assign new_n36957_ = ~new_n36514_ & ~new_n36517_;
  assign new_n36958_ = ~new_n36956_ & ~new_n36957_;
  assign new_n36959_ = new_n8519_ & ~new_n36958_;
  assign new_n36960_ = ~new_n36674_ & new_n36959_;
  assign new_n36961_ = ~new_n36954_ & ~new_n36960_;
  assign new_n36962_ = ~\b[3]  & ~new_n36961_;
  assign new_n36963_ = ~new_n36507_ & ~new_n36675_;
  assign new_n36964_ = new_n8353_ & ~new_n36510_;
  assign new_n36965_ = ~new_n36508_ & new_n36964_;
  assign new_n36966_ = new_n8519_ & ~new_n36965_;
  assign new_n36967_ = ~new_n36512_ & new_n36966_;
  assign new_n36968_ = ~new_n36674_ & new_n36967_;
  assign new_n36969_ = ~new_n36963_ & ~new_n36968_;
  assign new_n36970_ = ~\b[2]  & ~new_n36969_;
  assign new_n36971_ = new_n8820_ & ~new_n36674_;
  assign new_n36972_ = \a[30]  & ~new_n36971_;
  assign new_n36973_ = new_n8826_ & ~new_n36674_;
  assign new_n36974_ = ~new_n36972_ & ~new_n36973_;
  assign new_n36975_ = \b[1]  & ~new_n36974_;
  assign new_n36976_ = ~\b[1]  & ~new_n36973_;
  assign new_n36977_ = ~new_n36972_ & new_n36976_;
  assign new_n36978_ = ~new_n36975_ & ~new_n36977_;
  assign new_n36979_ = ~new_n8833_ & ~new_n36978_;
  assign new_n36980_ = ~\b[1]  & ~new_n36974_;
  assign new_n36981_ = ~new_n36979_ & ~new_n36980_;
  assign new_n36982_ = \b[2]  & ~new_n36968_;
  assign new_n36983_ = ~new_n36963_ & new_n36982_;
  assign new_n36984_ = ~new_n36970_ & ~new_n36983_;
  assign new_n36985_ = ~new_n36981_ & new_n36984_;
  assign new_n36986_ = ~new_n36970_ & ~new_n36985_;
  assign new_n36987_ = \b[3]  & ~new_n36960_;
  assign new_n36988_ = ~new_n36954_ & new_n36987_;
  assign new_n36989_ = ~new_n36962_ & ~new_n36988_;
  assign new_n36990_ = ~new_n36986_ & new_n36989_;
  assign new_n36991_ = ~new_n36962_ & ~new_n36990_;
  assign new_n36992_ = \b[4]  & ~new_n36951_;
  assign new_n36993_ = ~new_n36945_ & new_n36992_;
  assign new_n36994_ = ~new_n36953_ & ~new_n36993_;
  assign new_n36995_ = ~new_n36991_ & new_n36994_;
  assign new_n36996_ = ~new_n36953_ & ~new_n36995_;
  assign new_n36997_ = \b[5]  & ~new_n36942_;
  assign new_n36998_ = ~new_n36936_ & new_n36997_;
  assign new_n36999_ = ~new_n36944_ & ~new_n36998_;
  assign new_n37000_ = ~new_n36996_ & new_n36999_;
  assign new_n37001_ = ~new_n36944_ & ~new_n37000_;
  assign new_n37002_ = \b[6]  & ~new_n36933_;
  assign new_n37003_ = ~new_n36927_ & new_n37002_;
  assign new_n37004_ = ~new_n36935_ & ~new_n37003_;
  assign new_n37005_ = ~new_n37001_ & new_n37004_;
  assign new_n37006_ = ~new_n36935_ & ~new_n37005_;
  assign new_n37007_ = \b[7]  & ~new_n36924_;
  assign new_n37008_ = ~new_n36918_ & new_n37007_;
  assign new_n37009_ = ~new_n36926_ & ~new_n37008_;
  assign new_n37010_ = ~new_n37006_ & new_n37009_;
  assign new_n37011_ = ~new_n36926_ & ~new_n37010_;
  assign new_n37012_ = \b[8]  & ~new_n36915_;
  assign new_n37013_ = ~new_n36909_ & new_n37012_;
  assign new_n37014_ = ~new_n36917_ & ~new_n37013_;
  assign new_n37015_ = ~new_n37011_ & new_n37014_;
  assign new_n37016_ = ~new_n36917_ & ~new_n37015_;
  assign new_n37017_ = \b[9]  & ~new_n36906_;
  assign new_n37018_ = ~new_n36900_ & new_n37017_;
  assign new_n37019_ = ~new_n36908_ & ~new_n37018_;
  assign new_n37020_ = ~new_n37016_ & new_n37019_;
  assign new_n37021_ = ~new_n36908_ & ~new_n37020_;
  assign new_n37022_ = \b[10]  & ~new_n36897_;
  assign new_n37023_ = ~new_n36891_ & new_n37022_;
  assign new_n37024_ = ~new_n36899_ & ~new_n37023_;
  assign new_n37025_ = ~new_n37021_ & new_n37024_;
  assign new_n37026_ = ~new_n36899_ & ~new_n37025_;
  assign new_n37027_ = \b[11]  & ~new_n36888_;
  assign new_n37028_ = ~new_n36882_ & new_n37027_;
  assign new_n37029_ = ~new_n36890_ & ~new_n37028_;
  assign new_n37030_ = ~new_n37026_ & new_n37029_;
  assign new_n37031_ = ~new_n36890_ & ~new_n37030_;
  assign new_n37032_ = \b[12]  & ~new_n36879_;
  assign new_n37033_ = ~new_n36873_ & new_n37032_;
  assign new_n37034_ = ~new_n36881_ & ~new_n37033_;
  assign new_n37035_ = ~new_n37031_ & new_n37034_;
  assign new_n37036_ = ~new_n36881_ & ~new_n37035_;
  assign new_n37037_ = \b[13]  & ~new_n36870_;
  assign new_n37038_ = ~new_n36864_ & new_n37037_;
  assign new_n37039_ = ~new_n36872_ & ~new_n37038_;
  assign new_n37040_ = ~new_n37036_ & new_n37039_;
  assign new_n37041_ = ~new_n36872_ & ~new_n37040_;
  assign new_n37042_ = \b[14]  & ~new_n36861_;
  assign new_n37043_ = ~new_n36855_ & new_n37042_;
  assign new_n37044_ = ~new_n36863_ & ~new_n37043_;
  assign new_n37045_ = ~new_n37041_ & new_n37044_;
  assign new_n37046_ = ~new_n36863_ & ~new_n37045_;
  assign new_n37047_ = \b[15]  & ~new_n36852_;
  assign new_n37048_ = ~new_n36846_ & new_n37047_;
  assign new_n37049_ = ~new_n36854_ & ~new_n37048_;
  assign new_n37050_ = ~new_n37046_ & new_n37049_;
  assign new_n37051_ = ~new_n36854_ & ~new_n37050_;
  assign new_n37052_ = \b[16]  & ~new_n36843_;
  assign new_n37053_ = ~new_n36837_ & new_n37052_;
  assign new_n37054_ = ~new_n36845_ & ~new_n37053_;
  assign new_n37055_ = ~new_n37051_ & new_n37054_;
  assign new_n37056_ = ~new_n36845_ & ~new_n37055_;
  assign new_n37057_ = \b[17]  & ~new_n36834_;
  assign new_n37058_ = ~new_n36828_ & new_n37057_;
  assign new_n37059_ = ~new_n36836_ & ~new_n37058_;
  assign new_n37060_ = ~new_n37056_ & new_n37059_;
  assign new_n37061_ = ~new_n36836_ & ~new_n37060_;
  assign new_n37062_ = \b[18]  & ~new_n36825_;
  assign new_n37063_ = ~new_n36819_ & new_n37062_;
  assign new_n37064_ = ~new_n36827_ & ~new_n37063_;
  assign new_n37065_ = ~new_n37061_ & new_n37064_;
  assign new_n37066_ = ~new_n36827_ & ~new_n37065_;
  assign new_n37067_ = \b[19]  & ~new_n36816_;
  assign new_n37068_ = ~new_n36810_ & new_n37067_;
  assign new_n37069_ = ~new_n36818_ & ~new_n37068_;
  assign new_n37070_ = ~new_n37066_ & new_n37069_;
  assign new_n37071_ = ~new_n36818_ & ~new_n37070_;
  assign new_n37072_ = \b[20]  & ~new_n36807_;
  assign new_n37073_ = ~new_n36801_ & new_n37072_;
  assign new_n37074_ = ~new_n36809_ & ~new_n37073_;
  assign new_n37075_ = ~new_n37071_ & new_n37074_;
  assign new_n37076_ = ~new_n36809_ & ~new_n37075_;
  assign new_n37077_ = \b[21]  & ~new_n36798_;
  assign new_n37078_ = ~new_n36792_ & new_n37077_;
  assign new_n37079_ = ~new_n36800_ & ~new_n37078_;
  assign new_n37080_ = ~new_n37076_ & new_n37079_;
  assign new_n37081_ = ~new_n36800_ & ~new_n37080_;
  assign new_n37082_ = \b[22]  & ~new_n36789_;
  assign new_n37083_ = ~new_n36783_ & new_n37082_;
  assign new_n37084_ = ~new_n36791_ & ~new_n37083_;
  assign new_n37085_ = ~new_n37081_ & new_n37084_;
  assign new_n37086_ = ~new_n36791_ & ~new_n37085_;
  assign new_n37087_ = \b[23]  & ~new_n36780_;
  assign new_n37088_ = ~new_n36774_ & new_n37087_;
  assign new_n37089_ = ~new_n36782_ & ~new_n37088_;
  assign new_n37090_ = ~new_n37086_ & new_n37089_;
  assign new_n37091_ = ~new_n36782_ & ~new_n37090_;
  assign new_n37092_ = \b[24]  & ~new_n36771_;
  assign new_n37093_ = ~new_n36765_ & new_n37092_;
  assign new_n37094_ = ~new_n36773_ & ~new_n37093_;
  assign new_n37095_ = ~new_n37091_ & new_n37094_;
  assign new_n37096_ = ~new_n36773_ & ~new_n37095_;
  assign new_n37097_ = \b[25]  & ~new_n36762_;
  assign new_n37098_ = ~new_n36756_ & new_n37097_;
  assign new_n37099_ = ~new_n36764_ & ~new_n37098_;
  assign new_n37100_ = ~new_n37096_ & new_n37099_;
  assign new_n37101_ = ~new_n36764_ & ~new_n37100_;
  assign new_n37102_ = \b[26]  & ~new_n36753_;
  assign new_n37103_ = ~new_n36747_ & new_n37102_;
  assign new_n37104_ = ~new_n36755_ & ~new_n37103_;
  assign new_n37105_ = ~new_n37101_ & new_n37104_;
  assign new_n37106_ = ~new_n36755_ & ~new_n37105_;
  assign new_n37107_ = \b[27]  & ~new_n36744_;
  assign new_n37108_ = ~new_n36738_ & new_n37107_;
  assign new_n37109_ = ~new_n36746_ & ~new_n37108_;
  assign new_n37110_ = ~new_n37106_ & new_n37109_;
  assign new_n37111_ = ~new_n36746_ & ~new_n37110_;
  assign new_n37112_ = \b[28]  & ~new_n36735_;
  assign new_n37113_ = ~new_n36729_ & new_n37112_;
  assign new_n37114_ = ~new_n36737_ & ~new_n37113_;
  assign new_n37115_ = ~new_n37111_ & new_n37114_;
  assign new_n37116_ = ~new_n36737_ & ~new_n37115_;
  assign new_n37117_ = \b[29]  & ~new_n36726_;
  assign new_n37118_ = ~new_n36720_ & new_n37117_;
  assign new_n37119_ = ~new_n36728_ & ~new_n37118_;
  assign new_n37120_ = ~new_n37116_ & new_n37119_;
  assign new_n37121_ = ~new_n36728_ & ~new_n37120_;
  assign new_n37122_ = \b[30]  & ~new_n36717_;
  assign new_n37123_ = ~new_n36711_ & new_n37122_;
  assign new_n37124_ = ~new_n36719_ & ~new_n37123_;
  assign new_n37125_ = ~new_n37121_ & new_n37124_;
  assign new_n37126_ = ~new_n36719_ & ~new_n37125_;
  assign new_n37127_ = \b[31]  & ~new_n36708_;
  assign new_n37128_ = ~new_n36702_ & new_n37127_;
  assign new_n37129_ = ~new_n36710_ & ~new_n37128_;
  assign new_n37130_ = ~new_n37126_ & new_n37129_;
  assign new_n37131_ = ~new_n36710_ & ~new_n37130_;
  assign new_n37132_ = \b[32]  & ~new_n36699_;
  assign new_n37133_ = ~new_n36693_ & new_n37132_;
  assign new_n37134_ = ~new_n36701_ & ~new_n37133_;
  assign new_n37135_ = ~new_n37131_ & new_n37134_;
  assign new_n37136_ = ~new_n36701_ & ~new_n37135_;
  assign new_n37137_ = \b[33]  & ~new_n36682_;
  assign new_n37138_ = ~new_n36676_ & new_n37137_;
  assign new_n37139_ = ~new_n36692_ & ~new_n37138_;
  assign new_n37140_ = ~new_n37136_ & new_n37139_;
  assign new_n37141_ = ~new_n36692_ & ~new_n37140_;
  assign new_n37142_ = \b[34]  & ~new_n36684_;
  assign new_n37143_ = ~new_n36689_ & new_n37142_;
  assign new_n37144_ = ~new_n36691_ & ~new_n37143_;
  assign new_n37145_ = ~new_n37141_ & new_n37144_;
  assign new_n37146_ = ~new_n36691_ & ~new_n37145_;
  assign new_n37147_ = new_n9004_ & ~new_n37146_;
  assign new_n37148_ = ~new_n36683_ & ~new_n37147_;
  assign new_n37149_ = ~new_n36701_ & new_n37139_;
  assign new_n37150_ = ~new_n37135_ & new_n37149_;
  assign new_n37151_ = ~new_n37136_ & ~new_n37139_;
  assign new_n37152_ = ~new_n37150_ & ~new_n37151_;
  assign new_n37153_ = new_n9004_ & ~new_n37152_;
  assign new_n37154_ = ~new_n37146_ & new_n37153_;
  assign new_n37155_ = ~new_n37148_ & ~new_n37154_;
  assign new_n37156_ = ~\b[34]  & ~new_n37155_;
  assign new_n37157_ = ~new_n36700_ & ~new_n37147_;
  assign new_n37158_ = ~new_n36710_ & new_n37134_;
  assign new_n37159_ = ~new_n37130_ & new_n37158_;
  assign new_n37160_ = ~new_n37131_ & ~new_n37134_;
  assign new_n37161_ = ~new_n37159_ & ~new_n37160_;
  assign new_n37162_ = new_n9004_ & ~new_n37161_;
  assign new_n37163_ = ~new_n37146_ & new_n37162_;
  assign new_n37164_ = ~new_n37157_ & ~new_n37163_;
  assign new_n37165_ = ~\b[33]  & ~new_n37164_;
  assign new_n37166_ = ~new_n36709_ & ~new_n37147_;
  assign new_n37167_ = ~new_n36719_ & new_n37129_;
  assign new_n37168_ = ~new_n37125_ & new_n37167_;
  assign new_n37169_ = ~new_n37126_ & ~new_n37129_;
  assign new_n37170_ = ~new_n37168_ & ~new_n37169_;
  assign new_n37171_ = new_n9004_ & ~new_n37170_;
  assign new_n37172_ = ~new_n37146_ & new_n37171_;
  assign new_n37173_ = ~new_n37166_ & ~new_n37172_;
  assign new_n37174_ = ~\b[32]  & ~new_n37173_;
  assign new_n37175_ = ~new_n36718_ & ~new_n37147_;
  assign new_n37176_ = ~new_n36728_ & new_n37124_;
  assign new_n37177_ = ~new_n37120_ & new_n37176_;
  assign new_n37178_ = ~new_n37121_ & ~new_n37124_;
  assign new_n37179_ = ~new_n37177_ & ~new_n37178_;
  assign new_n37180_ = new_n9004_ & ~new_n37179_;
  assign new_n37181_ = ~new_n37146_ & new_n37180_;
  assign new_n37182_ = ~new_n37175_ & ~new_n37181_;
  assign new_n37183_ = ~\b[31]  & ~new_n37182_;
  assign new_n37184_ = ~new_n36727_ & ~new_n37147_;
  assign new_n37185_ = ~new_n36737_ & new_n37119_;
  assign new_n37186_ = ~new_n37115_ & new_n37185_;
  assign new_n37187_ = ~new_n37116_ & ~new_n37119_;
  assign new_n37188_ = ~new_n37186_ & ~new_n37187_;
  assign new_n37189_ = new_n9004_ & ~new_n37188_;
  assign new_n37190_ = ~new_n37146_ & new_n37189_;
  assign new_n37191_ = ~new_n37184_ & ~new_n37190_;
  assign new_n37192_ = ~\b[30]  & ~new_n37191_;
  assign new_n37193_ = ~new_n36736_ & ~new_n37147_;
  assign new_n37194_ = ~new_n36746_ & new_n37114_;
  assign new_n37195_ = ~new_n37110_ & new_n37194_;
  assign new_n37196_ = ~new_n37111_ & ~new_n37114_;
  assign new_n37197_ = ~new_n37195_ & ~new_n37196_;
  assign new_n37198_ = new_n9004_ & ~new_n37197_;
  assign new_n37199_ = ~new_n37146_ & new_n37198_;
  assign new_n37200_ = ~new_n37193_ & ~new_n37199_;
  assign new_n37201_ = ~\b[29]  & ~new_n37200_;
  assign new_n37202_ = ~new_n36745_ & ~new_n37147_;
  assign new_n37203_ = ~new_n36755_ & new_n37109_;
  assign new_n37204_ = ~new_n37105_ & new_n37203_;
  assign new_n37205_ = ~new_n37106_ & ~new_n37109_;
  assign new_n37206_ = ~new_n37204_ & ~new_n37205_;
  assign new_n37207_ = new_n9004_ & ~new_n37206_;
  assign new_n37208_ = ~new_n37146_ & new_n37207_;
  assign new_n37209_ = ~new_n37202_ & ~new_n37208_;
  assign new_n37210_ = ~\b[28]  & ~new_n37209_;
  assign new_n37211_ = ~new_n36754_ & ~new_n37147_;
  assign new_n37212_ = ~new_n36764_ & new_n37104_;
  assign new_n37213_ = ~new_n37100_ & new_n37212_;
  assign new_n37214_ = ~new_n37101_ & ~new_n37104_;
  assign new_n37215_ = ~new_n37213_ & ~new_n37214_;
  assign new_n37216_ = new_n9004_ & ~new_n37215_;
  assign new_n37217_ = ~new_n37146_ & new_n37216_;
  assign new_n37218_ = ~new_n37211_ & ~new_n37217_;
  assign new_n37219_ = ~\b[27]  & ~new_n37218_;
  assign new_n37220_ = ~new_n36763_ & ~new_n37147_;
  assign new_n37221_ = ~new_n36773_ & new_n37099_;
  assign new_n37222_ = ~new_n37095_ & new_n37221_;
  assign new_n37223_ = ~new_n37096_ & ~new_n37099_;
  assign new_n37224_ = ~new_n37222_ & ~new_n37223_;
  assign new_n37225_ = new_n9004_ & ~new_n37224_;
  assign new_n37226_ = ~new_n37146_ & new_n37225_;
  assign new_n37227_ = ~new_n37220_ & ~new_n37226_;
  assign new_n37228_ = ~\b[26]  & ~new_n37227_;
  assign new_n37229_ = ~new_n36772_ & ~new_n37147_;
  assign new_n37230_ = ~new_n36782_ & new_n37094_;
  assign new_n37231_ = ~new_n37090_ & new_n37230_;
  assign new_n37232_ = ~new_n37091_ & ~new_n37094_;
  assign new_n37233_ = ~new_n37231_ & ~new_n37232_;
  assign new_n37234_ = new_n9004_ & ~new_n37233_;
  assign new_n37235_ = ~new_n37146_ & new_n37234_;
  assign new_n37236_ = ~new_n37229_ & ~new_n37235_;
  assign new_n37237_ = ~\b[25]  & ~new_n37236_;
  assign new_n37238_ = ~new_n36781_ & ~new_n37147_;
  assign new_n37239_ = ~new_n36791_ & new_n37089_;
  assign new_n37240_ = ~new_n37085_ & new_n37239_;
  assign new_n37241_ = ~new_n37086_ & ~new_n37089_;
  assign new_n37242_ = ~new_n37240_ & ~new_n37241_;
  assign new_n37243_ = new_n9004_ & ~new_n37242_;
  assign new_n37244_ = ~new_n37146_ & new_n37243_;
  assign new_n37245_ = ~new_n37238_ & ~new_n37244_;
  assign new_n37246_ = ~\b[24]  & ~new_n37245_;
  assign new_n37247_ = ~new_n36790_ & ~new_n37147_;
  assign new_n37248_ = ~new_n36800_ & new_n37084_;
  assign new_n37249_ = ~new_n37080_ & new_n37248_;
  assign new_n37250_ = ~new_n37081_ & ~new_n37084_;
  assign new_n37251_ = ~new_n37249_ & ~new_n37250_;
  assign new_n37252_ = new_n9004_ & ~new_n37251_;
  assign new_n37253_ = ~new_n37146_ & new_n37252_;
  assign new_n37254_ = ~new_n37247_ & ~new_n37253_;
  assign new_n37255_ = ~\b[23]  & ~new_n37254_;
  assign new_n37256_ = ~new_n36799_ & ~new_n37147_;
  assign new_n37257_ = ~new_n36809_ & new_n37079_;
  assign new_n37258_ = ~new_n37075_ & new_n37257_;
  assign new_n37259_ = ~new_n37076_ & ~new_n37079_;
  assign new_n37260_ = ~new_n37258_ & ~new_n37259_;
  assign new_n37261_ = new_n9004_ & ~new_n37260_;
  assign new_n37262_ = ~new_n37146_ & new_n37261_;
  assign new_n37263_ = ~new_n37256_ & ~new_n37262_;
  assign new_n37264_ = ~\b[22]  & ~new_n37263_;
  assign new_n37265_ = ~new_n36808_ & ~new_n37147_;
  assign new_n37266_ = ~new_n36818_ & new_n37074_;
  assign new_n37267_ = ~new_n37070_ & new_n37266_;
  assign new_n37268_ = ~new_n37071_ & ~new_n37074_;
  assign new_n37269_ = ~new_n37267_ & ~new_n37268_;
  assign new_n37270_ = new_n9004_ & ~new_n37269_;
  assign new_n37271_ = ~new_n37146_ & new_n37270_;
  assign new_n37272_ = ~new_n37265_ & ~new_n37271_;
  assign new_n37273_ = ~\b[21]  & ~new_n37272_;
  assign new_n37274_ = ~new_n36817_ & ~new_n37147_;
  assign new_n37275_ = ~new_n36827_ & new_n37069_;
  assign new_n37276_ = ~new_n37065_ & new_n37275_;
  assign new_n37277_ = ~new_n37066_ & ~new_n37069_;
  assign new_n37278_ = ~new_n37276_ & ~new_n37277_;
  assign new_n37279_ = new_n9004_ & ~new_n37278_;
  assign new_n37280_ = ~new_n37146_ & new_n37279_;
  assign new_n37281_ = ~new_n37274_ & ~new_n37280_;
  assign new_n37282_ = ~\b[20]  & ~new_n37281_;
  assign new_n37283_ = ~new_n36826_ & ~new_n37147_;
  assign new_n37284_ = ~new_n36836_ & new_n37064_;
  assign new_n37285_ = ~new_n37060_ & new_n37284_;
  assign new_n37286_ = ~new_n37061_ & ~new_n37064_;
  assign new_n37287_ = ~new_n37285_ & ~new_n37286_;
  assign new_n37288_ = new_n9004_ & ~new_n37287_;
  assign new_n37289_ = ~new_n37146_ & new_n37288_;
  assign new_n37290_ = ~new_n37283_ & ~new_n37289_;
  assign new_n37291_ = ~\b[19]  & ~new_n37290_;
  assign new_n37292_ = ~new_n36835_ & ~new_n37147_;
  assign new_n37293_ = ~new_n36845_ & new_n37059_;
  assign new_n37294_ = ~new_n37055_ & new_n37293_;
  assign new_n37295_ = ~new_n37056_ & ~new_n37059_;
  assign new_n37296_ = ~new_n37294_ & ~new_n37295_;
  assign new_n37297_ = new_n9004_ & ~new_n37296_;
  assign new_n37298_ = ~new_n37146_ & new_n37297_;
  assign new_n37299_ = ~new_n37292_ & ~new_n37298_;
  assign new_n37300_ = ~\b[18]  & ~new_n37299_;
  assign new_n37301_ = ~new_n36844_ & ~new_n37147_;
  assign new_n37302_ = ~new_n36854_ & new_n37054_;
  assign new_n37303_ = ~new_n37050_ & new_n37302_;
  assign new_n37304_ = ~new_n37051_ & ~new_n37054_;
  assign new_n37305_ = ~new_n37303_ & ~new_n37304_;
  assign new_n37306_ = new_n9004_ & ~new_n37305_;
  assign new_n37307_ = ~new_n37146_ & new_n37306_;
  assign new_n37308_ = ~new_n37301_ & ~new_n37307_;
  assign new_n37309_ = ~\b[17]  & ~new_n37308_;
  assign new_n37310_ = ~new_n36853_ & ~new_n37147_;
  assign new_n37311_ = ~new_n36863_ & new_n37049_;
  assign new_n37312_ = ~new_n37045_ & new_n37311_;
  assign new_n37313_ = ~new_n37046_ & ~new_n37049_;
  assign new_n37314_ = ~new_n37312_ & ~new_n37313_;
  assign new_n37315_ = new_n9004_ & ~new_n37314_;
  assign new_n37316_ = ~new_n37146_ & new_n37315_;
  assign new_n37317_ = ~new_n37310_ & ~new_n37316_;
  assign new_n37318_ = ~\b[16]  & ~new_n37317_;
  assign new_n37319_ = ~new_n36862_ & ~new_n37147_;
  assign new_n37320_ = ~new_n36872_ & new_n37044_;
  assign new_n37321_ = ~new_n37040_ & new_n37320_;
  assign new_n37322_ = ~new_n37041_ & ~new_n37044_;
  assign new_n37323_ = ~new_n37321_ & ~new_n37322_;
  assign new_n37324_ = new_n9004_ & ~new_n37323_;
  assign new_n37325_ = ~new_n37146_ & new_n37324_;
  assign new_n37326_ = ~new_n37319_ & ~new_n37325_;
  assign new_n37327_ = ~\b[15]  & ~new_n37326_;
  assign new_n37328_ = ~new_n36871_ & ~new_n37147_;
  assign new_n37329_ = ~new_n36881_ & new_n37039_;
  assign new_n37330_ = ~new_n37035_ & new_n37329_;
  assign new_n37331_ = ~new_n37036_ & ~new_n37039_;
  assign new_n37332_ = ~new_n37330_ & ~new_n37331_;
  assign new_n37333_ = new_n9004_ & ~new_n37332_;
  assign new_n37334_ = ~new_n37146_ & new_n37333_;
  assign new_n37335_ = ~new_n37328_ & ~new_n37334_;
  assign new_n37336_ = ~\b[14]  & ~new_n37335_;
  assign new_n37337_ = ~new_n36880_ & ~new_n37147_;
  assign new_n37338_ = ~new_n36890_ & new_n37034_;
  assign new_n37339_ = ~new_n37030_ & new_n37338_;
  assign new_n37340_ = ~new_n37031_ & ~new_n37034_;
  assign new_n37341_ = ~new_n37339_ & ~new_n37340_;
  assign new_n37342_ = new_n9004_ & ~new_n37341_;
  assign new_n37343_ = ~new_n37146_ & new_n37342_;
  assign new_n37344_ = ~new_n37337_ & ~new_n37343_;
  assign new_n37345_ = ~\b[13]  & ~new_n37344_;
  assign new_n37346_ = ~new_n36889_ & ~new_n37147_;
  assign new_n37347_ = ~new_n36899_ & new_n37029_;
  assign new_n37348_ = ~new_n37025_ & new_n37347_;
  assign new_n37349_ = ~new_n37026_ & ~new_n37029_;
  assign new_n37350_ = ~new_n37348_ & ~new_n37349_;
  assign new_n37351_ = new_n9004_ & ~new_n37350_;
  assign new_n37352_ = ~new_n37146_ & new_n37351_;
  assign new_n37353_ = ~new_n37346_ & ~new_n37352_;
  assign new_n37354_ = ~\b[12]  & ~new_n37353_;
  assign new_n37355_ = ~new_n36898_ & ~new_n37147_;
  assign new_n37356_ = ~new_n36908_ & new_n37024_;
  assign new_n37357_ = ~new_n37020_ & new_n37356_;
  assign new_n37358_ = ~new_n37021_ & ~new_n37024_;
  assign new_n37359_ = ~new_n37357_ & ~new_n37358_;
  assign new_n37360_ = new_n9004_ & ~new_n37359_;
  assign new_n37361_ = ~new_n37146_ & new_n37360_;
  assign new_n37362_ = ~new_n37355_ & ~new_n37361_;
  assign new_n37363_ = ~\b[11]  & ~new_n37362_;
  assign new_n37364_ = ~new_n36907_ & ~new_n37147_;
  assign new_n37365_ = ~new_n36917_ & new_n37019_;
  assign new_n37366_ = ~new_n37015_ & new_n37365_;
  assign new_n37367_ = ~new_n37016_ & ~new_n37019_;
  assign new_n37368_ = ~new_n37366_ & ~new_n37367_;
  assign new_n37369_ = new_n9004_ & ~new_n37368_;
  assign new_n37370_ = ~new_n37146_ & new_n37369_;
  assign new_n37371_ = ~new_n37364_ & ~new_n37370_;
  assign new_n37372_ = ~\b[10]  & ~new_n37371_;
  assign new_n37373_ = ~new_n36916_ & ~new_n37147_;
  assign new_n37374_ = ~new_n36926_ & new_n37014_;
  assign new_n37375_ = ~new_n37010_ & new_n37374_;
  assign new_n37376_ = ~new_n37011_ & ~new_n37014_;
  assign new_n37377_ = ~new_n37375_ & ~new_n37376_;
  assign new_n37378_ = new_n9004_ & ~new_n37377_;
  assign new_n37379_ = ~new_n37146_ & new_n37378_;
  assign new_n37380_ = ~new_n37373_ & ~new_n37379_;
  assign new_n37381_ = ~\b[9]  & ~new_n37380_;
  assign new_n37382_ = ~new_n36925_ & ~new_n37147_;
  assign new_n37383_ = ~new_n36935_ & new_n37009_;
  assign new_n37384_ = ~new_n37005_ & new_n37383_;
  assign new_n37385_ = ~new_n37006_ & ~new_n37009_;
  assign new_n37386_ = ~new_n37384_ & ~new_n37385_;
  assign new_n37387_ = new_n9004_ & ~new_n37386_;
  assign new_n37388_ = ~new_n37146_ & new_n37387_;
  assign new_n37389_ = ~new_n37382_ & ~new_n37388_;
  assign new_n37390_ = ~\b[8]  & ~new_n37389_;
  assign new_n37391_ = ~new_n36934_ & ~new_n37147_;
  assign new_n37392_ = ~new_n36944_ & new_n37004_;
  assign new_n37393_ = ~new_n37000_ & new_n37392_;
  assign new_n37394_ = ~new_n37001_ & ~new_n37004_;
  assign new_n37395_ = ~new_n37393_ & ~new_n37394_;
  assign new_n37396_ = new_n9004_ & ~new_n37395_;
  assign new_n37397_ = ~new_n37146_ & new_n37396_;
  assign new_n37398_ = ~new_n37391_ & ~new_n37397_;
  assign new_n37399_ = ~\b[7]  & ~new_n37398_;
  assign new_n37400_ = ~new_n36943_ & ~new_n37147_;
  assign new_n37401_ = ~new_n36953_ & new_n36999_;
  assign new_n37402_ = ~new_n36995_ & new_n37401_;
  assign new_n37403_ = ~new_n36996_ & ~new_n36999_;
  assign new_n37404_ = ~new_n37402_ & ~new_n37403_;
  assign new_n37405_ = new_n9004_ & ~new_n37404_;
  assign new_n37406_ = ~new_n37146_ & new_n37405_;
  assign new_n37407_ = ~new_n37400_ & ~new_n37406_;
  assign new_n37408_ = ~\b[6]  & ~new_n37407_;
  assign new_n37409_ = ~new_n36952_ & ~new_n37147_;
  assign new_n37410_ = ~new_n36962_ & new_n36994_;
  assign new_n37411_ = ~new_n36990_ & new_n37410_;
  assign new_n37412_ = ~new_n36991_ & ~new_n36994_;
  assign new_n37413_ = ~new_n37411_ & ~new_n37412_;
  assign new_n37414_ = new_n9004_ & ~new_n37413_;
  assign new_n37415_ = ~new_n37146_ & new_n37414_;
  assign new_n37416_ = ~new_n37409_ & ~new_n37415_;
  assign new_n37417_ = ~\b[5]  & ~new_n37416_;
  assign new_n37418_ = ~new_n36961_ & ~new_n37147_;
  assign new_n37419_ = ~new_n36970_ & new_n36989_;
  assign new_n37420_ = ~new_n36985_ & new_n37419_;
  assign new_n37421_ = ~new_n36986_ & ~new_n36989_;
  assign new_n37422_ = ~new_n37420_ & ~new_n37421_;
  assign new_n37423_ = new_n9004_ & ~new_n37422_;
  assign new_n37424_ = ~new_n37146_ & new_n37423_;
  assign new_n37425_ = ~new_n37418_ & ~new_n37424_;
  assign new_n37426_ = ~\b[4]  & ~new_n37425_;
  assign new_n37427_ = ~new_n36969_ & ~new_n37147_;
  assign new_n37428_ = ~new_n36980_ & new_n36984_;
  assign new_n37429_ = ~new_n36979_ & new_n37428_;
  assign new_n37430_ = ~new_n36981_ & ~new_n36984_;
  assign new_n37431_ = ~new_n37429_ & ~new_n37430_;
  assign new_n37432_ = new_n9004_ & ~new_n37431_;
  assign new_n37433_ = ~new_n37146_ & new_n37432_;
  assign new_n37434_ = ~new_n37427_ & ~new_n37433_;
  assign new_n37435_ = ~\b[3]  & ~new_n37434_;
  assign new_n37436_ = ~new_n36974_ & ~new_n37147_;
  assign new_n37437_ = new_n8833_ & ~new_n36977_;
  assign new_n37438_ = ~new_n36975_ & new_n37437_;
  assign new_n37439_ = new_n9004_ & ~new_n37438_;
  assign new_n37440_ = ~new_n36979_ & new_n37439_;
  assign new_n37441_ = ~new_n37146_ & new_n37440_;
  assign new_n37442_ = ~new_n37436_ & ~new_n37441_;
  assign new_n37443_ = ~\b[2]  & ~new_n37442_;
  assign new_n37444_ = new_n9305_ & ~new_n37146_;
  assign new_n37445_ = \a[29]  & ~new_n37444_;
  assign new_n37446_ = new_n9311_ & ~new_n37146_;
  assign new_n37447_ = ~new_n37445_ & ~new_n37446_;
  assign new_n37448_ = \b[1]  & ~new_n37447_;
  assign new_n37449_ = ~\b[1]  & ~new_n37446_;
  assign new_n37450_ = ~new_n37445_ & new_n37449_;
  assign new_n37451_ = ~new_n37448_ & ~new_n37450_;
  assign new_n37452_ = ~new_n9318_ & ~new_n37451_;
  assign new_n37453_ = ~\b[1]  & ~new_n37447_;
  assign new_n37454_ = ~new_n37452_ & ~new_n37453_;
  assign new_n37455_ = \b[2]  & ~new_n37441_;
  assign new_n37456_ = ~new_n37436_ & new_n37455_;
  assign new_n37457_ = ~new_n37443_ & ~new_n37456_;
  assign new_n37458_ = ~new_n37454_ & new_n37457_;
  assign new_n37459_ = ~new_n37443_ & ~new_n37458_;
  assign new_n37460_ = \b[3]  & ~new_n37433_;
  assign new_n37461_ = ~new_n37427_ & new_n37460_;
  assign new_n37462_ = ~new_n37435_ & ~new_n37461_;
  assign new_n37463_ = ~new_n37459_ & new_n37462_;
  assign new_n37464_ = ~new_n37435_ & ~new_n37463_;
  assign new_n37465_ = \b[4]  & ~new_n37424_;
  assign new_n37466_ = ~new_n37418_ & new_n37465_;
  assign new_n37467_ = ~new_n37426_ & ~new_n37466_;
  assign new_n37468_ = ~new_n37464_ & new_n37467_;
  assign new_n37469_ = ~new_n37426_ & ~new_n37468_;
  assign new_n37470_ = \b[5]  & ~new_n37415_;
  assign new_n37471_ = ~new_n37409_ & new_n37470_;
  assign new_n37472_ = ~new_n37417_ & ~new_n37471_;
  assign new_n37473_ = ~new_n37469_ & new_n37472_;
  assign new_n37474_ = ~new_n37417_ & ~new_n37473_;
  assign new_n37475_ = \b[6]  & ~new_n37406_;
  assign new_n37476_ = ~new_n37400_ & new_n37475_;
  assign new_n37477_ = ~new_n37408_ & ~new_n37476_;
  assign new_n37478_ = ~new_n37474_ & new_n37477_;
  assign new_n37479_ = ~new_n37408_ & ~new_n37478_;
  assign new_n37480_ = \b[7]  & ~new_n37397_;
  assign new_n37481_ = ~new_n37391_ & new_n37480_;
  assign new_n37482_ = ~new_n37399_ & ~new_n37481_;
  assign new_n37483_ = ~new_n37479_ & new_n37482_;
  assign new_n37484_ = ~new_n37399_ & ~new_n37483_;
  assign new_n37485_ = \b[8]  & ~new_n37388_;
  assign new_n37486_ = ~new_n37382_ & new_n37485_;
  assign new_n37487_ = ~new_n37390_ & ~new_n37486_;
  assign new_n37488_ = ~new_n37484_ & new_n37487_;
  assign new_n37489_ = ~new_n37390_ & ~new_n37488_;
  assign new_n37490_ = \b[9]  & ~new_n37379_;
  assign new_n37491_ = ~new_n37373_ & new_n37490_;
  assign new_n37492_ = ~new_n37381_ & ~new_n37491_;
  assign new_n37493_ = ~new_n37489_ & new_n37492_;
  assign new_n37494_ = ~new_n37381_ & ~new_n37493_;
  assign new_n37495_ = \b[10]  & ~new_n37370_;
  assign new_n37496_ = ~new_n37364_ & new_n37495_;
  assign new_n37497_ = ~new_n37372_ & ~new_n37496_;
  assign new_n37498_ = ~new_n37494_ & new_n37497_;
  assign new_n37499_ = ~new_n37372_ & ~new_n37498_;
  assign new_n37500_ = \b[11]  & ~new_n37361_;
  assign new_n37501_ = ~new_n37355_ & new_n37500_;
  assign new_n37502_ = ~new_n37363_ & ~new_n37501_;
  assign new_n37503_ = ~new_n37499_ & new_n37502_;
  assign new_n37504_ = ~new_n37363_ & ~new_n37503_;
  assign new_n37505_ = \b[12]  & ~new_n37352_;
  assign new_n37506_ = ~new_n37346_ & new_n37505_;
  assign new_n37507_ = ~new_n37354_ & ~new_n37506_;
  assign new_n37508_ = ~new_n37504_ & new_n37507_;
  assign new_n37509_ = ~new_n37354_ & ~new_n37508_;
  assign new_n37510_ = \b[13]  & ~new_n37343_;
  assign new_n37511_ = ~new_n37337_ & new_n37510_;
  assign new_n37512_ = ~new_n37345_ & ~new_n37511_;
  assign new_n37513_ = ~new_n37509_ & new_n37512_;
  assign new_n37514_ = ~new_n37345_ & ~new_n37513_;
  assign new_n37515_ = \b[14]  & ~new_n37334_;
  assign new_n37516_ = ~new_n37328_ & new_n37515_;
  assign new_n37517_ = ~new_n37336_ & ~new_n37516_;
  assign new_n37518_ = ~new_n37514_ & new_n37517_;
  assign new_n37519_ = ~new_n37336_ & ~new_n37518_;
  assign new_n37520_ = \b[15]  & ~new_n37325_;
  assign new_n37521_ = ~new_n37319_ & new_n37520_;
  assign new_n37522_ = ~new_n37327_ & ~new_n37521_;
  assign new_n37523_ = ~new_n37519_ & new_n37522_;
  assign new_n37524_ = ~new_n37327_ & ~new_n37523_;
  assign new_n37525_ = \b[16]  & ~new_n37316_;
  assign new_n37526_ = ~new_n37310_ & new_n37525_;
  assign new_n37527_ = ~new_n37318_ & ~new_n37526_;
  assign new_n37528_ = ~new_n37524_ & new_n37527_;
  assign new_n37529_ = ~new_n37318_ & ~new_n37528_;
  assign new_n37530_ = \b[17]  & ~new_n37307_;
  assign new_n37531_ = ~new_n37301_ & new_n37530_;
  assign new_n37532_ = ~new_n37309_ & ~new_n37531_;
  assign new_n37533_ = ~new_n37529_ & new_n37532_;
  assign new_n37534_ = ~new_n37309_ & ~new_n37533_;
  assign new_n37535_ = \b[18]  & ~new_n37298_;
  assign new_n37536_ = ~new_n37292_ & new_n37535_;
  assign new_n37537_ = ~new_n37300_ & ~new_n37536_;
  assign new_n37538_ = ~new_n37534_ & new_n37537_;
  assign new_n37539_ = ~new_n37300_ & ~new_n37538_;
  assign new_n37540_ = \b[19]  & ~new_n37289_;
  assign new_n37541_ = ~new_n37283_ & new_n37540_;
  assign new_n37542_ = ~new_n37291_ & ~new_n37541_;
  assign new_n37543_ = ~new_n37539_ & new_n37542_;
  assign new_n37544_ = ~new_n37291_ & ~new_n37543_;
  assign new_n37545_ = \b[20]  & ~new_n37280_;
  assign new_n37546_ = ~new_n37274_ & new_n37545_;
  assign new_n37547_ = ~new_n37282_ & ~new_n37546_;
  assign new_n37548_ = ~new_n37544_ & new_n37547_;
  assign new_n37549_ = ~new_n37282_ & ~new_n37548_;
  assign new_n37550_ = \b[21]  & ~new_n37271_;
  assign new_n37551_ = ~new_n37265_ & new_n37550_;
  assign new_n37552_ = ~new_n37273_ & ~new_n37551_;
  assign new_n37553_ = ~new_n37549_ & new_n37552_;
  assign new_n37554_ = ~new_n37273_ & ~new_n37553_;
  assign new_n37555_ = \b[22]  & ~new_n37262_;
  assign new_n37556_ = ~new_n37256_ & new_n37555_;
  assign new_n37557_ = ~new_n37264_ & ~new_n37556_;
  assign new_n37558_ = ~new_n37554_ & new_n37557_;
  assign new_n37559_ = ~new_n37264_ & ~new_n37558_;
  assign new_n37560_ = \b[23]  & ~new_n37253_;
  assign new_n37561_ = ~new_n37247_ & new_n37560_;
  assign new_n37562_ = ~new_n37255_ & ~new_n37561_;
  assign new_n37563_ = ~new_n37559_ & new_n37562_;
  assign new_n37564_ = ~new_n37255_ & ~new_n37563_;
  assign new_n37565_ = \b[24]  & ~new_n37244_;
  assign new_n37566_ = ~new_n37238_ & new_n37565_;
  assign new_n37567_ = ~new_n37246_ & ~new_n37566_;
  assign new_n37568_ = ~new_n37564_ & new_n37567_;
  assign new_n37569_ = ~new_n37246_ & ~new_n37568_;
  assign new_n37570_ = \b[25]  & ~new_n37235_;
  assign new_n37571_ = ~new_n37229_ & new_n37570_;
  assign new_n37572_ = ~new_n37237_ & ~new_n37571_;
  assign new_n37573_ = ~new_n37569_ & new_n37572_;
  assign new_n37574_ = ~new_n37237_ & ~new_n37573_;
  assign new_n37575_ = \b[26]  & ~new_n37226_;
  assign new_n37576_ = ~new_n37220_ & new_n37575_;
  assign new_n37577_ = ~new_n37228_ & ~new_n37576_;
  assign new_n37578_ = ~new_n37574_ & new_n37577_;
  assign new_n37579_ = ~new_n37228_ & ~new_n37578_;
  assign new_n37580_ = \b[27]  & ~new_n37217_;
  assign new_n37581_ = ~new_n37211_ & new_n37580_;
  assign new_n37582_ = ~new_n37219_ & ~new_n37581_;
  assign new_n37583_ = ~new_n37579_ & new_n37582_;
  assign new_n37584_ = ~new_n37219_ & ~new_n37583_;
  assign new_n37585_ = \b[28]  & ~new_n37208_;
  assign new_n37586_ = ~new_n37202_ & new_n37585_;
  assign new_n37587_ = ~new_n37210_ & ~new_n37586_;
  assign new_n37588_ = ~new_n37584_ & new_n37587_;
  assign new_n37589_ = ~new_n37210_ & ~new_n37588_;
  assign new_n37590_ = \b[29]  & ~new_n37199_;
  assign new_n37591_ = ~new_n37193_ & new_n37590_;
  assign new_n37592_ = ~new_n37201_ & ~new_n37591_;
  assign new_n37593_ = ~new_n37589_ & new_n37592_;
  assign new_n37594_ = ~new_n37201_ & ~new_n37593_;
  assign new_n37595_ = \b[30]  & ~new_n37190_;
  assign new_n37596_ = ~new_n37184_ & new_n37595_;
  assign new_n37597_ = ~new_n37192_ & ~new_n37596_;
  assign new_n37598_ = ~new_n37594_ & new_n37597_;
  assign new_n37599_ = ~new_n37192_ & ~new_n37598_;
  assign new_n37600_ = \b[31]  & ~new_n37181_;
  assign new_n37601_ = ~new_n37175_ & new_n37600_;
  assign new_n37602_ = ~new_n37183_ & ~new_n37601_;
  assign new_n37603_ = ~new_n37599_ & new_n37602_;
  assign new_n37604_ = ~new_n37183_ & ~new_n37603_;
  assign new_n37605_ = \b[32]  & ~new_n37172_;
  assign new_n37606_ = ~new_n37166_ & new_n37605_;
  assign new_n37607_ = ~new_n37174_ & ~new_n37606_;
  assign new_n37608_ = ~new_n37604_ & new_n37607_;
  assign new_n37609_ = ~new_n37174_ & ~new_n37608_;
  assign new_n37610_ = \b[33]  & ~new_n37163_;
  assign new_n37611_ = ~new_n37157_ & new_n37610_;
  assign new_n37612_ = ~new_n37165_ & ~new_n37611_;
  assign new_n37613_ = ~new_n37609_ & new_n37612_;
  assign new_n37614_ = ~new_n37165_ & ~new_n37613_;
  assign new_n37615_ = \b[34]  & ~new_n37154_;
  assign new_n37616_ = ~new_n37148_ & new_n37615_;
  assign new_n37617_ = ~new_n37156_ & ~new_n37616_;
  assign new_n37618_ = ~new_n37614_ & new_n37617_;
  assign new_n37619_ = ~new_n37156_ & ~new_n37618_;
  assign new_n37620_ = ~new_n36690_ & ~new_n37147_;
  assign new_n37621_ = ~new_n36692_ & new_n37144_;
  assign new_n37622_ = ~new_n37140_ & new_n37621_;
  assign new_n37623_ = ~new_n37141_ & ~new_n37144_;
  assign new_n37624_ = ~new_n37622_ & ~new_n37623_;
  assign new_n37625_ = new_n37147_ & ~new_n37624_;
  assign new_n37626_ = ~new_n37620_ & ~new_n37625_;
  assign new_n37627_ = ~\b[35]  & ~new_n37626_;
  assign new_n37628_ = \b[35]  & ~new_n37620_;
  assign new_n37629_ = ~new_n37625_ & new_n37628_;
  assign new_n37630_ = new_n512_ & ~new_n37629_;
  assign new_n37631_ = ~new_n37627_ & new_n37630_;
  assign new_n37632_ = ~new_n37619_ & new_n37631_;
  assign new_n37633_ = new_n9004_ & ~new_n37626_;
  assign new_n37634_ = ~new_n37632_ & ~new_n37633_;
  assign new_n37635_ = ~new_n37165_ & new_n37617_;
  assign new_n37636_ = ~new_n37613_ & new_n37635_;
  assign new_n37637_ = ~new_n37614_ & ~new_n37617_;
  assign new_n37638_ = ~new_n37636_ & ~new_n37637_;
  assign new_n37639_ = ~new_n37634_ & ~new_n37638_;
  assign new_n37640_ = ~new_n37155_ & ~new_n37633_;
  assign new_n37641_ = ~new_n37632_ & new_n37640_;
  assign new_n37642_ = ~new_n37639_ & ~new_n37641_;
  assign new_n37643_ = ~new_n37156_ & ~new_n37629_;
  assign new_n37644_ = ~new_n37627_ & new_n37643_;
  assign new_n37645_ = ~new_n37618_ & new_n37644_;
  assign new_n37646_ = ~new_n37627_ & ~new_n37629_;
  assign new_n37647_ = ~new_n37619_ & ~new_n37646_;
  assign new_n37648_ = ~new_n37645_ & ~new_n37647_;
  assign new_n37649_ = ~new_n37634_ & ~new_n37648_;
  assign new_n37650_ = ~new_n37626_ & ~new_n37633_;
  assign new_n37651_ = ~new_n37632_ & new_n37650_;
  assign new_n37652_ = ~new_n37649_ & ~new_n37651_;
  assign new_n37653_ = ~\b[36]  & ~new_n37652_;
  assign new_n37654_ = ~\b[35]  & ~new_n37642_;
  assign new_n37655_ = ~new_n37174_ & new_n37612_;
  assign new_n37656_ = ~new_n37608_ & new_n37655_;
  assign new_n37657_ = ~new_n37609_ & ~new_n37612_;
  assign new_n37658_ = ~new_n37656_ & ~new_n37657_;
  assign new_n37659_ = ~new_n37634_ & ~new_n37658_;
  assign new_n37660_ = ~new_n37164_ & ~new_n37633_;
  assign new_n37661_ = ~new_n37632_ & new_n37660_;
  assign new_n37662_ = ~new_n37659_ & ~new_n37661_;
  assign new_n37663_ = ~\b[34]  & ~new_n37662_;
  assign new_n37664_ = ~new_n37183_ & new_n37607_;
  assign new_n37665_ = ~new_n37603_ & new_n37664_;
  assign new_n37666_ = ~new_n37604_ & ~new_n37607_;
  assign new_n37667_ = ~new_n37665_ & ~new_n37666_;
  assign new_n37668_ = ~new_n37634_ & ~new_n37667_;
  assign new_n37669_ = ~new_n37173_ & ~new_n37633_;
  assign new_n37670_ = ~new_n37632_ & new_n37669_;
  assign new_n37671_ = ~new_n37668_ & ~new_n37670_;
  assign new_n37672_ = ~\b[33]  & ~new_n37671_;
  assign new_n37673_ = ~new_n37192_ & new_n37602_;
  assign new_n37674_ = ~new_n37598_ & new_n37673_;
  assign new_n37675_ = ~new_n37599_ & ~new_n37602_;
  assign new_n37676_ = ~new_n37674_ & ~new_n37675_;
  assign new_n37677_ = ~new_n37634_ & ~new_n37676_;
  assign new_n37678_ = ~new_n37182_ & ~new_n37633_;
  assign new_n37679_ = ~new_n37632_ & new_n37678_;
  assign new_n37680_ = ~new_n37677_ & ~new_n37679_;
  assign new_n37681_ = ~\b[32]  & ~new_n37680_;
  assign new_n37682_ = ~new_n37201_ & new_n37597_;
  assign new_n37683_ = ~new_n37593_ & new_n37682_;
  assign new_n37684_ = ~new_n37594_ & ~new_n37597_;
  assign new_n37685_ = ~new_n37683_ & ~new_n37684_;
  assign new_n37686_ = ~new_n37634_ & ~new_n37685_;
  assign new_n37687_ = ~new_n37191_ & ~new_n37633_;
  assign new_n37688_ = ~new_n37632_ & new_n37687_;
  assign new_n37689_ = ~new_n37686_ & ~new_n37688_;
  assign new_n37690_ = ~\b[31]  & ~new_n37689_;
  assign new_n37691_ = ~new_n37210_ & new_n37592_;
  assign new_n37692_ = ~new_n37588_ & new_n37691_;
  assign new_n37693_ = ~new_n37589_ & ~new_n37592_;
  assign new_n37694_ = ~new_n37692_ & ~new_n37693_;
  assign new_n37695_ = ~new_n37634_ & ~new_n37694_;
  assign new_n37696_ = ~new_n37200_ & ~new_n37633_;
  assign new_n37697_ = ~new_n37632_ & new_n37696_;
  assign new_n37698_ = ~new_n37695_ & ~new_n37697_;
  assign new_n37699_ = ~\b[30]  & ~new_n37698_;
  assign new_n37700_ = ~new_n37219_ & new_n37587_;
  assign new_n37701_ = ~new_n37583_ & new_n37700_;
  assign new_n37702_ = ~new_n37584_ & ~new_n37587_;
  assign new_n37703_ = ~new_n37701_ & ~new_n37702_;
  assign new_n37704_ = ~new_n37634_ & ~new_n37703_;
  assign new_n37705_ = ~new_n37209_ & ~new_n37633_;
  assign new_n37706_ = ~new_n37632_ & new_n37705_;
  assign new_n37707_ = ~new_n37704_ & ~new_n37706_;
  assign new_n37708_ = ~\b[29]  & ~new_n37707_;
  assign new_n37709_ = ~new_n37228_ & new_n37582_;
  assign new_n37710_ = ~new_n37578_ & new_n37709_;
  assign new_n37711_ = ~new_n37579_ & ~new_n37582_;
  assign new_n37712_ = ~new_n37710_ & ~new_n37711_;
  assign new_n37713_ = ~new_n37634_ & ~new_n37712_;
  assign new_n37714_ = ~new_n37218_ & ~new_n37633_;
  assign new_n37715_ = ~new_n37632_ & new_n37714_;
  assign new_n37716_ = ~new_n37713_ & ~new_n37715_;
  assign new_n37717_ = ~\b[28]  & ~new_n37716_;
  assign new_n37718_ = ~new_n37237_ & new_n37577_;
  assign new_n37719_ = ~new_n37573_ & new_n37718_;
  assign new_n37720_ = ~new_n37574_ & ~new_n37577_;
  assign new_n37721_ = ~new_n37719_ & ~new_n37720_;
  assign new_n37722_ = ~new_n37634_ & ~new_n37721_;
  assign new_n37723_ = ~new_n37227_ & ~new_n37633_;
  assign new_n37724_ = ~new_n37632_ & new_n37723_;
  assign new_n37725_ = ~new_n37722_ & ~new_n37724_;
  assign new_n37726_ = ~\b[27]  & ~new_n37725_;
  assign new_n37727_ = ~new_n37246_ & new_n37572_;
  assign new_n37728_ = ~new_n37568_ & new_n37727_;
  assign new_n37729_ = ~new_n37569_ & ~new_n37572_;
  assign new_n37730_ = ~new_n37728_ & ~new_n37729_;
  assign new_n37731_ = ~new_n37634_ & ~new_n37730_;
  assign new_n37732_ = ~new_n37236_ & ~new_n37633_;
  assign new_n37733_ = ~new_n37632_ & new_n37732_;
  assign new_n37734_ = ~new_n37731_ & ~new_n37733_;
  assign new_n37735_ = ~\b[26]  & ~new_n37734_;
  assign new_n37736_ = ~new_n37255_ & new_n37567_;
  assign new_n37737_ = ~new_n37563_ & new_n37736_;
  assign new_n37738_ = ~new_n37564_ & ~new_n37567_;
  assign new_n37739_ = ~new_n37737_ & ~new_n37738_;
  assign new_n37740_ = ~new_n37634_ & ~new_n37739_;
  assign new_n37741_ = ~new_n37245_ & ~new_n37633_;
  assign new_n37742_ = ~new_n37632_ & new_n37741_;
  assign new_n37743_ = ~new_n37740_ & ~new_n37742_;
  assign new_n37744_ = ~\b[25]  & ~new_n37743_;
  assign new_n37745_ = ~new_n37264_ & new_n37562_;
  assign new_n37746_ = ~new_n37558_ & new_n37745_;
  assign new_n37747_ = ~new_n37559_ & ~new_n37562_;
  assign new_n37748_ = ~new_n37746_ & ~new_n37747_;
  assign new_n37749_ = ~new_n37634_ & ~new_n37748_;
  assign new_n37750_ = ~new_n37254_ & ~new_n37633_;
  assign new_n37751_ = ~new_n37632_ & new_n37750_;
  assign new_n37752_ = ~new_n37749_ & ~new_n37751_;
  assign new_n37753_ = ~\b[24]  & ~new_n37752_;
  assign new_n37754_ = ~new_n37273_ & new_n37557_;
  assign new_n37755_ = ~new_n37553_ & new_n37754_;
  assign new_n37756_ = ~new_n37554_ & ~new_n37557_;
  assign new_n37757_ = ~new_n37755_ & ~new_n37756_;
  assign new_n37758_ = ~new_n37634_ & ~new_n37757_;
  assign new_n37759_ = ~new_n37263_ & ~new_n37633_;
  assign new_n37760_ = ~new_n37632_ & new_n37759_;
  assign new_n37761_ = ~new_n37758_ & ~new_n37760_;
  assign new_n37762_ = ~\b[23]  & ~new_n37761_;
  assign new_n37763_ = ~new_n37282_ & new_n37552_;
  assign new_n37764_ = ~new_n37548_ & new_n37763_;
  assign new_n37765_ = ~new_n37549_ & ~new_n37552_;
  assign new_n37766_ = ~new_n37764_ & ~new_n37765_;
  assign new_n37767_ = ~new_n37634_ & ~new_n37766_;
  assign new_n37768_ = ~new_n37272_ & ~new_n37633_;
  assign new_n37769_ = ~new_n37632_ & new_n37768_;
  assign new_n37770_ = ~new_n37767_ & ~new_n37769_;
  assign new_n37771_ = ~\b[22]  & ~new_n37770_;
  assign new_n37772_ = ~new_n37291_ & new_n37547_;
  assign new_n37773_ = ~new_n37543_ & new_n37772_;
  assign new_n37774_ = ~new_n37544_ & ~new_n37547_;
  assign new_n37775_ = ~new_n37773_ & ~new_n37774_;
  assign new_n37776_ = ~new_n37634_ & ~new_n37775_;
  assign new_n37777_ = ~new_n37281_ & ~new_n37633_;
  assign new_n37778_ = ~new_n37632_ & new_n37777_;
  assign new_n37779_ = ~new_n37776_ & ~new_n37778_;
  assign new_n37780_ = ~\b[21]  & ~new_n37779_;
  assign new_n37781_ = ~new_n37300_ & new_n37542_;
  assign new_n37782_ = ~new_n37538_ & new_n37781_;
  assign new_n37783_ = ~new_n37539_ & ~new_n37542_;
  assign new_n37784_ = ~new_n37782_ & ~new_n37783_;
  assign new_n37785_ = ~new_n37634_ & ~new_n37784_;
  assign new_n37786_ = ~new_n37290_ & ~new_n37633_;
  assign new_n37787_ = ~new_n37632_ & new_n37786_;
  assign new_n37788_ = ~new_n37785_ & ~new_n37787_;
  assign new_n37789_ = ~\b[20]  & ~new_n37788_;
  assign new_n37790_ = ~new_n37309_ & new_n37537_;
  assign new_n37791_ = ~new_n37533_ & new_n37790_;
  assign new_n37792_ = ~new_n37534_ & ~new_n37537_;
  assign new_n37793_ = ~new_n37791_ & ~new_n37792_;
  assign new_n37794_ = ~new_n37634_ & ~new_n37793_;
  assign new_n37795_ = ~new_n37299_ & ~new_n37633_;
  assign new_n37796_ = ~new_n37632_ & new_n37795_;
  assign new_n37797_ = ~new_n37794_ & ~new_n37796_;
  assign new_n37798_ = ~\b[19]  & ~new_n37797_;
  assign new_n37799_ = ~new_n37318_ & new_n37532_;
  assign new_n37800_ = ~new_n37528_ & new_n37799_;
  assign new_n37801_ = ~new_n37529_ & ~new_n37532_;
  assign new_n37802_ = ~new_n37800_ & ~new_n37801_;
  assign new_n37803_ = ~new_n37634_ & ~new_n37802_;
  assign new_n37804_ = ~new_n37308_ & ~new_n37633_;
  assign new_n37805_ = ~new_n37632_ & new_n37804_;
  assign new_n37806_ = ~new_n37803_ & ~new_n37805_;
  assign new_n37807_ = ~\b[18]  & ~new_n37806_;
  assign new_n37808_ = ~new_n37327_ & new_n37527_;
  assign new_n37809_ = ~new_n37523_ & new_n37808_;
  assign new_n37810_ = ~new_n37524_ & ~new_n37527_;
  assign new_n37811_ = ~new_n37809_ & ~new_n37810_;
  assign new_n37812_ = ~new_n37634_ & ~new_n37811_;
  assign new_n37813_ = ~new_n37317_ & ~new_n37633_;
  assign new_n37814_ = ~new_n37632_ & new_n37813_;
  assign new_n37815_ = ~new_n37812_ & ~new_n37814_;
  assign new_n37816_ = ~\b[17]  & ~new_n37815_;
  assign new_n37817_ = ~new_n37336_ & new_n37522_;
  assign new_n37818_ = ~new_n37518_ & new_n37817_;
  assign new_n37819_ = ~new_n37519_ & ~new_n37522_;
  assign new_n37820_ = ~new_n37818_ & ~new_n37819_;
  assign new_n37821_ = ~new_n37634_ & ~new_n37820_;
  assign new_n37822_ = ~new_n37326_ & ~new_n37633_;
  assign new_n37823_ = ~new_n37632_ & new_n37822_;
  assign new_n37824_ = ~new_n37821_ & ~new_n37823_;
  assign new_n37825_ = ~\b[16]  & ~new_n37824_;
  assign new_n37826_ = ~new_n37345_ & new_n37517_;
  assign new_n37827_ = ~new_n37513_ & new_n37826_;
  assign new_n37828_ = ~new_n37514_ & ~new_n37517_;
  assign new_n37829_ = ~new_n37827_ & ~new_n37828_;
  assign new_n37830_ = ~new_n37634_ & ~new_n37829_;
  assign new_n37831_ = ~new_n37335_ & ~new_n37633_;
  assign new_n37832_ = ~new_n37632_ & new_n37831_;
  assign new_n37833_ = ~new_n37830_ & ~new_n37832_;
  assign new_n37834_ = ~\b[15]  & ~new_n37833_;
  assign new_n37835_ = ~new_n37354_ & new_n37512_;
  assign new_n37836_ = ~new_n37508_ & new_n37835_;
  assign new_n37837_ = ~new_n37509_ & ~new_n37512_;
  assign new_n37838_ = ~new_n37836_ & ~new_n37837_;
  assign new_n37839_ = ~new_n37634_ & ~new_n37838_;
  assign new_n37840_ = ~new_n37344_ & ~new_n37633_;
  assign new_n37841_ = ~new_n37632_ & new_n37840_;
  assign new_n37842_ = ~new_n37839_ & ~new_n37841_;
  assign new_n37843_ = ~\b[14]  & ~new_n37842_;
  assign new_n37844_ = ~new_n37363_ & new_n37507_;
  assign new_n37845_ = ~new_n37503_ & new_n37844_;
  assign new_n37846_ = ~new_n37504_ & ~new_n37507_;
  assign new_n37847_ = ~new_n37845_ & ~new_n37846_;
  assign new_n37848_ = ~new_n37634_ & ~new_n37847_;
  assign new_n37849_ = ~new_n37353_ & ~new_n37633_;
  assign new_n37850_ = ~new_n37632_ & new_n37849_;
  assign new_n37851_ = ~new_n37848_ & ~new_n37850_;
  assign new_n37852_ = ~\b[13]  & ~new_n37851_;
  assign new_n37853_ = ~new_n37372_ & new_n37502_;
  assign new_n37854_ = ~new_n37498_ & new_n37853_;
  assign new_n37855_ = ~new_n37499_ & ~new_n37502_;
  assign new_n37856_ = ~new_n37854_ & ~new_n37855_;
  assign new_n37857_ = ~new_n37634_ & ~new_n37856_;
  assign new_n37858_ = ~new_n37362_ & ~new_n37633_;
  assign new_n37859_ = ~new_n37632_ & new_n37858_;
  assign new_n37860_ = ~new_n37857_ & ~new_n37859_;
  assign new_n37861_ = ~\b[12]  & ~new_n37860_;
  assign new_n37862_ = ~new_n37381_ & new_n37497_;
  assign new_n37863_ = ~new_n37493_ & new_n37862_;
  assign new_n37864_ = ~new_n37494_ & ~new_n37497_;
  assign new_n37865_ = ~new_n37863_ & ~new_n37864_;
  assign new_n37866_ = ~new_n37634_ & ~new_n37865_;
  assign new_n37867_ = ~new_n37371_ & ~new_n37633_;
  assign new_n37868_ = ~new_n37632_ & new_n37867_;
  assign new_n37869_ = ~new_n37866_ & ~new_n37868_;
  assign new_n37870_ = ~\b[11]  & ~new_n37869_;
  assign new_n37871_ = ~new_n37390_ & new_n37492_;
  assign new_n37872_ = ~new_n37488_ & new_n37871_;
  assign new_n37873_ = ~new_n37489_ & ~new_n37492_;
  assign new_n37874_ = ~new_n37872_ & ~new_n37873_;
  assign new_n37875_ = ~new_n37634_ & ~new_n37874_;
  assign new_n37876_ = ~new_n37380_ & ~new_n37633_;
  assign new_n37877_ = ~new_n37632_ & new_n37876_;
  assign new_n37878_ = ~new_n37875_ & ~new_n37877_;
  assign new_n37879_ = ~\b[10]  & ~new_n37878_;
  assign new_n37880_ = ~new_n37399_ & new_n37487_;
  assign new_n37881_ = ~new_n37483_ & new_n37880_;
  assign new_n37882_ = ~new_n37484_ & ~new_n37487_;
  assign new_n37883_ = ~new_n37881_ & ~new_n37882_;
  assign new_n37884_ = ~new_n37634_ & ~new_n37883_;
  assign new_n37885_ = ~new_n37389_ & ~new_n37633_;
  assign new_n37886_ = ~new_n37632_ & new_n37885_;
  assign new_n37887_ = ~new_n37884_ & ~new_n37886_;
  assign new_n37888_ = ~\b[9]  & ~new_n37887_;
  assign new_n37889_ = ~new_n37408_ & new_n37482_;
  assign new_n37890_ = ~new_n37478_ & new_n37889_;
  assign new_n37891_ = ~new_n37479_ & ~new_n37482_;
  assign new_n37892_ = ~new_n37890_ & ~new_n37891_;
  assign new_n37893_ = ~new_n37634_ & ~new_n37892_;
  assign new_n37894_ = ~new_n37398_ & ~new_n37633_;
  assign new_n37895_ = ~new_n37632_ & new_n37894_;
  assign new_n37896_ = ~new_n37893_ & ~new_n37895_;
  assign new_n37897_ = ~\b[8]  & ~new_n37896_;
  assign new_n37898_ = ~new_n37417_ & new_n37477_;
  assign new_n37899_ = ~new_n37473_ & new_n37898_;
  assign new_n37900_ = ~new_n37474_ & ~new_n37477_;
  assign new_n37901_ = ~new_n37899_ & ~new_n37900_;
  assign new_n37902_ = ~new_n37634_ & ~new_n37901_;
  assign new_n37903_ = ~new_n37407_ & ~new_n37633_;
  assign new_n37904_ = ~new_n37632_ & new_n37903_;
  assign new_n37905_ = ~new_n37902_ & ~new_n37904_;
  assign new_n37906_ = ~\b[7]  & ~new_n37905_;
  assign new_n37907_ = ~new_n37426_ & new_n37472_;
  assign new_n37908_ = ~new_n37468_ & new_n37907_;
  assign new_n37909_ = ~new_n37469_ & ~new_n37472_;
  assign new_n37910_ = ~new_n37908_ & ~new_n37909_;
  assign new_n37911_ = ~new_n37634_ & ~new_n37910_;
  assign new_n37912_ = ~new_n37416_ & ~new_n37633_;
  assign new_n37913_ = ~new_n37632_ & new_n37912_;
  assign new_n37914_ = ~new_n37911_ & ~new_n37913_;
  assign new_n37915_ = ~\b[6]  & ~new_n37914_;
  assign new_n37916_ = ~new_n37435_ & new_n37467_;
  assign new_n37917_ = ~new_n37463_ & new_n37916_;
  assign new_n37918_ = ~new_n37464_ & ~new_n37467_;
  assign new_n37919_ = ~new_n37917_ & ~new_n37918_;
  assign new_n37920_ = ~new_n37634_ & ~new_n37919_;
  assign new_n37921_ = ~new_n37425_ & ~new_n37633_;
  assign new_n37922_ = ~new_n37632_ & new_n37921_;
  assign new_n37923_ = ~new_n37920_ & ~new_n37922_;
  assign new_n37924_ = ~\b[5]  & ~new_n37923_;
  assign new_n37925_ = ~new_n37443_ & new_n37462_;
  assign new_n37926_ = ~new_n37458_ & new_n37925_;
  assign new_n37927_ = ~new_n37459_ & ~new_n37462_;
  assign new_n37928_ = ~new_n37926_ & ~new_n37927_;
  assign new_n37929_ = ~new_n37634_ & ~new_n37928_;
  assign new_n37930_ = ~new_n37434_ & ~new_n37633_;
  assign new_n37931_ = ~new_n37632_ & new_n37930_;
  assign new_n37932_ = ~new_n37929_ & ~new_n37931_;
  assign new_n37933_ = ~\b[4]  & ~new_n37932_;
  assign new_n37934_ = ~new_n37453_ & new_n37457_;
  assign new_n37935_ = ~new_n37452_ & new_n37934_;
  assign new_n37936_ = ~new_n37454_ & ~new_n37457_;
  assign new_n37937_ = ~new_n37935_ & ~new_n37936_;
  assign new_n37938_ = ~new_n37634_ & ~new_n37937_;
  assign new_n37939_ = ~new_n37442_ & ~new_n37633_;
  assign new_n37940_ = ~new_n37632_ & new_n37939_;
  assign new_n37941_ = ~new_n37938_ & ~new_n37940_;
  assign new_n37942_ = ~\b[3]  & ~new_n37941_;
  assign new_n37943_ = new_n9318_ & ~new_n37450_;
  assign new_n37944_ = ~new_n37448_ & new_n37943_;
  assign new_n37945_ = ~new_n37452_ & ~new_n37944_;
  assign new_n37946_ = ~new_n37634_ & new_n37945_;
  assign new_n37947_ = ~new_n37447_ & ~new_n37633_;
  assign new_n37948_ = ~new_n37632_ & new_n37947_;
  assign new_n37949_ = ~new_n37946_ & ~new_n37948_;
  assign new_n37950_ = ~\b[2]  & ~new_n37949_;
  assign new_n37951_ = \b[0]  & ~new_n37634_;
  assign new_n37952_ = \a[28]  & ~new_n37951_;
  assign new_n37953_ = new_n9318_ & ~new_n37634_;
  assign new_n37954_ = ~new_n37952_ & ~new_n37953_;
  assign new_n37955_ = \b[1]  & ~new_n37954_;
  assign new_n37956_ = ~\b[1]  & ~new_n37953_;
  assign new_n37957_ = ~new_n37952_ & new_n37956_;
  assign new_n37958_ = ~new_n37955_ & ~new_n37957_;
  assign new_n37959_ = ~new_n9826_ & ~new_n37958_;
  assign new_n37960_ = ~\b[1]  & ~new_n37954_;
  assign new_n37961_ = ~new_n37959_ & ~new_n37960_;
  assign new_n37962_ = \b[2]  & ~new_n37948_;
  assign new_n37963_ = ~new_n37946_ & new_n37962_;
  assign new_n37964_ = ~new_n37950_ & ~new_n37963_;
  assign new_n37965_ = ~new_n37961_ & new_n37964_;
  assign new_n37966_ = ~new_n37950_ & ~new_n37965_;
  assign new_n37967_ = \b[3]  & ~new_n37940_;
  assign new_n37968_ = ~new_n37938_ & new_n37967_;
  assign new_n37969_ = ~new_n37942_ & ~new_n37968_;
  assign new_n37970_ = ~new_n37966_ & new_n37969_;
  assign new_n37971_ = ~new_n37942_ & ~new_n37970_;
  assign new_n37972_ = \b[4]  & ~new_n37931_;
  assign new_n37973_ = ~new_n37929_ & new_n37972_;
  assign new_n37974_ = ~new_n37933_ & ~new_n37973_;
  assign new_n37975_ = ~new_n37971_ & new_n37974_;
  assign new_n37976_ = ~new_n37933_ & ~new_n37975_;
  assign new_n37977_ = \b[5]  & ~new_n37922_;
  assign new_n37978_ = ~new_n37920_ & new_n37977_;
  assign new_n37979_ = ~new_n37924_ & ~new_n37978_;
  assign new_n37980_ = ~new_n37976_ & new_n37979_;
  assign new_n37981_ = ~new_n37924_ & ~new_n37980_;
  assign new_n37982_ = \b[6]  & ~new_n37913_;
  assign new_n37983_ = ~new_n37911_ & new_n37982_;
  assign new_n37984_ = ~new_n37915_ & ~new_n37983_;
  assign new_n37985_ = ~new_n37981_ & new_n37984_;
  assign new_n37986_ = ~new_n37915_ & ~new_n37985_;
  assign new_n37987_ = \b[7]  & ~new_n37904_;
  assign new_n37988_ = ~new_n37902_ & new_n37987_;
  assign new_n37989_ = ~new_n37906_ & ~new_n37988_;
  assign new_n37990_ = ~new_n37986_ & new_n37989_;
  assign new_n37991_ = ~new_n37906_ & ~new_n37990_;
  assign new_n37992_ = \b[8]  & ~new_n37895_;
  assign new_n37993_ = ~new_n37893_ & new_n37992_;
  assign new_n37994_ = ~new_n37897_ & ~new_n37993_;
  assign new_n37995_ = ~new_n37991_ & new_n37994_;
  assign new_n37996_ = ~new_n37897_ & ~new_n37995_;
  assign new_n37997_ = \b[9]  & ~new_n37886_;
  assign new_n37998_ = ~new_n37884_ & new_n37997_;
  assign new_n37999_ = ~new_n37888_ & ~new_n37998_;
  assign new_n38000_ = ~new_n37996_ & new_n37999_;
  assign new_n38001_ = ~new_n37888_ & ~new_n38000_;
  assign new_n38002_ = \b[10]  & ~new_n37877_;
  assign new_n38003_ = ~new_n37875_ & new_n38002_;
  assign new_n38004_ = ~new_n37879_ & ~new_n38003_;
  assign new_n38005_ = ~new_n38001_ & new_n38004_;
  assign new_n38006_ = ~new_n37879_ & ~new_n38005_;
  assign new_n38007_ = \b[11]  & ~new_n37868_;
  assign new_n38008_ = ~new_n37866_ & new_n38007_;
  assign new_n38009_ = ~new_n37870_ & ~new_n38008_;
  assign new_n38010_ = ~new_n38006_ & new_n38009_;
  assign new_n38011_ = ~new_n37870_ & ~new_n38010_;
  assign new_n38012_ = \b[12]  & ~new_n37859_;
  assign new_n38013_ = ~new_n37857_ & new_n38012_;
  assign new_n38014_ = ~new_n37861_ & ~new_n38013_;
  assign new_n38015_ = ~new_n38011_ & new_n38014_;
  assign new_n38016_ = ~new_n37861_ & ~new_n38015_;
  assign new_n38017_ = \b[13]  & ~new_n37850_;
  assign new_n38018_ = ~new_n37848_ & new_n38017_;
  assign new_n38019_ = ~new_n37852_ & ~new_n38018_;
  assign new_n38020_ = ~new_n38016_ & new_n38019_;
  assign new_n38021_ = ~new_n37852_ & ~new_n38020_;
  assign new_n38022_ = \b[14]  & ~new_n37841_;
  assign new_n38023_ = ~new_n37839_ & new_n38022_;
  assign new_n38024_ = ~new_n37843_ & ~new_n38023_;
  assign new_n38025_ = ~new_n38021_ & new_n38024_;
  assign new_n38026_ = ~new_n37843_ & ~new_n38025_;
  assign new_n38027_ = \b[15]  & ~new_n37832_;
  assign new_n38028_ = ~new_n37830_ & new_n38027_;
  assign new_n38029_ = ~new_n37834_ & ~new_n38028_;
  assign new_n38030_ = ~new_n38026_ & new_n38029_;
  assign new_n38031_ = ~new_n37834_ & ~new_n38030_;
  assign new_n38032_ = \b[16]  & ~new_n37823_;
  assign new_n38033_ = ~new_n37821_ & new_n38032_;
  assign new_n38034_ = ~new_n37825_ & ~new_n38033_;
  assign new_n38035_ = ~new_n38031_ & new_n38034_;
  assign new_n38036_ = ~new_n37825_ & ~new_n38035_;
  assign new_n38037_ = \b[17]  & ~new_n37814_;
  assign new_n38038_ = ~new_n37812_ & new_n38037_;
  assign new_n38039_ = ~new_n37816_ & ~new_n38038_;
  assign new_n38040_ = ~new_n38036_ & new_n38039_;
  assign new_n38041_ = ~new_n37816_ & ~new_n38040_;
  assign new_n38042_ = \b[18]  & ~new_n37805_;
  assign new_n38043_ = ~new_n37803_ & new_n38042_;
  assign new_n38044_ = ~new_n37807_ & ~new_n38043_;
  assign new_n38045_ = ~new_n38041_ & new_n38044_;
  assign new_n38046_ = ~new_n37807_ & ~new_n38045_;
  assign new_n38047_ = \b[19]  & ~new_n37796_;
  assign new_n38048_ = ~new_n37794_ & new_n38047_;
  assign new_n38049_ = ~new_n37798_ & ~new_n38048_;
  assign new_n38050_ = ~new_n38046_ & new_n38049_;
  assign new_n38051_ = ~new_n37798_ & ~new_n38050_;
  assign new_n38052_ = \b[20]  & ~new_n37787_;
  assign new_n38053_ = ~new_n37785_ & new_n38052_;
  assign new_n38054_ = ~new_n37789_ & ~new_n38053_;
  assign new_n38055_ = ~new_n38051_ & new_n38054_;
  assign new_n38056_ = ~new_n37789_ & ~new_n38055_;
  assign new_n38057_ = \b[21]  & ~new_n37778_;
  assign new_n38058_ = ~new_n37776_ & new_n38057_;
  assign new_n38059_ = ~new_n37780_ & ~new_n38058_;
  assign new_n38060_ = ~new_n38056_ & new_n38059_;
  assign new_n38061_ = ~new_n37780_ & ~new_n38060_;
  assign new_n38062_ = \b[22]  & ~new_n37769_;
  assign new_n38063_ = ~new_n37767_ & new_n38062_;
  assign new_n38064_ = ~new_n37771_ & ~new_n38063_;
  assign new_n38065_ = ~new_n38061_ & new_n38064_;
  assign new_n38066_ = ~new_n37771_ & ~new_n38065_;
  assign new_n38067_ = \b[23]  & ~new_n37760_;
  assign new_n38068_ = ~new_n37758_ & new_n38067_;
  assign new_n38069_ = ~new_n37762_ & ~new_n38068_;
  assign new_n38070_ = ~new_n38066_ & new_n38069_;
  assign new_n38071_ = ~new_n37762_ & ~new_n38070_;
  assign new_n38072_ = \b[24]  & ~new_n37751_;
  assign new_n38073_ = ~new_n37749_ & new_n38072_;
  assign new_n38074_ = ~new_n37753_ & ~new_n38073_;
  assign new_n38075_ = ~new_n38071_ & new_n38074_;
  assign new_n38076_ = ~new_n37753_ & ~new_n38075_;
  assign new_n38077_ = \b[25]  & ~new_n37742_;
  assign new_n38078_ = ~new_n37740_ & new_n38077_;
  assign new_n38079_ = ~new_n37744_ & ~new_n38078_;
  assign new_n38080_ = ~new_n38076_ & new_n38079_;
  assign new_n38081_ = ~new_n37744_ & ~new_n38080_;
  assign new_n38082_ = \b[26]  & ~new_n37733_;
  assign new_n38083_ = ~new_n37731_ & new_n38082_;
  assign new_n38084_ = ~new_n37735_ & ~new_n38083_;
  assign new_n38085_ = ~new_n38081_ & new_n38084_;
  assign new_n38086_ = ~new_n37735_ & ~new_n38085_;
  assign new_n38087_ = \b[27]  & ~new_n37724_;
  assign new_n38088_ = ~new_n37722_ & new_n38087_;
  assign new_n38089_ = ~new_n37726_ & ~new_n38088_;
  assign new_n38090_ = ~new_n38086_ & new_n38089_;
  assign new_n38091_ = ~new_n37726_ & ~new_n38090_;
  assign new_n38092_ = \b[28]  & ~new_n37715_;
  assign new_n38093_ = ~new_n37713_ & new_n38092_;
  assign new_n38094_ = ~new_n37717_ & ~new_n38093_;
  assign new_n38095_ = ~new_n38091_ & new_n38094_;
  assign new_n38096_ = ~new_n37717_ & ~new_n38095_;
  assign new_n38097_ = \b[29]  & ~new_n37706_;
  assign new_n38098_ = ~new_n37704_ & new_n38097_;
  assign new_n38099_ = ~new_n37708_ & ~new_n38098_;
  assign new_n38100_ = ~new_n38096_ & new_n38099_;
  assign new_n38101_ = ~new_n37708_ & ~new_n38100_;
  assign new_n38102_ = \b[30]  & ~new_n37697_;
  assign new_n38103_ = ~new_n37695_ & new_n38102_;
  assign new_n38104_ = ~new_n37699_ & ~new_n38103_;
  assign new_n38105_ = ~new_n38101_ & new_n38104_;
  assign new_n38106_ = ~new_n37699_ & ~new_n38105_;
  assign new_n38107_ = \b[31]  & ~new_n37688_;
  assign new_n38108_ = ~new_n37686_ & new_n38107_;
  assign new_n38109_ = ~new_n37690_ & ~new_n38108_;
  assign new_n38110_ = ~new_n38106_ & new_n38109_;
  assign new_n38111_ = ~new_n37690_ & ~new_n38110_;
  assign new_n38112_ = \b[32]  & ~new_n37679_;
  assign new_n38113_ = ~new_n37677_ & new_n38112_;
  assign new_n38114_ = ~new_n37681_ & ~new_n38113_;
  assign new_n38115_ = ~new_n38111_ & new_n38114_;
  assign new_n38116_ = ~new_n37681_ & ~new_n38115_;
  assign new_n38117_ = \b[33]  & ~new_n37670_;
  assign new_n38118_ = ~new_n37668_ & new_n38117_;
  assign new_n38119_ = ~new_n37672_ & ~new_n38118_;
  assign new_n38120_ = ~new_n38116_ & new_n38119_;
  assign new_n38121_ = ~new_n37672_ & ~new_n38120_;
  assign new_n38122_ = \b[34]  & ~new_n37661_;
  assign new_n38123_ = ~new_n37659_ & new_n38122_;
  assign new_n38124_ = ~new_n37663_ & ~new_n38123_;
  assign new_n38125_ = ~new_n38121_ & new_n38124_;
  assign new_n38126_ = ~new_n37663_ & ~new_n38125_;
  assign new_n38127_ = \b[35]  & ~new_n37641_;
  assign new_n38128_ = ~new_n37639_ & new_n38127_;
  assign new_n38129_ = ~new_n37654_ & ~new_n38128_;
  assign new_n38130_ = ~new_n38126_ & new_n38129_;
  assign new_n38131_ = ~new_n37654_ & ~new_n38130_;
  assign new_n38132_ = \b[36]  & ~new_n37651_;
  assign new_n38133_ = ~new_n37649_ & new_n38132_;
  assign new_n38134_ = ~new_n37653_ & ~new_n38133_;
  assign new_n38135_ = ~new_n38131_ & new_n38134_;
  assign new_n38136_ = ~new_n37653_ & ~new_n38135_;
  assign new_n38137_ = new_n599_ & ~new_n38136_;
  assign new_n38138_ = ~new_n37642_ & ~new_n38137_;
  assign new_n38139_ = ~new_n37663_ & new_n38129_;
  assign new_n38140_ = ~new_n38125_ & new_n38139_;
  assign new_n38141_ = ~new_n38126_ & ~new_n38129_;
  assign new_n38142_ = ~new_n38140_ & ~new_n38141_;
  assign new_n38143_ = new_n599_ & ~new_n38142_;
  assign new_n38144_ = ~new_n38136_ & new_n38143_;
  assign new_n38145_ = ~new_n38138_ & ~new_n38144_;
  assign new_n38146_ = ~new_n37652_ & ~new_n38137_;
  assign new_n38147_ = ~new_n37654_ & new_n38134_;
  assign new_n38148_ = ~new_n38130_ & new_n38147_;
  assign new_n38149_ = ~new_n38131_ & ~new_n38134_;
  assign new_n38150_ = ~new_n38148_ & ~new_n38149_;
  assign new_n38151_ = new_n38137_ & ~new_n38150_;
  assign new_n38152_ = ~new_n38146_ & ~new_n38151_;
  assign new_n38153_ = ~\b[37]  & ~new_n38152_;
  assign new_n38154_ = ~\b[36]  & ~new_n38145_;
  assign new_n38155_ = ~new_n37662_ & ~new_n38137_;
  assign new_n38156_ = ~new_n37672_ & new_n38124_;
  assign new_n38157_ = ~new_n38120_ & new_n38156_;
  assign new_n38158_ = ~new_n38121_ & ~new_n38124_;
  assign new_n38159_ = ~new_n38157_ & ~new_n38158_;
  assign new_n38160_ = new_n599_ & ~new_n38159_;
  assign new_n38161_ = ~new_n38136_ & new_n38160_;
  assign new_n38162_ = ~new_n38155_ & ~new_n38161_;
  assign new_n38163_ = ~\b[35]  & ~new_n38162_;
  assign new_n38164_ = ~new_n37671_ & ~new_n38137_;
  assign new_n38165_ = ~new_n37681_ & new_n38119_;
  assign new_n38166_ = ~new_n38115_ & new_n38165_;
  assign new_n38167_ = ~new_n38116_ & ~new_n38119_;
  assign new_n38168_ = ~new_n38166_ & ~new_n38167_;
  assign new_n38169_ = new_n599_ & ~new_n38168_;
  assign new_n38170_ = ~new_n38136_ & new_n38169_;
  assign new_n38171_ = ~new_n38164_ & ~new_n38170_;
  assign new_n38172_ = ~\b[34]  & ~new_n38171_;
  assign new_n38173_ = ~new_n37680_ & ~new_n38137_;
  assign new_n38174_ = ~new_n37690_ & new_n38114_;
  assign new_n38175_ = ~new_n38110_ & new_n38174_;
  assign new_n38176_ = ~new_n38111_ & ~new_n38114_;
  assign new_n38177_ = ~new_n38175_ & ~new_n38176_;
  assign new_n38178_ = new_n599_ & ~new_n38177_;
  assign new_n38179_ = ~new_n38136_ & new_n38178_;
  assign new_n38180_ = ~new_n38173_ & ~new_n38179_;
  assign new_n38181_ = ~\b[33]  & ~new_n38180_;
  assign new_n38182_ = ~new_n37689_ & ~new_n38137_;
  assign new_n38183_ = ~new_n37699_ & new_n38109_;
  assign new_n38184_ = ~new_n38105_ & new_n38183_;
  assign new_n38185_ = ~new_n38106_ & ~new_n38109_;
  assign new_n38186_ = ~new_n38184_ & ~new_n38185_;
  assign new_n38187_ = new_n599_ & ~new_n38186_;
  assign new_n38188_ = ~new_n38136_ & new_n38187_;
  assign new_n38189_ = ~new_n38182_ & ~new_n38188_;
  assign new_n38190_ = ~\b[32]  & ~new_n38189_;
  assign new_n38191_ = ~new_n37698_ & ~new_n38137_;
  assign new_n38192_ = ~new_n37708_ & new_n38104_;
  assign new_n38193_ = ~new_n38100_ & new_n38192_;
  assign new_n38194_ = ~new_n38101_ & ~new_n38104_;
  assign new_n38195_ = ~new_n38193_ & ~new_n38194_;
  assign new_n38196_ = new_n599_ & ~new_n38195_;
  assign new_n38197_ = ~new_n38136_ & new_n38196_;
  assign new_n38198_ = ~new_n38191_ & ~new_n38197_;
  assign new_n38199_ = ~\b[31]  & ~new_n38198_;
  assign new_n38200_ = ~new_n37707_ & ~new_n38137_;
  assign new_n38201_ = ~new_n37717_ & new_n38099_;
  assign new_n38202_ = ~new_n38095_ & new_n38201_;
  assign new_n38203_ = ~new_n38096_ & ~new_n38099_;
  assign new_n38204_ = ~new_n38202_ & ~new_n38203_;
  assign new_n38205_ = new_n599_ & ~new_n38204_;
  assign new_n38206_ = ~new_n38136_ & new_n38205_;
  assign new_n38207_ = ~new_n38200_ & ~new_n38206_;
  assign new_n38208_ = ~\b[30]  & ~new_n38207_;
  assign new_n38209_ = ~new_n37716_ & ~new_n38137_;
  assign new_n38210_ = ~new_n37726_ & new_n38094_;
  assign new_n38211_ = ~new_n38090_ & new_n38210_;
  assign new_n38212_ = ~new_n38091_ & ~new_n38094_;
  assign new_n38213_ = ~new_n38211_ & ~new_n38212_;
  assign new_n38214_ = new_n599_ & ~new_n38213_;
  assign new_n38215_ = ~new_n38136_ & new_n38214_;
  assign new_n38216_ = ~new_n38209_ & ~new_n38215_;
  assign new_n38217_ = ~\b[29]  & ~new_n38216_;
  assign new_n38218_ = ~new_n37725_ & ~new_n38137_;
  assign new_n38219_ = ~new_n37735_ & new_n38089_;
  assign new_n38220_ = ~new_n38085_ & new_n38219_;
  assign new_n38221_ = ~new_n38086_ & ~new_n38089_;
  assign new_n38222_ = ~new_n38220_ & ~new_n38221_;
  assign new_n38223_ = new_n599_ & ~new_n38222_;
  assign new_n38224_ = ~new_n38136_ & new_n38223_;
  assign new_n38225_ = ~new_n38218_ & ~new_n38224_;
  assign new_n38226_ = ~\b[28]  & ~new_n38225_;
  assign new_n38227_ = ~new_n37734_ & ~new_n38137_;
  assign new_n38228_ = ~new_n37744_ & new_n38084_;
  assign new_n38229_ = ~new_n38080_ & new_n38228_;
  assign new_n38230_ = ~new_n38081_ & ~new_n38084_;
  assign new_n38231_ = ~new_n38229_ & ~new_n38230_;
  assign new_n38232_ = new_n599_ & ~new_n38231_;
  assign new_n38233_ = ~new_n38136_ & new_n38232_;
  assign new_n38234_ = ~new_n38227_ & ~new_n38233_;
  assign new_n38235_ = ~\b[27]  & ~new_n38234_;
  assign new_n38236_ = ~new_n37743_ & ~new_n38137_;
  assign new_n38237_ = ~new_n37753_ & new_n38079_;
  assign new_n38238_ = ~new_n38075_ & new_n38237_;
  assign new_n38239_ = ~new_n38076_ & ~new_n38079_;
  assign new_n38240_ = ~new_n38238_ & ~new_n38239_;
  assign new_n38241_ = new_n599_ & ~new_n38240_;
  assign new_n38242_ = ~new_n38136_ & new_n38241_;
  assign new_n38243_ = ~new_n38236_ & ~new_n38242_;
  assign new_n38244_ = ~\b[26]  & ~new_n38243_;
  assign new_n38245_ = ~new_n37752_ & ~new_n38137_;
  assign new_n38246_ = ~new_n37762_ & new_n38074_;
  assign new_n38247_ = ~new_n38070_ & new_n38246_;
  assign new_n38248_ = ~new_n38071_ & ~new_n38074_;
  assign new_n38249_ = ~new_n38247_ & ~new_n38248_;
  assign new_n38250_ = new_n599_ & ~new_n38249_;
  assign new_n38251_ = ~new_n38136_ & new_n38250_;
  assign new_n38252_ = ~new_n38245_ & ~new_n38251_;
  assign new_n38253_ = ~\b[25]  & ~new_n38252_;
  assign new_n38254_ = ~new_n37761_ & ~new_n38137_;
  assign new_n38255_ = ~new_n37771_ & new_n38069_;
  assign new_n38256_ = ~new_n38065_ & new_n38255_;
  assign new_n38257_ = ~new_n38066_ & ~new_n38069_;
  assign new_n38258_ = ~new_n38256_ & ~new_n38257_;
  assign new_n38259_ = new_n599_ & ~new_n38258_;
  assign new_n38260_ = ~new_n38136_ & new_n38259_;
  assign new_n38261_ = ~new_n38254_ & ~new_n38260_;
  assign new_n38262_ = ~\b[24]  & ~new_n38261_;
  assign new_n38263_ = ~new_n37770_ & ~new_n38137_;
  assign new_n38264_ = ~new_n37780_ & new_n38064_;
  assign new_n38265_ = ~new_n38060_ & new_n38264_;
  assign new_n38266_ = ~new_n38061_ & ~new_n38064_;
  assign new_n38267_ = ~new_n38265_ & ~new_n38266_;
  assign new_n38268_ = new_n599_ & ~new_n38267_;
  assign new_n38269_ = ~new_n38136_ & new_n38268_;
  assign new_n38270_ = ~new_n38263_ & ~new_n38269_;
  assign new_n38271_ = ~\b[23]  & ~new_n38270_;
  assign new_n38272_ = ~new_n37779_ & ~new_n38137_;
  assign new_n38273_ = ~new_n37789_ & new_n38059_;
  assign new_n38274_ = ~new_n38055_ & new_n38273_;
  assign new_n38275_ = ~new_n38056_ & ~new_n38059_;
  assign new_n38276_ = ~new_n38274_ & ~new_n38275_;
  assign new_n38277_ = new_n599_ & ~new_n38276_;
  assign new_n38278_ = ~new_n38136_ & new_n38277_;
  assign new_n38279_ = ~new_n38272_ & ~new_n38278_;
  assign new_n38280_ = ~\b[22]  & ~new_n38279_;
  assign new_n38281_ = ~new_n37788_ & ~new_n38137_;
  assign new_n38282_ = ~new_n37798_ & new_n38054_;
  assign new_n38283_ = ~new_n38050_ & new_n38282_;
  assign new_n38284_ = ~new_n38051_ & ~new_n38054_;
  assign new_n38285_ = ~new_n38283_ & ~new_n38284_;
  assign new_n38286_ = new_n599_ & ~new_n38285_;
  assign new_n38287_ = ~new_n38136_ & new_n38286_;
  assign new_n38288_ = ~new_n38281_ & ~new_n38287_;
  assign new_n38289_ = ~\b[21]  & ~new_n38288_;
  assign new_n38290_ = ~new_n37797_ & ~new_n38137_;
  assign new_n38291_ = ~new_n37807_ & new_n38049_;
  assign new_n38292_ = ~new_n38045_ & new_n38291_;
  assign new_n38293_ = ~new_n38046_ & ~new_n38049_;
  assign new_n38294_ = ~new_n38292_ & ~new_n38293_;
  assign new_n38295_ = new_n599_ & ~new_n38294_;
  assign new_n38296_ = ~new_n38136_ & new_n38295_;
  assign new_n38297_ = ~new_n38290_ & ~new_n38296_;
  assign new_n38298_ = ~\b[20]  & ~new_n38297_;
  assign new_n38299_ = ~new_n37806_ & ~new_n38137_;
  assign new_n38300_ = ~new_n37816_ & new_n38044_;
  assign new_n38301_ = ~new_n38040_ & new_n38300_;
  assign new_n38302_ = ~new_n38041_ & ~new_n38044_;
  assign new_n38303_ = ~new_n38301_ & ~new_n38302_;
  assign new_n38304_ = new_n599_ & ~new_n38303_;
  assign new_n38305_ = ~new_n38136_ & new_n38304_;
  assign new_n38306_ = ~new_n38299_ & ~new_n38305_;
  assign new_n38307_ = ~\b[19]  & ~new_n38306_;
  assign new_n38308_ = ~new_n37815_ & ~new_n38137_;
  assign new_n38309_ = ~new_n37825_ & new_n38039_;
  assign new_n38310_ = ~new_n38035_ & new_n38309_;
  assign new_n38311_ = ~new_n38036_ & ~new_n38039_;
  assign new_n38312_ = ~new_n38310_ & ~new_n38311_;
  assign new_n38313_ = new_n599_ & ~new_n38312_;
  assign new_n38314_ = ~new_n38136_ & new_n38313_;
  assign new_n38315_ = ~new_n38308_ & ~new_n38314_;
  assign new_n38316_ = ~\b[18]  & ~new_n38315_;
  assign new_n38317_ = ~new_n37824_ & ~new_n38137_;
  assign new_n38318_ = ~new_n37834_ & new_n38034_;
  assign new_n38319_ = ~new_n38030_ & new_n38318_;
  assign new_n38320_ = ~new_n38031_ & ~new_n38034_;
  assign new_n38321_ = ~new_n38319_ & ~new_n38320_;
  assign new_n38322_ = new_n599_ & ~new_n38321_;
  assign new_n38323_ = ~new_n38136_ & new_n38322_;
  assign new_n38324_ = ~new_n38317_ & ~new_n38323_;
  assign new_n38325_ = ~\b[17]  & ~new_n38324_;
  assign new_n38326_ = ~new_n37833_ & ~new_n38137_;
  assign new_n38327_ = ~new_n37843_ & new_n38029_;
  assign new_n38328_ = ~new_n38025_ & new_n38327_;
  assign new_n38329_ = ~new_n38026_ & ~new_n38029_;
  assign new_n38330_ = ~new_n38328_ & ~new_n38329_;
  assign new_n38331_ = new_n599_ & ~new_n38330_;
  assign new_n38332_ = ~new_n38136_ & new_n38331_;
  assign new_n38333_ = ~new_n38326_ & ~new_n38332_;
  assign new_n38334_ = ~\b[16]  & ~new_n38333_;
  assign new_n38335_ = ~new_n37842_ & ~new_n38137_;
  assign new_n38336_ = ~new_n37852_ & new_n38024_;
  assign new_n38337_ = ~new_n38020_ & new_n38336_;
  assign new_n38338_ = ~new_n38021_ & ~new_n38024_;
  assign new_n38339_ = ~new_n38337_ & ~new_n38338_;
  assign new_n38340_ = new_n599_ & ~new_n38339_;
  assign new_n38341_ = ~new_n38136_ & new_n38340_;
  assign new_n38342_ = ~new_n38335_ & ~new_n38341_;
  assign new_n38343_ = ~\b[15]  & ~new_n38342_;
  assign new_n38344_ = ~new_n37851_ & ~new_n38137_;
  assign new_n38345_ = ~new_n37861_ & new_n38019_;
  assign new_n38346_ = ~new_n38015_ & new_n38345_;
  assign new_n38347_ = ~new_n38016_ & ~new_n38019_;
  assign new_n38348_ = ~new_n38346_ & ~new_n38347_;
  assign new_n38349_ = new_n599_ & ~new_n38348_;
  assign new_n38350_ = ~new_n38136_ & new_n38349_;
  assign new_n38351_ = ~new_n38344_ & ~new_n38350_;
  assign new_n38352_ = ~\b[14]  & ~new_n38351_;
  assign new_n38353_ = ~new_n37860_ & ~new_n38137_;
  assign new_n38354_ = ~new_n37870_ & new_n38014_;
  assign new_n38355_ = ~new_n38010_ & new_n38354_;
  assign new_n38356_ = ~new_n38011_ & ~new_n38014_;
  assign new_n38357_ = ~new_n38355_ & ~new_n38356_;
  assign new_n38358_ = new_n599_ & ~new_n38357_;
  assign new_n38359_ = ~new_n38136_ & new_n38358_;
  assign new_n38360_ = ~new_n38353_ & ~new_n38359_;
  assign new_n38361_ = ~\b[13]  & ~new_n38360_;
  assign new_n38362_ = ~new_n37869_ & ~new_n38137_;
  assign new_n38363_ = ~new_n37879_ & new_n38009_;
  assign new_n38364_ = ~new_n38005_ & new_n38363_;
  assign new_n38365_ = ~new_n38006_ & ~new_n38009_;
  assign new_n38366_ = ~new_n38364_ & ~new_n38365_;
  assign new_n38367_ = new_n599_ & ~new_n38366_;
  assign new_n38368_ = ~new_n38136_ & new_n38367_;
  assign new_n38369_ = ~new_n38362_ & ~new_n38368_;
  assign new_n38370_ = ~\b[12]  & ~new_n38369_;
  assign new_n38371_ = ~new_n37878_ & ~new_n38137_;
  assign new_n38372_ = ~new_n37888_ & new_n38004_;
  assign new_n38373_ = ~new_n38000_ & new_n38372_;
  assign new_n38374_ = ~new_n38001_ & ~new_n38004_;
  assign new_n38375_ = ~new_n38373_ & ~new_n38374_;
  assign new_n38376_ = new_n599_ & ~new_n38375_;
  assign new_n38377_ = ~new_n38136_ & new_n38376_;
  assign new_n38378_ = ~new_n38371_ & ~new_n38377_;
  assign new_n38379_ = ~\b[11]  & ~new_n38378_;
  assign new_n38380_ = ~new_n37887_ & ~new_n38137_;
  assign new_n38381_ = ~new_n37897_ & new_n37999_;
  assign new_n38382_ = ~new_n37995_ & new_n38381_;
  assign new_n38383_ = ~new_n37996_ & ~new_n37999_;
  assign new_n38384_ = ~new_n38382_ & ~new_n38383_;
  assign new_n38385_ = new_n599_ & ~new_n38384_;
  assign new_n38386_ = ~new_n38136_ & new_n38385_;
  assign new_n38387_ = ~new_n38380_ & ~new_n38386_;
  assign new_n38388_ = ~\b[10]  & ~new_n38387_;
  assign new_n38389_ = ~new_n37896_ & ~new_n38137_;
  assign new_n38390_ = ~new_n37906_ & new_n37994_;
  assign new_n38391_ = ~new_n37990_ & new_n38390_;
  assign new_n38392_ = ~new_n37991_ & ~new_n37994_;
  assign new_n38393_ = ~new_n38391_ & ~new_n38392_;
  assign new_n38394_ = new_n599_ & ~new_n38393_;
  assign new_n38395_ = ~new_n38136_ & new_n38394_;
  assign new_n38396_ = ~new_n38389_ & ~new_n38395_;
  assign new_n38397_ = ~\b[9]  & ~new_n38396_;
  assign new_n38398_ = ~new_n37905_ & ~new_n38137_;
  assign new_n38399_ = ~new_n37915_ & new_n37989_;
  assign new_n38400_ = ~new_n37985_ & new_n38399_;
  assign new_n38401_ = ~new_n37986_ & ~new_n37989_;
  assign new_n38402_ = ~new_n38400_ & ~new_n38401_;
  assign new_n38403_ = new_n599_ & ~new_n38402_;
  assign new_n38404_ = ~new_n38136_ & new_n38403_;
  assign new_n38405_ = ~new_n38398_ & ~new_n38404_;
  assign new_n38406_ = ~\b[8]  & ~new_n38405_;
  assign new_n38407_ = ~new_n37914_ & ~new_n38137_;
  assign new_n38408_ = ~new_n37924_ & new_n37984_;
  assign new_n38409_ = ~new_n37980_ & new_n38408_;
  assign new_n38410_ = ~new_n37981_ & ~new_n37984_;
  assign new_n38411_ = ~new_n38409_ & ~new_n38410_;
  assign new_n38412_ = new_n599_ & ~new_n38411_;
  assign new_n38413_ = ~new_n38136_ & new_n38412_;
  assign new_n38414_ = ~new_n38407_ & ~new_n38413_;
  assign new_n38415_ = ~\b[7]  & ~new_n38414_;
  assign new_n38416_ = ~new_n37923_ & ~new_n38137_;
  assign new_n38417_ = ~new_n37933_ & new_n37979_;
  assign new_n38418_ = ~new_n37975_ & new_n38417_;
  assign new_n38419_ = ~new_n37976_ & ~new_n37979_;
  assign new_n38420_ = ~new_n38418_ & ~new_n38419_;
  assign new_n38421_ = new_n599_ & ~new_n38420_;
  assign new_n38422_ = ~new_n38136_ & new_n38421_;
  assign new_n38423_ = ~new_n38416_ & ~new_n38422_;
  assign new_n38424_ = ~\b[6]  & ~new_n38423_;
  assign new_n38425_ = ~new_n37932_ & ~new_n38137_;
  assign new_n38426_ = ~new_n37942_ & new_n37974_;
  assign new_n38427_ = ~new_n37970_ & new_n38426_;
  assign new_n38428_ = ~new_n37971_ & ~new_n37974_;
  assign new_n38429_ = ~new_n38427_ & ~new_n38428_;
  assign new_n38430_ = new_n599_ & ~new_n38429_;
  assign new_n38431_ = ~new_n38136_ & new_n38430_;
  assign new_n38432_ = ~new_n38425_ & ~new_n38431_;
  assign new_n38433_ = ~\b[5]  & ~new_n38432_;
  assign new_n38434_ = ~new_n37941_ & ~new_n38137_;
  assign new_n38435_ = ~new_n37950_ & new_n37969_;
  assign new_n38436_ = ~new_n37965_ & new_n38435_;
  assign new_n38437_ = ~new_n37966_ & ~new_n37969_;
  assign new_n38438_ = ~new_n38436_ & ~new_n38437_;
  assign new_n38439_ = new_n599_ & ~new_n38438_;
  assign new_n38440_ = ~new_n38136_ & new_n38439_;
  assign new_n38441_ = ~new_n38434_ & ~new_n38440_;
  assign new_n38442_ = ~\b[4]  & ~new_n38441_;
  assign new_n38443_ = ~new_n37949_ & ~new_n38137_;
  assign new_n38444_ = ~new_n37960_ & new_n37964_;
  assign new_n38445_ = ~new_n37959_ & new_n38444_;
  assign new_n38446_ = ~new_n37961_ & ~new_n37964_;
  assign new_n38447_ = ~new_n38445_ & ~new_n38446_;
  assign new_n38448_ = new_n599_ & ~new_n38447_;
  assign new_n38449_ = ~new_n38136_ & new_n38448_;
  assign new_n38450_ = ~new_n38443_ & ~new_n38449_;
  assign new_n38451_ = ~\b[3]  & ~new_n38450_;
  assign new_n38452_ = ~new_n37954_ & ~new_n38137_;
  assign new_n38453_ = new_n9826_ & ~new_n37957_;
  assign new_n38454_ = ~new_n37955_ & new_n38453_;
  assign new_n38455_ = new_n599_ & ~new_n38454_;
  assign new_n38456_ = ~new_n37959_ & new_n38455_;
  assign new_n38457_ = ~new_n38136_ & new_n38456_;
  assign new_n38458_ = ~new_n38452_ & ~new_n38457_;
  assign new_n38459_ = ~\b[2]  & ~new_n38458_;
  assign new_n38460_ = new_n10332_ & ~new_n38136_;
  assign new_n38461_ = \a[27]  & ~new_n38460_;
  assign new_n38462_ = new_n10337_ & ~new_n38136_;
  assign new_n38463_ = ~new_n38461_ & ~new_n38462_;
  assign new_n38464_ = \b[1]  & ~new_n38463_;
  assign new_n38465_ = ~\b[1]  & ~new_n38462_;
  assign new_n38466_ = ~new_n38461_ & new_n38465_;
  assign new_n38467_ = ~new_n38464_ & ~new_n38466_;
  assign new_n38468_ = ~new_n10344_ & ~new_n38467_;
  assign new_n38469_ = ~\b[1]  & ~new_n38463_;
  assign new_n38470_ = ~new_n38468_ & ~new_n38469_;
  assign new_n38471_ = \b[2]  & ~new_n38457_;
  assign new_n38472_ = ~new_n38452_ & new_n38471_;
  assign new_n38473_ = ~new_n38459_ & ~new_n38472_;
  assign new_n38474_ = ~new_n38470_ & new_n38473_;
  assign new_n38475_ = ~new_n38459_ & ~new_n38474_;
  assign new_n38476_ = \b[3]  & ~new_n38449_;
  assign new_n38477_ = ~new_n38443_ & new_n38476_;
  assign new_n38478_ = ~new_n38451_ & ~new_n38477_;
  assign new_n38479_ = ~new_n38475_ & new_n38478_;
  assign new_n38480_ = ~new_n38451_ & ~new_n38479_;
  assign new_n38481_ = \b[4]  & ~new_n38440_;
  assign new_n38482_ = ~new_n38434_ & new_n38481_;
  assign new_n38483_ = ~new_n38442_ & ~new_n38482_;
  assign new_n38484_ = ~new_n38480_ & new_n38483_;
  assign new_n38485_ = ~new_n38442_ & ~new_n38484_;
  assign new_n38486_ = \b[5]  & ~new_n38431_;
  assign new_n38487_ = ~new_n38425_ & new_n38486_;
  assign new_n38488_ = ~new_n38433_ & ~new_n38487_;
  assign new_n38489_ = ~new_n38485_ & new_n38488_;
  assign new_n38490_ = ~new_n38433_ & ~new_n38489_;
  assign new_n38491_ = \b[6]  & ~new_n38422_;
  assign new_n38492_ = ~new_n38416_ & new_n38491_;
  assign new_n38493_ = ~new_n38424_ & ~new_n38492_;
  assign new_n38494_ = ~new_n38490_ & new_n38493_;
  assign new_n38495_ = ~new_n38424_ & ~new_n38494_;
  assign new_n38496_ = \b[7]  & ~new_n38413_;
  assign new_n38497_ = ~new_n38407_ & new_n38496_;
  assign new_n38498_ = ~new_n38415_ & ~new_n38497_;
  assign new_n38499_ = ~new_n38495_ & new_n38498_;
  assign new_n38500_ = ~new_n38415_ & ~new_n38499_;
  assign new_n38501_ = \b[8]  & ~new_n38404_;
  assign new_n38502_ = ~new_n38398_ & new_n38501_;
  assign new_n38503_ = ~new_n38406_ & ~new_n38502_;
  assign new_n38504_ = ~new_n38500_ & new_n38503_;
  assign new_n38505_ = ~new_n38406_ & ~new_n38504_;
  assign new_n38506_ = \b[9]  & ~new_n38395_;
  assign new_n38507_ = ~new_n38389_ & new_n38506_;
  assign new_n38508_ = ~new_n38397_ & ~new_n38507_;
  assign new_n38509_ = ~new_n38505_ & new_n38508_;
  assign new_n38510_ = ~new_n38397_ & ~new_n38509_;
  assign new_n38511_ = \b[10]  & ~new_n38386_;
  assign new_n38512_ = ~new_n38380_ & new_n38511_;
  assign new_n38513_ = ~new_n38388_ & ~new_n38512_;
  assign new_n38514_ = ~new_n38510_ & new_n38513_;
  assign new_n38515_ = ~new_n38388_ & ~new_n38514_;
  assign new_n38516_ = \b[11]  & ~new_n38377_;
  assign new_n38517_ = ~new_n38371_ & new_n38516_;
  assign new_n38518_ = ~new_n38379_ & ~new_n38517_;
  assign new_n38519_ = ~new_n38515_ & new_n38518_;
  assign new_n38520_ = ~new_n38379_ & ~new_n38519_;
  assign new_n38521_ = \b[12]  & ~new_n38368_;
  assign new_n38522_ = ~new_n38362_ & new_n38521_;
  assign new_n38523_ = ~new_n38370_ & ~new_n38522_;
  assign new_n38524_ = ~new_n38520_ & new_n38523_;
  assign new_n38525_ = ~new_n38370_ & ~new_n38524_;
  assign new_n38526_ = \b[13]  & ~new_n38359_;
  assign new_n38527_ = ~new_n38353_ & new_n38526_;
  assign new_n38528_ = ~new_n38361_ & ~new_n38527_;
  assign new_n38529_ = ~new_n38525_ & new_n38528_;
  assign new_n38530_ = ~new_n38361_ & ~new_n38529_;
  assign new_n38531_ = \b[14]  & ~new_n38350_;
  assign new_n38532_ = ~new_n38344_ & new_n38531_;
  assign new_n38533_ = ~new_n38352_ & ~new_n38532_;
  assign new_n38534_ = ~new_n38530_ & new_n38533_;
  assign new_n38535_ = ~new_n38352_ & ~new_n38534_;
  assign new_n38536_ = \b[15]  & ~new_n38341_;
  assign new_n38537_ = ~new_n38335_ & new_n38536_;
  assign new_n38538_ = ~new_n38343_ & ~new_n38537_;
  assign new_n38539_ = ~new_n38535_ & new_n38538_;
  assign new_n38540_ = ~new_n38343_ & ~new_n38539_;
  assign new_n38541_ = \b[16]  & ~new_n38332_;
  assign new_n38542_ = ~new_n38326_ & new_n38541_;
  assign new_n38543_ = ~new_n38334_ & ~new_n38542_;
  assign new_n38544_ = ~new_n38540_ & new_n38543_;
  assign new_n38545_ = ~new_n38334_ & ~new_n38544_;
  assign new_n38546_ = \b[17]  & ~new_n38323_;
  assign new_n38547_ = ~new_n38317_ & new_n38546_;
  assign new_n38548_ = ~new_n38325_ & ~new_n38547_;
  assign new_n38549_ = ~new_n38545_ & new_n38548_;
  assign new_n38550_ = ~new_n38325_ & ~new_n38549_;
  assign new_n38551_ = \b[18]  & ~new_n38314_;
  assign new_n38552_ = ~new_n38308_ & new_n38551_;
  assign new_n38553_ = ~new_n38316_ & ~new_n38552_;
  assign new_n38554_ = ~new_n38550_ & new_n38553_;
  assign new_n38555_ = ~new_n38316_ & ~new_n38554_;
  assign new_n38556_ = \b[19]  & ~new_n38305_;
  assign new_n38557_ = ~new_n38299_ & new_n38556_;
  assign new_n38558_ = ~new_n38307_ & ~new_n38557_;
  assign new_n38559_ = ~new_n38555_ & new_n38558_;
  assign new_n38560_ = ~new_n38307_ & ~new_n38559_;
  assign new_n38561_ = \b[20]  & ~new_n38296_;
  assign new_n38562_ = ~new_n38290_ & new_n38561_;
  assign new_n38563_ = ~new_n38298_ & ~new_n38562_;
  assign new_n38564_ = ~new_n38560_ & new_n38563_;
  assign new_n38565_ = ~new_n38298_ & ~new_n38564_;
  assign new_n38566_ = \b[21]  & ~new_n38287_;
  assign new_n38567_ = ~new_n38281_ & new_n38566_;
  assign new_n38568_ = ~new_n38289_ & ~new_n38567_;
  assign new_n38569_ = ~new_n38565_ & new_n38568_;
  assign new_n38570_ = ~new_n38289_ & ~new_n38569_;
  assign new_n38571_ = \b[22]  & ~new_n38278_;
  assign new_n38572_ = ~new_n38272_ & new_n38571_;
  assign new_n38573_ = ~new_n38280_ & ~new_n38572_;
  assign new_n38574_ = ~new_n38570_ & new_n38573_;
  assign new_n38575_ = ~new_n38280_ & ~new_n38574_;
  assign new_n38576_ = \b[23]  & ~new_n38269_;
  assign new_n38577_ = ~new_n38263_ & new_n38576_;
  assign new_n38578_ = ~new_n38271_ & ~new_n38577_;
  assign new_n38579_ = ~new_n38575_ & new_n38578_;
  assign new_n38580_ = ~new_n38271_ & ~new_n38579_;
  assign new_n38581_ = \b[24]  & ~new_n38260_;
  assign new_n38582_ = ~new_n38254_ & new_n38581_;
  assign new_n38583_ = ~new_n38262_ & ~new_n38582_;
  assign new_n38584_ = ~new_n38580_ & new_n38583_;
  assign new_n38585_ = ~new_n38262_ & ~new_n38584_;
  assign new_n38586_ = \b[25]  & ~new_n38251_;
  assign new_n38587_ = ~new_n38245_ & new_n38586_;
  assign new_n38588_ = ~new_n38253_ & ~new_n38587_;
  assign new_n38589_ = ~new_n38585_ & new_n38588_;
  assign new_n38590_ = ~new_n38253_ & ~new_n38589_;
  assign new_n38591_ = \b[26]  & ~new_n38242_;
  assign new_n38592_ = ~new_n38236_ & new_n38591_;
  assign new_n38593_ = ~new_n38244_ & ~new_n38592_;
  assign new_n38594_ = ~new_n38590_ & new_n38593_;
  assign new_n38595_ = ~new_n38244_ & ~new_n38594_;
  assign new_n38596_ = \b[27]  & ~new_n38233_;
  assign new_n38597_ = ~new_n38227_ & new_n38596_;
  assign new_n38598_ = ~new_n38235_ & ~new_n38597_;
  assign new_n38599_ = ~new_n38595_ & new_n38598_;
  assign new_n38600_ = ~new_n38235_ & ~new_n38599_;
  assign new_n38601_ = \b[28]  & ~new_n38224_;
  assign new_n38602_ = ~new_n38218_ & new_n38601_;
  assign new_n38603_ = ~new_n38226_ & ~new_n38602_;
  assign new_n38604_ = ~new_n38600_ & new_n38603_;
  assign new_n38605_ = ~new_n38226_ & ~new_n38604_;
  assign new_n38606_ = \b[29]  & ~new_n38215_;
  assign new_n38607_ = ~new_n38209_ & new_n38606_;
  assign new_n38608_ = ~new_n38217_ & ~new_n38607_;
  assign new_n38609_ = ~new_n38605_ & new_n38608_;
  assign new_n38610_ = ~new_n38217_ & ~new_n38609_;
  assign new_n38611_ = \b[30]  & ~new_n38206_;
  assign new_n38612_ = ~new_n38200_ & new_n38611_;
  assign new_n38613_ = ~new_n38208_ & ~new_n38612_;
  assign new_n38614_ = ~new_n38610_ & new_n38613_;
  assign new_n38615_ = ~new_n38208_ & ~new_n38614_;
  assign new_n38616_ = \b[31]  & ~new_n38197_;
  assign new_n38617_ = ~new_n38191_ & new_n38616_;
  assign new_n38618_ = ~new_n38199_ & ~new_n38617_;
  assign new_n38619_ = ~new_n38615_ & new_n38618_;
  assign new_n38620_ = ~new_n38199_ & ~new_n38619_;
  assign new_n38621_ = \b[32]  & ~new_n38188_;
  assign new_n38622_ = ~new_n38182_ & new_n38621_;
  assign new_n38623_ = ~new_n38190_ & ~new_n38622_;
  assign new_n38624_ = ~new_n38620_ & new_n38623_;
  assign new_n38625_ = ~new_n38190_ & ~new_n38624_;
  assign new_n38626_ = \b[33]  & ~new_n38179_;
  assign new_n38627_ = ~new_n38173_ & new_n38626_;
  assign new_n38628_ = ~new_n38181_ & ~new_n38627_;
  assign new_n38629_ = ~new_n38625_ & new_n38628_;
  assign new_n38630_ = ~new_n38181_ & ~new_n38629_;
  assign new_n38631_ = \b[34]  & ~new_n38170_;
  assign new_n38632_ = ~new_n38164_ & new_n38631_;
  assign new_n38633_ = ~new_n38172_ & ~new_n38632_;
  assign new_n38634_ = ~new_n38630_ & new_n38633_;
  assign new_n38635_ = ~new_n38172_ & ~new_n38634_;
  assign new_n38636_ = \b[35]  & ~new_n38161_;
  assign new_n38637_ = ~new_n38155_ & new_n38636_;
  assign new_n38638_ = ~new_n38163_ & ~new_n38637_;
  assign new_n38639_ = ~new_n38635_ & new_n38638_;
  assign new_n38640_ = ~new_n38163_ & ~new_n38639_;
  assign new_n38641_ = \b[36]  & ~new_n38144_;
  assign new_n38642_ = ~new_n38138_ & new_n38641_;
  assign new_n38643_ = ~new_n38154_ & ~new_n38642_;
  assign new_n38644_ = ~new_n38640_ & new_n38643_;
  assign new_n38645_ = ~new_n38154_ & ~new_n38644_;
  assign new_n38646_ = \b[37]  & ~new_n38146_;
  assign new_n38647_ = ~new_n38151_ & new_n38646_;
  assign new_n38648_ = ~new_n38153_ & ~new_n38647_;
  assign new_n38649_ = ~new_n38645_ & new_n38648_;
  assign new_n38650_ = ~new_n38153_ & ~new_n38649_;
  assign new_n38651_ = new_n10530_ & ~new_n38650_;
  assign new_n38652_ = ~new_n38145_ & ~new_n38651_;
  assign new_n38653_ = ~new_n38163_ & new_n38643_;
  assign new_n38654_ = ~new_n38639_ & new_n38653_;
  assign new_n38655_ = ~new_n38640_ & ~new_n38643_;
  assign new_n38656_ = ~new_n38654_ & ~new_n38655_;
  assign new_n38657_ = new_n10530_ & ~new_n38656_;
  assign new_n38658_ = ~new_n38650_ & new_n38657_;
  assign new_n38659_ = ~new_n38652_ & ~new_n38658_;
  assign new_n38660_ = ~\b[37]  & ~new_n38659_;
  assign new_n38661_ = ~new_n38162_ & ~new_n38651_;
  assign new_n38662_ = ~new_n38172_ & new_n38638_;
  assign new_n38663_ = ~new_n38634_ & new_n38662_;
  assign new_n38664_ = ~new_n38635_ & ~new_n38638_;
  assign new_n38665_ = ~new_n38663_ & ~new_n38664_;
  assign new_n38666_ = new_n10530_ & ~new_n38665_;
  assign new_n38667_ = ~new_n38650_ & new_n38666_;
  assign new_n38668_ = ~new_n38661_ & ~new_n38667_;
  assign new_n38669_ = ~\b[36]  & ~new_n38668_;
  assign new_n38670_ = ~new_n38171_ & ~new_n38651_;
  assign new_n38671_ = ~new_n38181_ & new_n38633_;
  assign new_n38672_ = ~new_n38629_ & new_n38671_;
  assign new_n38673_ = ~new_n38630_ & ~new_n38633_;
  assign new_n38674_ = ~new_n38672_ & ~new_n38673_;
  assign new_n38675_ = new_n10530_ & ~new_n38674_;
  assign new_n38676_ = ~new_n38650_ & new_n38675_;
  assign new_n38677_ = ~new_n38670_ & ~new_n38676_;
  assign new_n38678_ = ~\b[35]  & ~new_n38677_;
  assign new_n38679_ = ~new_n38180_ & ~new_n38651_;
  assign new_n38680_ = ~new_n38190_ & new_n38628_;
  assign new_n38681_ = ~new_n38624_ & new_n38680_;
  assign new_n38682_ = ~new_n38625_ & ~new_n38628_;
  assign new_n38683_ = ~new_n38681_ & ~new_n38682_;
  assign new_n38684_ = new_n10530_ & ~new_n38683_;
  assign new_n38685_ = ~new_n38650_ & new_n38684_;
  assign new_n38686_ = ~new_n38679_ & ~new_n38685_;
  assign new_n38687_ = ~\b[34]  & ~new_n38686_;
  assign new_n38688_ = ~new_n38189_ & ~new_n38651_;
  assign new_n38689_ = ~new_n38199_ & new_n38623_;
  assign new_n38690_ = ~new_n38619_ & new_n38689_;
  assign new_n38691_ = ~new_n38620_ & ~new_n38623_;
  assign new_n38692_ = ~new_n38690_ & ~new_n38691_;
  assign new_n38693_ = new_n10530_ & ~new_n38692_;
  assign new_n38694_ = ~new_n38650_ & new_n38693_;
  assign new_n38695_ = ~new_n38688_ & ~new_n38694_;
  assign new_n38696_ = ~\b[33]  & ~new_n38695_;
  assign new_n38697_ = ~new_n38198_ & ~new_n38651_;
  assign new_n38698_ = ~new_n38208_ & new_n38618_;
  assign new_n38699_ = ~new_n38614_ & new_n38698_;
  assign new_n38700_ = ~new_n38615_ & ~new_n38618_;
  assign new_n38701_ = ~new_n38699_ & ~new_n38700_;
  assign new_n38702_ = new_n10530_ & ~new_n38701_;
  assign new_n38703_ = ~new_n38650_ & new_n38702_;
  assign new_n38704_ = ~new_n38697_ & ~new_n38703_;
  assign new_n38705_ = ~\b[32]  & ~new_n38704_;
  assign new_n38706_ = ~new_n38207_ & ~new_n38651_;
  assign new_n38707_ = ~new_n38217_ & new_n38613_;
  assign new_n38708_ = ~new_n38609_ & new_n38707_;
  assign new_n38709_ = ~new_n38610_ & ~new_n38613_;
  assign new_n38710_ = ~new_n38708_ & ~new_n38709_;
  assign new_n38711_ = new_n10530_ & ~new_n38710_;
  assign new_n38712_ = ~new_n38650_ & new_n38711_;
  assign new_n38713_ = ~new_n38706_ & ~new_n38712_;
  assign new_n38714_ = ~\b[31]  & ~new_n38713_;
  assign new_n38715_ = ~new_n38216_ & ~new_n38651_;
  assign new_n38716_ = ~new_n38226_ & new_n38608_;
  assign new_n38717_ = ~new_n38604_ & new_n38716_;
  assign new_n38718_ = ~new_n38605_ & ~new_n38608_;
  assign new_n38719_ = ~new_n38717_ & ~new_n38718_;
  assign new_n38720_ = new_n10530_ & ~new_n38719_;
  assign new_n38721_ = ~new_n38650_ & new_n38720_;
  assign new_n38722_ = ~new_n38715_ & ~new_n38721_;
  assign new_n38723_ = ~\b[30]  & ~new_n38722_;
  assign new_n38724_ = ~new_n38225_ & ~new_n38651_;
  assign new_n38725_ = ~new_n38235_ & new_n38603_;
  assign new_n38726_ = ~new_n38599_ & new_n38725_;
  assign new_n38727_ = ~new_n38600_ & ~new_n38603_;
  assign new_n38728_ = ~new_n38726_ & ~new_n38727_;
  assign new_n38729_ = new_n10530_ & ~new_n38728_;
  assign new_n38730_ = ~new_n38650_ & new_n38729_;
  assign new_n38731_ = ~new_n38724_ & ~new_n38730_;
  assign new_n38732_ = ~\b[29]  & ~new_n38731_;
  assign new_n38733_ = ~new_n38234_ & ~new_n38651_;
  assign new_n38734_ = ~new_n38244_ & new_n38598_;
  assign new_n38735_ = ~new_n38594_ & new_n38734_;
  assign new_n38736_ = ~new_n38595_ & ~new_n38598_;
  assign new_n38737_ = ~new_n38735_ & ~new_n38736_;
  assign new_n38738_ = new_n10530_ & ~new_n38737_;
  assign new_n38739_ = ~new_n38650_ & new_n38738_;
  assign new_n38740_ = ~new_n38733_ & ~new_n38739_;
  assign new_n38741_ = ~\b[28]  & ~new_n38740_;
  assign new_n38742_ = ~new_n38243_ & ~new_n38651_;
  assign new_n38743_ = ~new_n38253_ & new_n38593_;
  assign new_n38744_ = ~new_n38589_ & new_n38743_;
  assign new_n38745_ = ~new_n38590_ & ~new_n38593_;
  assign new_n38746_ = ~new_n38744_ & ~new_n38745_;
  assign new_n38747_ = new_n10530_ & ~new_n38746_;
  assign new_n38748_ = ~new_n38650_ & new_n38747_;
  assign new_n38749_ = ~new_n38742_ & ~new_n38748_;
  assign new_n38750_ = ~\b[27]  & ~new_n38749_;
  assign new_n38751_ = ~new_n38252_ & ~new_n38651_;
  assign new_n38752_ = ~new_n38262_ & new_n38588_;
  assign new_n38753_ = ~new_n38584_ & new_n38752_;
  assign new_n38754_ = ~new_n38585_ & ~new_n38588_;
  assign new_n38755_ = ~new_n38753_ & ~new_n38754_;
  assign new_n38756_ = new_n10530_ & ~new_n38755_;
  assign new_n38757_ = ~new_n38650_ & new_n38756_;
  assign new_n38758_ = ~new_n38751_ & ~new_n38757_;
  assign new_n38759_ = ~\b[26]  & ~new_n38758_;
  assign new_n38760_ = ~new_n38261_ & ~new_n38651_;
  assign new_n38761_ = ~new_n38271_ & new_n38583_;
  assign new_n38762_ = ~new_n38579_ & new_n38761_;
  assign new_n38763_ = ~new_n38580_ & ~new_n38583_;
  assign new_n38764_ = ~new_n38762_ & ~new_n38763_;
  assign new_n38765_ = new_n10530_ & ~new_n38764_;
  assign new_n38766_ = ~new_n38650_ & new_n38765_;
  assign new_n38767_ = ~new_n38760_ & ~new_n38766_;
  assign new_n38768_ = ~\b[25]  & ~new_n38767_;
  assign new_n38769_ = ~new_n38270_ & ~new_n38651_;
  assign new_n38770_ = ~new_n38280_ & new_n38578_;
  assign new_n38771_ = ~new_n38574_ & new_n38770_;
  assign new_n38772_ = ~new_n38575_ & ~new_n38578_;
  assign new_n38773_ = ~new_n38771_ & ~new_n38772_;
  assign new_n38774_ = new_n10530_ & ~new_n38773_;
  assign new_n38775_ = ~new_n38650_ & new_n38774_;
  assign new_n38776_ = ~new_n38769_ & ~new_n38775_;
  assign new_n38777_ = ~\b[24]  & ~new_n38776_;
  assign new_n38778_ = ~new_n38279_ & ~new_n38651_;
  assign new_n38779_ = ~new_n38289_ & new_n38573_;
  assign new_n38780_ = ~new_n38569_ & new_n38779_;
  assign new_n38781_ = ~new_n38570_ & ~new_n38573_;
  assign new_n38782_ = ~new_n38780_ & ~new_n38781_;
  assign new_n38783_ = new_n10530_ & ~new_n38782_;
  assign new_n38784_ = ~new_n38650_ & new_n38783_;
  assign new_n38785_ = ~new_n38778_ & ~new_n38784_;
  assign new_n38786_ = ~\b[23]  & ~new_n38785_;
  assign new_n38787_ = ~new_n38288_ & ~new_n38651_;
  assign new_n38788_ = ~new_n38298_ & new_n38568_;
  assign new_n38789_ = ~new_n38564_ & new_n38788_;
  assign new_n38790_ = ~new_n38565_ & ~new_n38568_;
  assign new_n38791_ = ~new_n38789_ & ~new_n38790_;
  assign new_n38792_ = new_n10530_ & ~new_n38791_;
  assign new_n38793_ = ~new_n38650_ & new_n38792_;
  assign new_n38794_ = ~new_n38787_ & ~new_n38793_;
  assign new_n38795_ = ~\b[22]  & ~new_n38794_;
  assign new_n38796_ = ~new_n38297_ & ~new_n38651_;
  assign new_n38797_ = ~new_n38307_ & new_n38563_;
  assign new_n38798_ = ~new_n38559_ & new_n38797_;
  assign new_n38799_ = ~new_n38560_ & ~new_n38563_;
  assign new_n38800_ = ~new_n38798_ & ~new_n38799_;
  assign new_n38801_ = new_n10530_ & ~new_n38800_;
  assign new_n38802_ = ~new_n38650_ & new_n38801_;
  assign new_n38803_ = ~new_n38796_ & ~new_n38802_;
  assign new_n38804_ = ~\b[21]  & ~new_n38803_;
  assign new_n38805_ = ~new_n38306_ & ~new_n38651_;
  assign new_n38806_ = ~new_n38316_ & new_n38558_;
  assign new_n38807_ = ~new_n38554_ & new_n38806_;
  assign new_n38808_ = ~new_n38555_ & ~new_n38558_;
  assign new_n38809_ = ~new_n38807_ & ~new_n38808_;
  assign new_n38810_ = new_n10530_ & ~new_n38809_;
  assign new_n38811_ = ~new_n38650_ & new_n38810_;
  assign new_n38812_ = ~new_n38805_ & ~new_n38811_;
  assign new_n38813_ = ~\b[20]  & ~new_n38812_;
  assign new_n38814_ = ~new_n38315_ & ~new_n38651_;
  assign new_n38815_ = ~new_n38325_ & new_n38553_;
  assign new_n38816_ = ~new_n38549_ & new_n38815_;
  assign new_n38817_ = ~new_n38550_ & ~new_n38553_;
  assign new_n38818_ = ~new_n38816_ & ~new_n38817_;
  assign new_n38819_ = new_n10530_ & ~new_n38818_;
  assign new_n38820_ = ~new_n38650_ & new_n38819_;
  assign new_n38821_ = ~new_n38814_ & ~new_n38820_;
  assign new_n38822_ = ~\b[19]  & ~new_n38821_;
  assign new_n38823_ = ~new_n38324_ & ~new_n38651_;
  assign new_n38824_ = ~new_n38334_ & new_n38548_;
  assign new_n38825_ = ~new_n38544_ & new_n38824_;
  assign new_n38826_ = ~new_n38545_ & ~new_n38548_;
  assign new_n38827_ = ~new_n38825_ & ~new_n38826_;
  assign new_n38828_ = new_n10530_ & ~new_n38827_;
  assign new_n38829_ = ~new_n38650_ & new_n38828_;
  assign new_n38830_ = ~new_n38823_ & ~new_n38829_;
  assign new_n38831_ = ~\b[18]  & ~new_n38830_;
  assign new_n38832_ = ~new_n38333_ & ~new_n38651_;
  assign new_n38833_ = ~new_n38343_ & new_n38543_;
  assign new_n38834_ = ~new_n38539_ & new_n38833_;
  assign new_n38835_ = ~new_n38540_ & ~new_n38543_;
  assign new_n38836_ = ~new_n38834_ & ~new_n38835_;
  assign new_n38837_ = new_n10530_ & ~new_n38836_;
  assign new_n38838_ = ~new_n38650_ & new_n38837_;
  assign new_n38839_ = ~new_n38832_ & ~new_n38838_;
  assign new_n38840_ = ~\b[17]  & ~new_n38839_;
  assign new_n38841_ = ~new_n38342_ & ~new_n38651_;
  assign new_n38842_ = ~new_n38352_ & new_n38538_;
  assign new_n38843_ = ~new_n38534_ & new_n38842_;
  assign new_n38844_ = ~new_n38535_ & ~new_n38538_;
  assign new_n38845_ = ~new_n38843_ & ~new_n38844_;
  assign new_n38846_ = new_n10530_ & ~new_n38845_;
  assign new_n38847_ = ~new_n38650_ & new_n38846_;
  assign new_n38848_ = ~new_n38841_ & ~new_n38847_;
  assign new_n38849_ = ~\b[16]  & ~new_n38848_;
  assign new_n38850_ = ~new_n38351_ & ~new_n38651_;
  assign new_n38851_ = ~new_n38361_ & new_n38533_;
  assign new_n38852_ = ~new_n38529_ & new_n38851_;
  assign new_n38853_ = ~new_n38530_ & ~new_n38533_;
  assign new_n38854_ = ~new_n38852_ & ~new_n38853_;
  assign new_n38855_ = new_n10530_ & ~new_n38854_;
  assign new_n38856_ = ~new_n38650_ & new_n38855_;
  assign new_n38857_ = ~new_n38850_ & ~new_n38856_;
  assign new_n38858_ = ~\b[15]  & ~new_n38857_;
  assign new_n38859_ = ~new_n38360_ & ~new_n38651_;
  assign new_n38860_ = ~new_n38370_ & new_n38528_;
  assign new_n38861_ = ~new_n38524_ & new_n38860_;
  assign new_n38862_ = ~new_n38525_ & ~new_n38528_;
  assign new_n38863_ = ~new_n38861_ & ~new_n38862_;
  assign new_n38864_ = new_n10530_ & ~new_n38863_;
  assign new_n38865_ = ~new_n38650_ & new_n38864_;
  assign new_n38866_ = ~new_n38859_ & ~new_n38865_;
  assign new_n38867_ = ~\b[14]  & ~new_n38866_;
  assign new_n38868_ = ~new_n38369_ & ~new_n38651_;
  assign new_n38869_ = ~new_n38379_ & new_n38523_;
  assign new_n38870_ = ~new_n38519_ & new_n38869_;
  assign new_n38871_ = ~new_n38520_ & ~new_n38523_;
  assign new_n38872_ = ~new_n38870_ & ~new_n38871_;
  assign new_n38873_ = new_n10530_ & ~new_n38872_;
  assign new_n38874_ = ~new_n38650_ & new_n38873_;
  assign new_n38875_ = ~new_n38868_ & ~new_n38874_;
  assign new_n38876_ = ~\b[13]  & ~new_n38875_;
  assign new_n38877_ = ~new_n38378_ & ~new_n38651_;
  assign new_n38878_ = ~new_n38388_ & new_n38518_;
  assign new_n38879_ = ~new_n38514_ & new_n38878_;
  assign new_n38880_ = ~new_n38515_ & ~new_n38518_;
  assign new_n38881_ = ~new_n38879_ & ~new_n38880_;
  assign new_n38882_ = new_n10530_ & ~new_n38881_;
  assign new_n38883_ = ~new_n38650_ & new_n38882_;
  assign new_n38884_ = ~new_n38877_ & ~new_n38883_;
  assign new_n38885_ = ~\b[12]  & ~new_n38884_;
  assign new_n38886_ = ~new_n38387_ & ~new_n38651_;
  assign new_n38887_ = ~new_n38397_ & new_n38513_;
  assign new_n38888_ = ~new_n38509_ & new_n38887_;
  assign new_n38889_ = ~new_n38510_ & ~new_n38513_;
  assign new_n38890_ = ~new_n38888_ & ~new_n38889_;
  assign new_n38891_ = new_n10530_ & ~new_n38890_;
  assign new_n38892_ = ~new_n38650_ & new_n38891_;
  assign new_n38893_ = ~new_n38886_ & ~new_n38892_;
  assign new_n38894_ = ~\b[11]  & ~new_n38893_;
  assign new_n38895_ = ~new_n38396_ & ~new_n38651_;
  assign new_n38896_ = ~new_n38406_ & new_n38508_;
  assign new_n38897_ = ~new_n38504_ & new_n38896_;
  assign new_n38898_ = ~new_n38505_ & ~new_n38508_;
  assign new_n38899_ = ~new_n38897_ & ~new_n38898_;
  assign new_n38900_ = new_n10530_ & ~new_n38899_;
  assign new_n38901_ = ~new_n38650_ & new_n38900_;
  assign new_n38902_ = ~new_n38895_ & ~new_n38901_;
  assign new_n38903_ = ~\b[10]  & ~new_n38902_;
  assign new_n38904_ = ~new_n38405_ & ~new_n38651_;
  assign new_n38905_ = ~new_n38415_ & new_n38503_;
  assign new_n38906_ = ~new_n38499_ & new_n38905_;
  assign new_n38907_ = ~new_n38500_ & ~new_n38503_;
  assign new_n38908_ = ~new_n38906_ & ~new_n38907_;
  assign new_n38909_ = new_n10530_ & ~new_n38908_;
  assign new_n38910_ = ~new_n38650_ & new_n38909_;
  assign new_n38911_ = ~new_n38904_ & ~new_n38910_;
  assign new_n38912_ = ~\b[9]  & ~new_n38911_;
  assign new_n38913_ = ~new_n38414_ & ~new_n38651_;
  assign new_n38914_ = ~new_n38424_ & new_n38498_;
  assign new_n38915_ = ~new_n38494_ & new_n38914_;
  assign new_n38916_ = ~new_n38495_ & ~new_n38498_;
  assign new_n38917_ = ~new_n38915_ & ~new_n38916_;
  assign new_n38918_ = new_n10530_ & ~new_n38917_;
  assign new_n38919_ = ~new_n38650_ & new_n38918_;
  assign new_n38920_ = ~new_n38913_ & ~new_n38919_;
  assign new_n38921_ = ~\b[8]  & ~new_n38920_;
  assign new_n38922_ = ~new_n38423_ & ~new_n38651_;
  assign new_n38923_ = ~new_n38433_ & new_n38493_;
  assign new_n38924_ = ~new_n38489_ & new_n38923_;
  assign new_n38925_ = ~new_n38490_ & ~new_n38493_;
  assign new_n38926_ = ~new_n38924_ & ~new_n38925_;
  assign new_n38927_ = new_n10530_ & ~new_n38926_;
  assign new_n38928_ = ~new_n38650_ & new_n38927_;
  assign new_n38929_ = ~new_n38922_ & ~new_n38928_;
  assign new_n38930_ = ~\b[7]  & ~new_n38929_;
  assign new_n38931_ = ~new_n38432_ & ~new_n38651_;
  assign new_n38932_ = ~new_n38442_ & new_n38488_;
  assign new_n38933_ = ~new_n38484_ & new_n38932_;
  assign new_n38934_ = ~new_n38485_ & ~new_n38488_;
  assign new_n38935_ = ~new_n38933_ & ~new_n38934_;
  assign new_n38936_ = new_n10530_ & ~new_n38935_;
  assign new_n38937_ = ~new_n38650_ & new_n38936_;
  assign new_n38938_ = ~new_n38931_ & ~new_n38937_;
  assign new_n38939_ = ~\b[6]  & ~new_n38938_;
  assign new_n38940_ = ~new_n38441_ & ~new_n38651_;
  assign new_n38941_ = ~new_n38451_ & new_n38483_;
  assign new_n38942_ = ~new_n38479_ & new_n38941_;
  assign new_n38943_ = ~new_n38480_ & ~new_n38483_;
  assign new_n38944_ = ~new_n38942_ & ~new_n38943_;
  assign new_n38945_ = new_n10530_ & ~new_n38944_;
  assign new_n38946_ = ~new_n38650_ & new_n38945_;
  assign new_n38947_ = ~new_n38940_ & ~new_n38946_;
  assign new_n38948_ = ~\b[5]  & ~new_n38947_;
  assign new_n38949_ = ~new_n38450_ & ~new_n38651_;
  assign new_n38950_ = ~new_n38459_ & new_n38478_;
  assign new_n38951_ = ~new_n38474_ & new_n38950_;
  assign new_n38952_ = ~new_n38475_ & ~new_n38478_;
  assign new_n38953_ = ~new_n38951_ & ~new_n38952_;
  assign new_n38954_ = new_n10530_ & ~new_n38953_;
  assign new_n38955_ = ~new_n38650_ & new_n38954_;
  assign new_n38956_ = ~new_n38949_ & ~new_n38955_;
  assign new_n38957_ = ~\b[4]  & ~new_n38956_;
  assign new_n38958_ = ~new_n38458_ & ~new_n38651_;
  assign new_n38959_ = ~new_n38469_ & new_n38473_;
  assign new_n38960_ = ~new_n38468_ & new_n38959_;
  assign new_n38961_ = ~new_n38470_ & ~new_n38473_;
  assign new_n38962_ = ~new_n38960_ & ~new_n38961_;
  assign new_n38963_ = new_n10530_ & ~new_n38962_;
  assign new_n38964_ = ~new_n38650_ & new_n38963_;
  assign new_n38965_ = ~new_n38958_ & ~new_n38964_;
  assign new_n38966_ = ~\b[3]  & ~new_n38965_;
  assign new_n38967_ = ~new_n38463_ & ~new_n38651_;
  assign new_n38968_ = new_n10344_ & ~new_n38466_;
  assign new_n38969_ = ~new_n38464_ & new_n38968_;
  assign new_n38970_ = new_n10530_ & ~new_n38969_;
  assign new_n38971_ = ~new_n38468_ & new_n38970_;
  assign new_n38972_ = ~new_n38650_ & new_n38971_;
  assign new_n38973_ = ~new_n38967_ & ~new_n38972_;
  assign new_n38974_ = ~\b[2]  & ~new_n38973_;
  assign new_n38975_ = new_n10859_ & ~new_n38650_;
  assign new_n38976_ = \a[26]  & ~new_n38975_;
  assign new_n38977_ = new_n10865_ & ~new_n38650_;
  assign new_n38978_ = ~new_n38976_ & ~new_n38977_;
  assign new_n38979_ = \b[1]  & ~new_n38978_;
  assign new_n38980_ = ~\b[1]  & ~new_n38977_;
  assign new_n38981_ = ~new_n38976_ & new_n38980_;
  assign new_n38982_ = ~new_n38979_ & ~new_n38981_;
  assign new_n38983_ = ~new_n10872_ & ~new_n38982_;
  assign new_n38984_ = ~\b[1]  & ~new_n38978_;
  assign new_n38985_ = ~new_n38983_ & ~new_n38984_;
  assign new_n38986_ = \b[2]  & ~new_n38972_;
  assign new_n38987_ = ~new_n38967_ & new_n38986_;
  assign new_n38988_ = ~new_n38974_ & ~new_n38987_;
  assign new_n38989_ = ~new_n38985_ & new_n38988_;
  assign new_n38990_ = ~new_n38974_ & ~new_n38989_;
  assign new_n38991_ = \b[3]  & ~new_n38964_;
  assign new_n38992_ = ~new_n38958_ & new_n38991_;
  assign new_n38993_ = ~new_n38966_ & ~new_n38992_;
  assign new_n38994_ = ~new_n38990_ & new_n38993_;
  assign new_n38995_ = ~new_n38966_ & ~new_n38994_;
  assign new_n38996_ = \b[4]  & ~new_n38955_;
  assign new_n38997_ = ~new_n38949_ & new_n38996_;
  assign new_n38998_ = ~new_n38957_ & ~new_n38997_;
  assign new_n38999_ = ~new_n38995_ & new_n38998_;
  assign new_n39000_ = ~new_n38957_ & ~new_n38999_;
  assign new_n39001_ = \b[5]  & ~new_n38946_;
  assign new_n39002_ = ~new_n38940_ & new_n39001_;
  assign new_n39003_ = ~new_n38948_ & ~new_n39002_;
  assign new_n39004_ = ~new_n39000_ & new_n39003_;
  assign new_n39005_ = ~new_n38948_ & ~new_n39004_;
  assign new_n39006_ = \b[6]  & ~new_n38937_;
  assign new_n39007_ = ~new_n38931_ & new_n39006_;
  assign new_n39008_ = ~new_n38939_ & ~new_n39007_;
  assign new_n39009_ = ~new_n39005_ & new_n39008_;
  assign new_n39010_ = ~new_n38939_ & ~new_n39009_;
  assign new_n39011_ = \b[7]  & ~new_n38928_;
  assign new_n39012_ = ~new_n38922_ & new_n39011_;
  assign new_n39013_ = ~new_n38930_ & ~new_n39012_;
  assign new_n39014_ = ~new_n39010_ & new_n39013_;
  assign new_n39015_ = ~new_n38930_ & ~new_n39014_;
  assign new_n39016_ = \b[8]  & ~new_n38919_;
  assign new_n39017_ = ~new_n38913_ & new_n39016_;
  assign new_n39018_ = ~new_n38921_ & ~new_n39017_;
  assign new_n39019_ = ~new_n39015_ & new_n39018_;
  assign new_n39020_ = ~new_n38921_ & ~new_n39019_;
  assign new_n39021_ = \b[9]  & ~new_n38910_;
  assign new_n39022_ = ~new_n38904_ & new_n39021_;
  assign new_n39023_ = ~new_n38912_ & ~new_n39022_;
  assign new_n39024_ = ~new_n39020_ & new_n39023_;
  assign new_n39025_ = ~new_n38912_ & ~new_n39024_;
  assign new_n39026_ = \b[10]  & ~new_n38901_;
  assign new_n39027_ = ~new_n38895_ & new_n39026_;
  assign new_n39028_ = ~new_n38903_ & ~new_n39027_;
  assign new_n39029_ = ~new_n39025_ & new_n39028_;
  assign new_n39030_ = ~new_n38903_ & ~new_n39029_;
  assign new_n39031_ = \b[11]  & ~new_n38892_;
  assign new_n39032_ = ~new_n38886_ & new_n39031_;
  assign new_n39033_ = ~new_n38894_ & ~new_n39032_;
  assign new_n39034_ = ~new_n39030_ & new_n39033_;
  assign new_n39035_ = ~new_n38894_ & ~new_n39034_;
  assign new_n39036_ = \b[12]  & ~new_n38883_;
  assign new_n39037_ = ~new_n38877_ & new_n39036_;
  assign new_n39038_ = ~new_n38885_ & ~new_n39037_;
  assign new_n39039_ = ~new_n39035_ & new_n39038_;
  assign new_n39040_ = ~new_n38885_ & ~new_n39039_;
  assign new_n39041_ = \b[13]  & ~new_n38874_;
  assign new_n39042_ = ~new_n38868_ & new_n39041_;
  assign new_n39043_ = ~new_n38876_ & ~new_n39042_;
  assign new_n39044_ = ~new_n39040_ & new_n39043_;
  assign new_n39045_ = ~new_n38876_ & ~new_n39044_;
  assign new_n39046_ = \b[14]  & ~new_n38865_;
  assign new_n39047_ = ~new_n38859_ & new_n39046_;
  assign new_n39048_ = ~new_n38867_ & ~new_n39047_;
  assign new_n39049_ = ~new_n39045_ & new_n39048_;
  assign new_n39050_ = ~new_n38867_ & ~new_n39049_;
  assign new_n39051_ = \b[15]  & ~new_n38856_;
  assign new_n39052_ = ~new_n38850_ & new_n39051_;
  assign new_n39053_ = ~new_n38858_ & ~new_n39052_;
  assign new_n39054_ = ~new_n39050_ & new_n39053_;
  assign new_n39055_ = ~new_n38858_ & ~new_n39054_;
  assign new_n39056_ = \b[16]  & ~new_n38847_;
  assign new_n39057_ = ~new_n38841_ & new_n39056_;
  assign new_n39058_ = ~new_n38849_ & ~new_n39057_;
  assign new_n39059_ = ~new_n39055_ & new_n39058_;
  assign new_n39060_ = ~new_n38849_ & ~new_n39059_;
  assign new_n39061_ = \b[17]  & ~new_n38838_;
  assign new_n39062_ = ~new_n38832_ & new_n39061_;
  assign new_n39063_ = ~new_n38840_ & ~new_n39062_;
  assign new_n39064_ = ~new_n39060_ & new_n39063_;
  assign new_n39065_ = ~new_n38840_ & ~new_n39064_;
  assign new_n39066_ = \b[18]  & ~new_n38829_;
  assign new_n39067_ = ~new_n38823_ & new_n39066_;
  assign new_n39068_ = ~new_n38831_ & ~new_n39067_;
  assign new_n39069_ = ~new_n39065_ & new_n39068_;
  assign new_n39070_ = ~new_n38831_ & ~new_n39069_;
  assign new_n39071_ = \b[19]  & ~new_n38820_;
  assign new_n39072_ = ~new_n38814_ & new_n39071_;
  assign new_n39073_ = ~new_n38822_ & ~new_n39072_;
  assign new_n39074_ = ~new_n39070_ & new_n39073_;
  assign new_n39075_ = ~new_n38822_ & ~new_n39074_;
  assign new_n39076_ = \b[20]  & ~new_n38811_;
  assign new_n39077_ = ~new_n38805_ & new_n39076_;
  assign new_n39078_ = ~new_n38813_ & ~new_n39077_;
  assign new_n39079_ = ~new_n39075_ & new_n39078_;
  assign new_n39080_ = ~new_n38813_ & ~new_n39079_;
  assign new_n39081_ = \b[21]  & ~new_n38802_;
  assign new_n39082_ = ~new_n38796_ & new_n39081_;
  assign new_n39083_ = ~new_n38804_ & ~new_n39082_;
  assign new_n39084_ = ~new_n39080_ & new_n39083_;
  assign new_n39085_ = ~new_n38804_ & ~new_n39084_;
  assign new_n39086_ = \b[22]  & ~new_n38793_;
  assign new_n39087_ = ~new_n38787_ & new_n39086_;
  assign new_n39088_ = ~new_n38795_ & ~new_n39087_;
  assign new_n39089_ = ~new_n39085_ & new_n39088_;
  assign new_n39090_ = ~new_n38795_ & ~new_n39089_;
  assign new_n39091_ = \b[23]  & ~new_n38784_;
  assign new_n39092_ = ~new_n38778_ & new_n39091_;
  assign new_n39093_ = ~new_n38786_ & ~new_n39092_;
  assign new_n39094_ = ~new_n39090_ & new_n39093_;
  assign new_n39095_ = ~new_n38786_ & ~new_n39094_;
  assign new_n39096_ = \b[24]  & ~new_n38775_;
  assign new_n39097_ = ~new_n38769_ & new_n39096_;
  assign new_n39098_ = ~new_n38777_ & ~new_n39097_;
  assign new_n39099_ = ~new_n39095_ & new_n39098_;
  assign new_n39100_ = ~new_n38777_ & ~new_n39099_;
  assign new_n39101_ = \b[25]  & ~new_n38766_;
  assign new_n39102_ = ~new_n38760_ & new_n39101_;
  assign new_n39103_ = ~new_n38768_ & ~new_n39102_;
  assign new_n39104_ = ~new_n39100_ & new_n39103_;
  assign new_n39105_ = ~new_n38768_ & ~new_n39104_;
  assign new_n39106_ = \b[26]  & ~new_n38757_;
  assign new_n39107_ = ~new_n38751_ & new_n39106_;
  assign new_n39108_ = ~new_n38759_ & ~new_n39107_;
  assign new_n39109_ = ~new_n39105_ & new_n39108_;
  assign new_n39110_ = ~new_n38759_ & ~new_n39109_;
  assign new_n39111_ = \b[27]  & ~new_n38748_;
  assign new_n39112_ = ~new_n38742_ & new_n39111_;
  assign new_n39113_ = ~new_n38750_ & ~new_n39112_;
  assign new_n39114_ = ~new_n39110_ & new_n39113_;
  assign new_n39115_ = ~new_n38750_ & ~new_n39114_;
  assign new_n39116_ = \b[28]  & ~new_n38739_;
  assign new_n39117_ = ~new_n38733_ & new_n39116_;
  assign new_n39118_ = ~new_n38741_ & ~new_n39117_;
  assign new_n39119_ = ~new_n39115_ & new_n39118_;
  assign new_n39120_ = ~new_n38741_ & ~new_n39119_;
  assign new_n39121_ = \b[29]  & ~new_n38730_;
  assign new_n39122_ = ~new_n38724_ & new_n39121_;
  assign new_n39123_ = ~new_n38732_ & ~new_n39122_;
  assign new_n39124_ = ~new_n39120_ & new_n39123_;
  assign new_n39125_ = ~new_n38732_ & ~new_n39124_;
  assign new_n39126_ = \b[30]  & ~new_n38721_;
  assign new_n39127_ = ~new_n38715_ & new_n39126_;
  assign new_n39128_ = ~new_n38723_ & ~new_n39127_;
  assign new_n39129_ = ~new_n39125_ & new_n39128_;
  assign new_n39130_ = ~new_n38723_ & ~new_n39129_;
  assign new_n39131_ = \b[31]  & ~new_n38712_;
  assign new_n39132_ = ~new_n38706_ & new_n39131_;
  assign new_n39133_ = ~new_n38714_ & ~new_n39132_;
  assign new_n39134_ = ~new_n39130_ & new_n39133_;
  assign new_n39135_ = ~new_n38714_ & ~new_n39134_;
  assign new_n39136_ = \b[32]  & ~new_n38703_;
  assign new_n39137_ = ~new_n38697_ & new_n39136_;
  assign new_n39138_ = ~new_n38705_ & ~new_n39137_;
  assign new_n39139_ = ~new_n39135_ & new_n39138_;
  assign new_n39140_ = ~new_n38705_ & ~new_n39139_;
  assign new_n39141_ = \b[33]  & ~new_n38694_;
  assign new_n39142_ = ~new_n38688_ & new_n39141_;
  assign new_n39143_ = ~new_n38696_ & ~new_n39142_;
  assign new_n39144_ = ~new_n39140_ & new_n39143_;
  assign new_n39145_ = ~new_n38696_ & ~new_n39144_;
  assign new_n39146_ = \b[34]  & ~new_n38685_;
  assign new_n39147_ = ~new_n38679_ & new_n39146_;
  assign new_n39148_ = ~new_n38687_ & ~new_n39147_;
  assign new_n39149_ = ~new_n39145_ & new_n39148_;
  assign new_n39150_ = ~new_n38687_ & ~new_n39149_;
  assign new_n39151_ = \b[35]  & ~new_n38676_;
  assign new_n39152_ = ~new_n38670_ & new_n39151_;
  assign new_n39153_ = ~new_n38678_ & ~new_n39152_;
  assign new_n39154_ = ~new_n39150_ & new_n39153_;
  assign new_n39155_ = ~new_n38678_ & ~new_n39154_;
  assign new_n39156_ = \b[36]  & ~new_n38667_;
  assign new_n39157_ = ~new_n38661_ & new_n39156_;
  assign new_n39158_ = ~new_n38669_ & ~new_n39157_;
  assign new_n39159_ = ~new_n39155_ & new_n39158_;
  assign new_n39160_ = ~new_n38669_ & ~new_n39159_;
  assign new_n39161_ = \b[37]  & ~new_n38658_;
  assign new_n39162_ = ~new_n38652_ & new_n39161_;
  assign new_n39163_ = ~new_n38660_ & ~new_n39162_;
  assign new_n39164_ = ~new_n39160_ & new_n39163_;
  assign new_n39165_ = ~new_n38660_ & ~new_n39164_;
  assign new_n39166_ = ~new_n38152_ & ~new_n38651_;
  assign new_n39167_ = ~new_n38154_ & new_n38648_;
  assign new_n39168_ = ~new_n38644_ & new_n39167_;
  assign new_n39169_ = ~new_n38645_ & ~new_n38648_;
  assign new_n39170_ = ~new_n39168_ & ~new_n39169_;
  assign new_n39171_ = new_n38651_ & ~new_n39170_;
  assign new_n39172_ = ~new_n39166_ & ~new_n39171_;
  assign new_n39173_ = ~\b[38]  & ~new_n39172_;
  assign new_n39174_ = \b[38]  & ~new_n39166_;
  assign new_n39175_ = ~new_n39171_ & new_n39174_;
  assign new_n39176_ = new_n11068_ & ~new_n39175_;
  assign new_n39177_ = ~new_n39173_ & new_n39176_;
  assign new_n39178_ = ~new_n39165_ & new_n39177_;
  assign new_n39179_ = new_n10530_ & ~new_n39172_;
  assign new_n39180_ = ~new_n39178_ & ~new_n39179_;
  assign new_n39181_ = ~new_n38669_ & new_n39163_;
  assign new_n39182_ = ~new_n39159_ & new_n39181_;
  assign new_n39183_ = ~new_n39160_ & ~new_n39163_;
  assign new_n39184_ = ~new_n39182_ & ~new_n39183_;
  assign new_n39185_ = ~new_n39180_ & ~new_n39184_;
  assign new_n39186_ = ~new_n38659_ & ~new_n39179_;
  assign new_n39187_ = ~new_n39178_ & new_n39186_;
  assign new_n39188_ = ~new_n39185_ & ~new_n39187_;
  assign new_n39189_ = ~new_n38660_ & ~new_n39175_;
  assign new_n39190_ = ~new_n39173_ & new_n39189_;
  assign new_n39191_ = ~new_n39164_ & new_n39190_;
  assign new_n39192_ = ~new_n39173_ & ~new_n39175_;
  assign new_n39193_ = ~new_n39165_ & ~new_n39192_;
  assign new_n39194_ = ~new_n39191_ & ~new_n39193_;
  assign new_n39195_ = ~new_n39180_ & ~new_n39194_;
  assign new_n39196_ = ~new_n39172_ & ~new_n39179_;
  assign new_n39197_ = ~new_n39178_ & new_n39196_;
  assign new_n39198_ = ~new_n39195_ & ~new_n39197_;
  assign new_n39199_ = ~\b[39]  & ~new_n39198_;
  assign new_n39200_ = ~\b[38]  & ~new_n39188_;
  assign new_n39201_ = ~new_n38678_ & new_n39158_;
  assign new_n39202_ = ~new_n39154_ & new_n39201_;
  assign new_n39203_ = ~new_n39155_ & ~new_n39158_;
  assign new_n39204_ = ~new_n39202_ & ~new_n39203_;
  assign new_n39205_ = ~new_n39180_ & ~new_n39204_;
  assign new_n39206_ = ~new_n38668_ & ~new_n39179_;
  assign new_n39207_ = ~new_n39178_ & new_n39206_;
  assign new_n39208_ = ~new_n39205_ & ~new_n39207_;
  assign new_n39209_ = ~\b[37]  & ~new_n39208_;
  assign new_n39210_ = ~new_n38687_ & new_n39153_;
  assign new_n39211_ = ~new_n39149_ & new_n39210_;
  assign new_n39212_ = ~new_n39150_ & ~new_n39153_;
  assign new_n39213_ = ~new_n39211_ & ~new_n39212_;
  assign new_n39214_ = ~new_n39180_ & ~new_n39213_;
  assign new_n39215_ = ~new_n38677_ & ~new_n39179_;
  assign new_n39216_ = ~new_n39178_ & new_n39215_;
  assign new_n39217_ = ~new_n39214_ & ~new_n39216_;
  assign new_n39218_ = ~\b[36]  & ~new_n39217_;
  assign new_n39219_ = ~new_n38696_ & new_n39148_;
  assign new_n39220_ = ~new_n39144_ & new_n39219_;
  assign new_n39221_ = ~new_n39145_ & ~new_n39148_;
  assign new_n39222_ = ~new_n39220_ & ~new_n39221_;
  assign new_n39223_ = ~new_n39180_ & ~new_n39222_;
  assign new_n39224_ = ~new_n38686_ & ~new_n39179_;
  assign new_n39225_ = ~new_n39178_ & new_n39224_;
  assign new_n39226_ = ~new_n39223_ & ~new_n39225_;
  assign new_n39227_ = ~\b[35]  & ~new_n39226_;
  assign new_n39228_ = ~new_n38705_ & new_n39143_;
  assign new_n39229_ = ~new_n39139_ & new_n39228_;
  assign new_n39230_ = ~new_n39140_ & ~new_n39143_;
  assign new_n39231_ = ~new_n39229_ & ~new_n39230_;
  assign new_n39232_ = ~new_n39180_ & ~new_n39231_;
  assign new_n39233_ = ~new_n38695_ & ~new_n39179_;
  assign new_n39234_ = ~new_n39178_ & new_n39233_;
  assign new_n39235_ = ~new_n39232_ & ~new_n39234_;
  assign new_n39236_ = ~\b[34]  & ~new_n39235_;
  assign new_n39237_ = ~new_n38714_ & new_n39138_;
  assign new_n39238_ = ~new_n39134_ & new_n39237_;
  assign new_n39239_ = ~new_n39135_ & ~new_n39138_;
  assign new_n39240_ = ~new_n39238_ & ~new_n39239_;
  assign new_n39241_ = ~new_n39180_ & ~new_n39240_;
  assign new_n39242_ = ~new_n38704_ & ~new_n39179_;
  assign new_n39243_ = ~new_n39178_ & new_n39242_;
  assign new_n39244_ = ~new_n39241_ & ~new_n39243_;
  assign new_n39245_ = ~\b[33]  & ~new_n39244_;
  assign new_n39246_ = ~new_n38723_ & new_n39133_;
  assign new_n39247_ = ~new_n39129_ & new_n39246_;
  assign new_n39248_ = ~new_n39130_ & ~new_n39133_;
  assign new_n39249_ = ~new_n39247_ & ~new_n39248_;
  assign new_n39250_ = ~new_n39180_ & ~new_n39249_;
  assign new_n39251_ = ~new_n38713_ & ~new_n39179_;
  assign new_n39252_ = ~new_n39178_ & new_n39251_;
  assign new_n39253_ = ~new_n39250_ & ~new_n39252_;
  assign new_n39254_ = ~\b[32]  & ~new_n39253_;
  assign new_n39255_ = ~new_n38732_ & new_n39128_;
  assign new_n39256_ = ~new_n39124_ & new_n39255_;
  assign new_n39257_ = ~new_n39125_ & ~new_n39128_;
  assign new_n39258_ = ~new_n39256_ & ~new_n39257_;
  assign new_n39259_ = ~new_n39180_ & ~new_n39258_;
  assign new_n39260_ = ~new_n38722_ & ~new_n39179_;
  assign new_n39261_ = ~new_n39178_ & new_n39260_;
  assign new_n39262_ = ~new_n39259_ & ~new_n39261_;
  assign new_n39263_ = ~\b[31]  & ~new_n39262_;
  assign new_n39264_ = ~new_n38741_ & new_n39123_;
  assign new_n39265_ = ~new_n39119_ & new_n39264_;
  assign new_n39266_ = ~new_n39120_ & ~new_n39123_;
  assign new_n39267_ = ~new_n39265_ & ~new_n39266_;
  assign new_n39268_ = ~new_n39180_ & ~new_n39267_;
  assign new_n39269_ = ~new_n38731_ & ~new_n39179_;
  assign new_n39270_ = ~new_n39178_ & new_n39269_;
  assign new_n39271_ = ~new_n39268_ & ~new_n39270_;
  assign new_n39272_ = ~\b[30]  & ~new_n39271_;
  assign new_n39273_ = ~new_n38750_ & new_n39118_;
  assign new_n39274_ = ~new_n39114_ & new_n39273_;
  assign new_n39275_ = ~new_n39115_ & ~new_n39118_;
  assign new_n39276_ = ~new_n39274_ & ~new_n39275_;
  assign new_n39277_ = ~new_n39180_ & ~new_n39276_;
  assign new_n39278_ = ~new_n38740_ & ~new_n39179_;
  assign new_n39279_ = ~new_n39178_ & new_n39278_;
  assign new_n39280_ = ~new_n39277_ & ~new_n39279_;
  assign new_n39281_ = ~\b[29]  & ~new_n39280_;
  assign new_n39282_ = ~new_n38759_ & new_n39113_;
  assign new_n39283_ = ~new_n39109_ & new_n39282_;
  assign new_n39284_ = ~new_n39110_ & ~new_n39113_;
  assign new_n39285_ = ~new_n39283_ & ~new_n39284_;
  assign new_n39286_ = ~new_n39180_ & ~new_n39285_;
  assign new_n39287_ = ~new_n38749_ & ~new_n39179_;
  assign new_n39288_ = ~new_n39178_ & new_n39287_;
  assign new_n39289_ = ~new_n39286_ & ~new_n39288_;
  assign new_n39290_ = ~\b[28]  & ~new_n39289_;
  assign new_n39291_ = ~new_n38768_ & new_n39108_;
  assign new_n39292_ = ~new_n39104_ & new_n39291_;
  assign new_n39293_ = ~new_n39105_ & ~new_n39108_;
  assign new_n39294_ = ~new_n39292_ & ~new_n39293_;
  assign new_n39295_ = ~new_n39180_ & ~new_n39294_;
  assign new_n39296_ = ~new_n38758_ & ~new_n39179_;
  assign new_n39297_ = ~new_n39178_ & new_n39296_;
  assign new_n39298_ = ~new_n39295_ & ~new_n39297_;
  assign new_n39299_ = ~\b[27]  & ~new_n39298_;
  assign new_n39300_ = ~new_n38777_ & new_n39103_;
  assign new_n39301_ = ~new_n39099_ & new_n39300_;
  assign new_n39302_ = ~new_n39100_ & ~new_n39103_;
  assign new_n39303_ = ~new_n39301_ & ~new_n39302_;
  assign new_n39304_ = ~new_n39180_ & ~new_n39303_;
  assign new_n39305_ = ~new_n38767_ & ~new_n39179_;
  assign new_n39306_ = ~new_n39178_ & new_n39305_;
  assign new_n39307_ = ~new_n39304_ & ~new_n39306_;
  assign new_n39308_ = ~\b[26]  & ~new_n39307_;
  assign new_n39309_ = ~new_n38786_ & new_n39098_;
  assign new_n39310_ = ~new_n39094_ & new_n39309_;
  assign new_n39311_ = ~new_n39095_ & ~new_n39098_;
  assign new_n39312_ = ~new_n39310_ & ~new_n39311_;
  assign new_n39313_ = ~new_n39180_ & ~new_n39312_;
  assign new_n39314_ = ~new_n38776_ & ~new_n39179_;
  assign new_n39315_ = ~new_n39178_ & new_n39314_;
  assign new_n39316_ = ~new_n39313_ & ~new_n39315_;
  assign new_n39317_ = ~\b[25]  & ~new_n39316_;
  assign new_n39318_ = ~new_n38795_ & new_n39093_;
  assign new_n39319_ = ~new_n39089_ & new_n39318_;
  assign new_n39320_ = ~new_n39090_ & ~new_n39093_;
  assign new_n39321_ = ~new_n39319_ & ~new_n39320_;
  assign new_n39322_ = ~new_n39180_ & ~new_n39321_;
  assign new_n39323_ = ~new_n38785_ & ~new_n39179_;
  assign new_n39324_ = ~new_n39178_ & new_n39323_;
  assign new_n39325_ = ~new_n39322_ & ~new_n39324_;
  assign new_n39326_ = ~\b[24]  & ~new_n39325_;
  assign new_n39327_ = ~new_n38804_ & new_n39088_;
  assign new_n39328_ = ~new_n39084_ & new_n39327_;
  assign new_n39329_ = ~new_n39085_ & ~new_n39088_;
  assign new_n39330_ = ~new_n39328_ & ~new_n39329_;
  assign new_n39331_ = ~new_n39180_ & ~new_n39330_;
  assign new_n39332_ = ~new_n38794_ & ~new_n39179_;
  assign new_n39333_ = ~new_n39178_ & new_n39332_;
  assign new_n39334_ = ~new_n39331_ & ~new_n39333_;
  assign new_n39335_ = ~\b[23]  & ~new_n39334_;
  assign new_n39336_ = ~new_n38813_ & new_n39083_;
  assign new_n39337_ = ~new_n39079_ & new_n39336_;
  assign new_n39338_ = ~new_n39080_ & ~new_n39083_;
  assign new_n39339_ = ~new_n39337_ & ~new_n39338_;
  assign new_n39340_ = ~new_n39180_ & ~new_n39339_;
  assign new_n39341_ = ~new_n38803_ & ~new_n39179_;
  assign new_n39342_ = ~new_n39178_ & new_n39341_;
  assign new_n39343_ = ~new_n39340_ & ~new_n39342_;
  assign new_n39344_ = ~\b[22]  & ~new_n39343_;
  assign new_n39345_ = ~new_n38822_ & new_n39078_;
  assign new_n39346_ = ~new_n39074_ & new_n39345_;
  assign new_n39347_ = ~new_n39075_ & ~new_n39078_;
  assign new_n39348_ = ~new_n39346_ & ~new_n39347_;
  assign new_n39349_ = ~new_n39180_ & ~new_n39348_;
  assign new_n39350_ = ~new_n38812_ & ~new_n39179_;
  assign new_n39351_ = ~new_n39178_ & new_n39350_;
  assign new_n39352_ = ~new_n39349_ & ~new_n39351_;
  assign new_n39353_ = ~\b[21]  & ~new_n39352_;
  assign new_n39354_ = ~new_n38831_ & new_n39073_;
  assign new_n39355_ = ~new_n39069_ & new_n39354_;
  assign new_n39356_ = ~new_n39070_ & ~new_n39073_;
  assign new_n39357_ = ~new_n39355_ & ~new_n39356_;
  assign new_n39358_ = ~new_n39180_ & ~new_n39357_;
  assign new_n39359_ = ~new_n38821_ & ~new_n39179_;
  assign new_n39360_ = ~new_n39178_ & new_n39359_;
  assign new_n39361_ = ~new_n39358_ & ~new_n39360_;
  assign new_n39362_ = ~\b[20]  & ~new_n39361_;
  assign new_n39363_ = ~new_n38840_ & new_n39068_;
  assign new_n39364_ = ~new_n39064_ & new_n39363_;
  assign new_n39365_ = ~new_n39065_ & ~new_n39068_;
  assign new_n39366_ = ~new_n39364_ & ~new_n39365_;
  assign new_n39367_ = ~new_n39180_ & ~new_n39366_;
  assign new_n39368_ = ~new_n38830_ & ~new_n39179_;
  assign new_n39369_ = ~new_n39178_ & new_n39368_;
  assign new_n39370_ = ~new_n39367_ & ~new_n39369_;
  assign new_n39371_ = ~\b[19]  & ~new_n39370_;
  assign new_n39372_ = ~new_n38849_ & new_n39063_;
  assign new_n39373_ = ~new_n39059_ & new_n39372_;
  assign new_n39374_ = ~new_n39060_ & ~new_n39063_;
  assign new_n39375_ = ~new_n39373_ & ~new_n39374_;
  assign new_n39376_ = ~new_n39180_ & ~new_n39375_;
  assign new_n39377_ = ~new_n38839_ & ~new_n39179_;
  assign new_n39378_ = ~new_n39178_ & new_n39377_;
  assign new_n39379_ = ~new_n39376_ & ~new_n39378_;
  assign new_n39380_ = ~\b[18]  & ~new_n39379_;
  assign new_n39381_ = ~new_n38858_ & new_n39058_;
  assign new_n39382_ = ~new_n39054_ & new_n39381_;
  assign new_n39383_ = ~new_n39055_ & ~new_n39058_;
  assign new_n39384_ = ~new_n39382_ & ~new_n39383_;
  assign new_n39385_ = ~new_n39180_ & ~new_n39384_;
  assign new_n39386_ = ~new_n38848_ & ~new_n39179_;
  assign new_n39387_ = ~new_n39178_ & new_n39386_;
  assign new_n39388_ = ~new_n39385_ & ~new_n39387_;
  assign new_n39389_ = ~\b[17]  & ~new_n39388_;
  assign new_n39390_ = ~new_n38867_ & new_n39053_;
  assign new_n39391_ = ~new_n39049_ & new_n39390_;
  assign new_n39392_ = ~new_n39050_ & ~new_n39053_;
  assign new_n39393_ = ~new_n39391_ & ~new_n39392_;
  assign new_n39394_ = ~new_n39180_ & ~new_n39393_;
  assign new_n39395_ = ~new_n38857_ & ~new_n39179_;
  assign new_n39396_ = ~new_n39178_ & new_n39395_;
  assign new_n39397_ = ~new_n39394_ & ~new_n39396_;
  assign new_n39398_ = ~\b[16]  & ~new_n39397_;
  assign new_n39399_ = ~new_n38876_ & new_n39048_;
  assign new_n39400_ = ~new_n39044_ & new_n39399_;
  assign new_n39401_ = ~new_n39045_ & ~new_n39048_;
  assign new_n39402_ = ~new_n39400_ & ~new_n39401_;
  assign new_n39403_ = ~new_n39180_ & ~new_n39402_;
  assign new_n39404_ = ~new_n38866_ & ~new_n39179_;
  assign new_n39405_ = ~new_n39178_ & new_n39404_;
  assign new_n39406_ = ~new_n39403_ & ~new_n39405_;
  assign new_n39407_ = ~\b[15]  & ~new_n39406_;
  assign new_n39408_ = ~new_n38885_ & new_n39043_;
  assign new_n39409_ = ~new_n39039_ & new_n39408_;
  assign new_n39410_ = ~new_n39040_ & ~new_n39043_;
  assign new_n39411_ = ~new_n39409_ & ~new_n39410_;
  assign new_n39412_ = ~new_n39180_ & ~new_n39411_;
  assign new_n39413_ = ~new_n38875_ & ~new_n39179_;
  assign new_n39414_ = ~new_n39178_ & new_n39413_;
  assign new_n39415_ = ~new_n39412_ & ~new_n39414_;
  assign new_n39416_ = ~\b[14]  & ~new_n39415_;
  assign new_n39417_ = ~new_n38894_ & new_n39038_;
  assign new_n39418_ = ~new_n39034_ & new_n39417_;
  assign new_n39419_ = ~new_n39035_ & ~new_n39038_;
  assign new_n39420_ = ~new_n39418_ & ~new_n39419_;
  assign new_n39421_ = ~new_n39180_ & ~new_n39420_;
  assign new_n39422_ = ~new_n38884_ & ~new_n39179_;
  assign new_n39423_ = ~new_n39178_ & new_n39422_;
  assign new_n39424_ = ~new_n39421_ & ~new_n39423_;
  assign new_n39425_ = ~\b[13]  & ~new_n39424_;
  assign new_n39426_ = ~new_n38903_ & new_n39033_;
  assign new_n39427_ = ~new_n39029_ & new_n39426_;
  assign new_n39428_ = ~new_n39030_ & ~new_n39033_;
  assign new_n39429_ = ~new_n39427_ & ~new_n39428_;
  assign new_n39430_ = ~new_n39180_ & ~new_n39429_;
  assign new_n39431_ = ~new_n38893_ & ~new_n39179_;
  assign new_n39432_ = ~new_n39178_ & new_n39431_;
  assign new_n39433_ = ~new_n39430_ & ~new_n39432_;
  assign new_n39434_ = ~\b[12]  & ~new_n39433_;
  assign new_n39435_ = ~new_n38912_ & new_n39028_;
  assign new_n39436_ = ~new_n39024_ & new_n39435_;
  assign new_n39437_ = ~new_n39025_ & ~new_n39028_;
  assign new_n39438_ = ~new_n39436_ & ~new_n39437_;
  assign new_n39439_ = ~new_n39180_ & ~new_n39438_;
  assign new_n39440_ = ~new_n38902_ & ~new_n39179_;
  assign new_n39441_ = ~new_n39178_ & new_n39440_;
  assign new_n39442_ = ~new_n39439_ & ~new_n39441_;
  assign new_n39443_ = ~\b[11]  & ~new_n39442_;
  assign new_n39444_ = ~new_n38921_ & new_n39023_;
  assign new_n39445_ = ~new_n39019_ & new_n39444_;
  assign new_n39446_ = ~new_n39020_ & ~new_n39023_;
  assign new_n39447_ = ~new_n39445_ & ~new_n39446_;
  assign new_n39448_ = ~new_n39180_ & ~new_n39447_;
  assign new_n39449_ = ~new_n38911_ & ~new_n39179_;
  assign new_n39450_ = ~new_n39178_ & new_n39449_;
  assign new_n39451_ = ~new_n39448_ & ~new_n39450_;
  assign new_n39452_ = ~\b[10]  & ~new_n39451_;
  assign new_n39453_ = ~new_n38930_ & new_n39018_;
  assign new_n39454_ = ~new_n39014_ & new_n39453_;
  assign new_n39455_ = ~new_n39015_ & ~new_n39018_;
  assign new_n39456_ = ~new_n39454_ & ~new_n39455_;
  assign new_n39457_ = ~new_n39180_ & ~new_n39456_;
  assign new_n39458_ = ~new_n38920_ & ~new_n39179_;
  assign new_n39459_ = ~new_n39178_ & new_n39458_;
  assign new_n39460_ = ~new_n39457_ & ~new_n39459_;
  assign new_n39461_ = ~\b[9]  & ~new_n39460_;
  assign new_n39462_ = ~new_n38939_ & new_n39013_;
  assign new_n39463_ = ~new_n39009_ & new_n39462_;
  assign new_n39464_ = ~new_n39010_ & ~new_n39013_;
  assign new_n39465_ = ~new_n39463_ & ~new_n39464_;
  assign new_n39466_ = ~new_n39180_ & ~new_n39465_;
  assign new_n39467_ = ~new_n38929_ & ~new_n39179_;
  assign new_n39468_ = ~new_n39178_ & new_n39467_;
  assign new_n39469_ = ~new_n39466_ & ~new_n39468_;
  assign new_n39470_ = ~\b[8]  & ~new_n39469_;
  assign new_n39471_ = ~new_n38948_ & new_n39008_;
  assign new_n39472_ = ~new_n39004_ & new_n39471_;
  assign new_n39473_ = ~new_n39005_ & ~new_n39008_;
  assign new_n39474_ = ~new_n39472_ & ~new_n39473_;
  assign new_n39475_ = ~new_n39180_ & ~new_n39474_;
  assign new_n39476_ = ~new_n38938_ & ~new_n39179_;
  assign new_n39477_ = ~new_n39178_ & new_n39476_;
  assign new_n39478_ = ~new_n39475_ & ~new_n39477_;
  assign new_n39479_ = ~\b[7]  & ~new_n39478_;
  assign new_n39480_ = ~new_n38957_ & new_n39003_;
  assign new_n39481_ = ~new_n38999_ & new_n39480_;
  assign new_n39482_ = ~new_n39000_ & ~new_n39003_;
  assign new_n39483_ = ~new_n39481_ & ~new_n39482_;
  assign new_n39484_ = ~new_n39180_ & ~new_n39483_;
  assign new_n39485_ = ~new_n38947_ & ~new_n39179_;
  assign new_n39486_ = ~new_n39178_ & new_n39485_;
  assign new_n39487_ = ~new_n39484_ & ~new_n39486_;
  assign new_n39488_ = ~\b[6]  & ~new_n39487_;
  assign new_n39489_ = ~new_n38966_ & new_n38998_;
  assign new_n39490_ = ~new_n38994_ & new_n39489_;
  assign new_n39491_ = ~new_n38995_ & ~new_n38998_;
  assign new_n39492_ = ~new_n39490_ & ~new_n39491_;
  assign new_n39493_ = ~new_n39180_ & ~new_n39492_;
  assign new_n39494_ = ~new_n38956_ & ~new_n39179_;
  assign new_n39495_ = ~new_n39178_ & new_n39494_;
  assign new_n39496_ = ~new_n39493_ & ~new_n39495_;
  assign new_n39497_ = ~\b[5]  & ~new_n39496_;
  assign new_n39498_ = ~new_n38974_ & new_n38993_;
  assign new_n39499_ = ~new_n38989_ & new_n39498_;
  assign new_n39500_ = ~new_n38990_ & ~new_n38993_;
  assign new_n39501_ = ~new_n39499_ & ~new_n39500_;
  assign new_n39502_ = ~new_n39180_ & ~new_n39501_;
  assign new_n39503_ = ~new_n38965_ & ~new_n39179_;
  assign new_n39504_ = ~new_n39178_ & new_n39503_;
  assign new_n39505_ = ~new_n39502_ & ~new_n39504_;
  assign new_n39506_ = ~\b[4]  & ~new_n39505_;
  assign new_n39507_ = ~new_n38984_ & new_n38988_;
  assign new_n39508_ = ~new_n38983_ & new_n39507_;
  assign new_n39509_ = ~new_n38985_ & ~new_n38988_;
  assign new_n39510_ = ~new_n39508_ & ~new_n39509_;
  assign new_n39511_ = ~new_n39180_ & ~new_n39510_;
  assign new_n39512_ = ~new_n38973_ & ~new_n39179_;
  assign new_n39513_ = ~new_n39178_ & new_n39512_;
  assign new_n39514_ = ~new_n39511_ & ~new_n39513_;
  assign new_n39515_ = ~\b[3]  & ~new_n39514_;
  assign new_n39516_ = new_n10872_ & ~new_n38981_;
  assign new_n39517_ = ~new_n38979_ & new_n39516_;
  assign new_n39518_ = ~new_n38983_ & ~new_n39517_;
  assign new_n39519_ = ~new_n39180_ & new_n39518_;
  assign new_n39520_ = ~new_n38978_ & ~new_n39179_;
  assign new_n39521_ = ~new_n39178_ & new_n39520_;
  assign new_n39522_ = ~new_n39519_ & ~new_n39521_;
  assign new_n39523_ = ~\b[2]  & ~new_n39522_;
  assign new_n39524_ = \b[0]  & ~new_n39180_;
  assign new_n39525_ = \a[25]  & ~new_n39524_;
  assign new_n39526_ = new_n10872_ & ~new_n39180_;
  assign new_n39527_ = ~new_n39525_ & ~new_n39526_;
  assign new_n39528_ = \b[1]  & ~new_n39527_;
  assign new_n39529_ = ~\b[1]  & ~new_n39526_;
  assign new_n39530_ = ~new_n39525_ & new_n39529_;
  assign new_n39531_ = ~new_n39528_ & ~new_n39530_;
  assign new_n39532_ = ~new_n11425_ & ~new_n39531_;
  assign new_n39533_ = ~\b[1]  & ~new_n39527_;
  assign new_n39534_ = ~new_n39532_ & ~new_n39533_;
  assign new_n39535_ = \b[2]  & ~new_n39521_;
  assign new_n39536_ = ~new_n39519_ & new_n39535_;
  assign new_n39537_ = ~new_n39523_ & ~new_n39536_;
  assign new_n39538_ = ~new_n39534_ & new_n39537_;
  assign new_n39539_ = ~new_n39523_ & ~new_n39538_;
  assign new_n39540_ = \b[3]  & ~new_n39513_;
  assign new_n39541_ = ~new_n39511_ & new_n39540_;
  assign new_n39542_ = ~new_n39515_ & ~new_n39541_;
  assign new_n39543_ = ~new_n39539_ & new_n39542_;
  assign new_n39544_ = ~new_n39515_ & ~new_n39543_;
  assign new_n39545_ = \b[4]  & ~new_n39504_;
  assign new_n39546_ = ~new_n39502_ & new_n39545_;
  assign new_n39547_ = ~new_n39506_ & ~new_n39546_;
  assign new_n39548_ = ~new_n39544_ & new_n39547_;
  assign new_n39549_ = ~new_n39506_ & ~new_n39548_;
  assign new_n39550_ = \b[5]  & ~new_n39495_;
  assign new_n39551_ = ~new_n39493_ & new_n39550_;
  assign new_n39552_ = ~new_n39497_ & ~new_n39551_;
  assign new_n39553_ = ~new_n39549_ & new_n39552_;
  assign new_n39554_ = ~new_n39497_ & ~new_n39553_;
  assign new_n39555_ = \b[6]  & ~new_n39486_;
  assign new_n39556_ = ~new_n39484_ & new_n39555_;
  assign new_n39557_ = ~new_n39488_ & ~new_n39556_;
  assign new_n39558_ = ~new_n39554_ & new_n39557_;
  assign new_n39559_ = ~new_n39488_ & ~new_n39558_;
  assign new_n39560_ = \b[7]  & ~new_n39477_;
  assign new_n39561_ = ~new_n39475_ & new_n39560_;
  assign new_n39562_ = ~new_n39479_ & ~new_n39561_;
  assign new_n39563_ = ~new_n39559_ & new_n39562_;
  assign new_n39564_ = ~new_n39479_ & ~new_n39563_;
  assign new_n39565_ = \b[8]  & ~new_n39468_;
  assign new_n39566_ = ~new_n39466_ & new_n39565_;
  assign new_n39567_ = ~new_n39470_ & ~new_n39566_;
  assign new_n39568_ = ~new_n39564_ & new_n39567_;
  assign new_n39569_ = ~new_n39470_ & ~new_n39568_;
  assign new_n39570_ = \b[9]  & ~new_n39459_;
  assign new_n39571_ = ~new_n39457_ & new_n39570_;
  assign new_n39572_ = ~new_n39461_ & ~new_n39571_;
  assign new_n39573_ = ~new_n39569_ & new_n39572_;
  assign new_n39574_ = ~new_n39461_ & ~new_n39573_;
  assign new_n39575_ = \b[10]  & ~new_n39450_;
  assign new_n39576_ = ~new_n39448_ & new_n39575_;
  assign new_n39577_ = ~new_n39452_ & ~new_n39576_;
  assign new_n39578_ = ~new_n39574_ & new_n39577_;
  assign new_n39579_ = ~new_n39452_ & ~new_n39578_;
  assign new_n39580_ = \b[11]  & ~new_n39441_;
  assign new_n39581_ = ~new_n39439_ & new_n39580_;
  assign new_n39582_ = ~new_n39443_ & ~new_n39581_;
  assign new_n39583_ = ~new_n39579_ & new_n39582_;
  assign new_n39584_ = ~new_n39443_ & ~new_n39583_;
  assign new_n39585_ = \b[12]  & ~new_n39432_;
  assign new_n39586_ = ~new_n39430_ & new_n39585_;
  assign new_n39587_ = ~new_n39434_ & ~new_n39586_;
  assign new_n39588_ = ~new_n39584_ & new_n39587_;
  assign new_n39589_ = ~new_n39434_ & ~new_n39588_;
  assign new_n39590_ = \b[13]  & ~new_n39423_;
  assign new_n39591_ = ~new_n39421_ & new_n39590_;
  assign new_n39592_ = ~new_n39425_ & ~new_n39591_;
  assign new_n39593_ = ~new_n39589_ & new_n39592_;
  assign new_n39594_ = ~new_n39425_ & ~new_n39593_;
  assign new_n39595_ = \b[14]  & ~new_n39414_;
  assign new_n39596_ = ~new_n39412_ & new_n39595_;
  assign new_n39597_ = ~new_n39416_ & ~new_n39596_;
  assign new_n39598_ = ~new_n39594_ & new_n39597_;
  assign new_n39599_ = ~new_n39416_ & ~new_n39598_;
  assign new_n39600_ = \b[15]  & ~new_n39405_;
  assign new_n39601_ = ~new_n39403_ & new_n39600_;
  assign new_n39602_ = ~new_n39407_ & ~new_n39601_;
  assign new_n39603_ = ~new_n39599_ & new_n39602_;
  assign new_n39604_ = ~new_n39407_ & ~new_n39603_;
  assign new_n39605_ = \b[16]  & ~new_n39396_;
  assign new_n39606_ = ~new_n39394_ & new_n39605_;
  assign new_n39607_ = ~new_n39398_ & ~new_n39606_;
  assign new_n39608_ = ~new_n39604_ & new_n39607_;
  assign new_n39609_ = ~new_n39398_ & ~new_n39608_;
  assign new_n39610_ = \b[17]  & ~new_n39387_;
  assign new_n39611_ = ~new_n39385_ & new_n39610_;
  assign new_n39612_ = ~new_n39389_ & ~new_n39611_;
  assign new_n39613_ = ~new_n39609_ & new_n39612_;
  assign new_n39614_ = ~new_n39389_ & ~new_n39613_;
  assign new_n39615_ = \b[18]  & ~new_n39378_;
  assign new_n39616_ = ~new_n39376_ & new_n39615_;
  assign new_n39617_ = ~new_n39380_ & ~new_n39616_;
  assign new_n39618_ = ~new_n39614_ & new_n39617_;
  assign new_n39619_ = ~new_n39380_ & ~new_n39618_;
  assign new_n39620_ = \b[19]  & ~new_n39369_;
  assign new_n39621_ = ~new_n39367_ & new_n39620_;
  assign new_n39622_ = ~new_n39371_ & ~new_n39621_;
  assign new_n39623_ = ~new_n39619_ & new_n39622_;
  assign new_n39624_ = ~new_n39371_ & ~new_n39623_;
  assign new_n39625_ = \b[20]  & ~new_n39360_;
  assign new_n39626_ = ~new_n39358_ & new_n39625_;
  assign new_n39627_ = ~new_n39362_ & ~new_n39626_;
  assign new_n39628_ = ~new_n39624_ & new_n39627_;
  assign new_n39629_ = ~new_n39362_ & ~new_n39628_;
  assign new_n39630_ = \b[21]  & ~new_n39351_;
  assign new_n39631_ = ~new_n39349_ & new_n39630_;
  assign new_n39632_ = ~new_n39353_ & ~new_n39631_;
  assign new_n39633_ = ~new_n39629_ & new_n39632_;
  assign new_n39634_ = ~new_n39353_ & ~new_n39633_;
  assign new_n39635_ = \b[22]  & ~new_n39342_;
  assign new_n39636_ = ~new_n39340_ & new_n39635_;
  assign new_n39637_ = ~new_n39344_ & ~new_n39636_;
  assign new_n39638_ = ~new_n39634_ & new_n39637_;
  assign new_n39639_ = ~new_n39344_ & ~new_n39638_;
  assign new_n39640_ = \b[23]  & ~new_n39333_;
  assign new_n39641_ = ~new_n39331_ & new_n39640_;
  assign new_n39642_ = ~new_n39335_ & ~new_n39641_;
  assign new_n39643_ = ~new_n39639_ & new_n39642_;
  assign new_n39644_ = ~new_n39335_ & ~new_n39643_;
  assign new_n39645_ = \b[24]  & ~new_n39324_;
  assign new_n39646_ = ~new_n39322_ & new_n39645_;
  assign new_n39647_ = ~new_n39326_ & ~new_n39646_;
  assign new_n39648_ = ~new_n39644_ & new_n39647_;
  assign new_n39649_ = ~new_n39326_ & ~new_n39648_;
  assign new_n39650_ = \b[25]  & ~new_n39315_;
  assign new_n39651_ = ~new_n39313_ & new_n39650_;
  assign new_n39652_ = ~new_n39317_ & ~new_n39651_;
  assign new_n39653_ = ~new_n39649_ & new_n39652_;
  assign new_n39654_ = ~new_n39317_ & ~new_n39653_;
  assign new_n39655_ = \b[26]  & ~new_n39306_;
  assign new_n39656_ = ~new_n39304_ & new_n39655_;
  assign new_n39657_ = ~new_n39308_ & ~new_n39656_;
  assign new_n39658_ = ~new_n39654_ & new_n39657_;
  assign new_n39659_ = ~new_n39308_ & ~new_n39658_;
  assign new_n39660_ = \b[27]  & ~new_n39297_;
  assign new_n39661_ = ~new_n39295_ & new_n39660_;
  assign new_n39662_ = ~new_n39299_ & ~new_n39661_;
  assign new_n39663_ = ~new_n39659_ & new_n39662_;
  assign new_n39664_ = ~new_n39299_ & ~new_n39663_;
  assign new_n39665_ = \b[28]  & ~new_n39288_;
  assign new_n39666_ = ~new_n39286_ & new_n39665_;
  assign new_n39667_ = ~new_n39290_ & ~new_n39666_;
  assign new_n39668_ = ~new_n39664_ & new_n39667_;
  assign new_n39669_ = ~new_n39290_ & ~new_n39668_;
  assign new_n39670_ = \b[29]  & ~new_n39279_;
  assign new_n39671_ = ~new_n39277_ & new_n39670_;
  assign new_n39672_ = ~new_n39281_ & ~new_n39671_;
  assign new_n39673_ = ~new_n39669_ & new_n39672_;
  assign new_n39674_ = ~new_n39281_ & ~new_n39673_;
  assign new_n39675_ = \b[30]  & ~new_n39270_;
  assign new_n39676_ = ~new_n39268_ & new_n39675_;
  assign new_n39677_ = ~new_n39272_ & ~new_n39676_;
  assign new_n39678_ = ~new_n39674_ & new_n39677_;
  assign new_n39679_ = ~new_n39272_ & ~new_n39678_;
  assign new_n39680_ = \b[31]  & ~new_n39261_;
  assign new_n39681_ = ~new_n39259_ & new_n39680_;
  assign new_n39682_ = ~new_n39263_ & ~new_n39681_;
  assign new_n39683_ = ~new_n39679_ & new_n39682_;
  assign new_n39684_ = ~new_n39263_ & ~new_n39683_;
  assign new_n39685_ = \b[32]  & ~new_n39252_;
  assign new_n39686_ = ~new_n39250_ & new_n39685_;
  assign new_n39687_ = ~new_n39254_ & ~new_n39686_;
  assign new_n39688_ = ~new_n39684_ & new_n39687_;
  assign new_n39689_ = ~new_n39254_ & ~new_n39688_;
  assign new_n39690_ = \b[33]  & ~new_n39243_;
  assign new_n39691_ = ~new_n39241_ & new_n39690_;
  assign new_n39692_ = ~new_n39245_ & ~new_n39691_;
  assign new_n39693_ = ~new_n39689_ & new_n39692_;
  assign new_n39694_ = ~new_n39245_ & ~new_n39693_;
  assign new_n39695_ = \b[34]  & ~new_n39234_;
  assign new_n39696_ = ~new_n39232_ & new_n39695_;
  assign new_n39697_ = ~new_n39236_ & ~new_n39696_;
  assign new_n39698_ = ~new_n39694_ & new_n39697_;
  assign new_n39699_ = ~new_n39236_ & ~new_n39698_;
  assign new_n39700_ = \b[35]  & ~new_n39225_;
  assign new_n39701_ = ~new_n39223_ & new_n39700_;
  assign new_n39702_ = ~new_n39227_ & ~new_n39701_;
  assign new_n39703_ = ~new_n39699_ & new_n39702_;
  assign new_n39704_ = ~new_n39227_ & ~new_n39703_;
  assign new_n39705_ = \b[36]  & ~new_n39216_;
  assign new_n39706_ = ~new_n39214_ & new_n39705_;
  assign new_n39707_ = ~new_n39218_ & ~new_n39706_;
  assign new_n39708_ = ~new_n39704_ & new_n39707_;
  assign new_n39709_ = ~new_n39218_ & ~new_n39708_;
  assign new_n39710_ = \b[37]  & ~new_n39207_;
  assign new_n39711_ = ~new_n39205_ & new_n39710_;
  assign new_n39712_ = ~new_n39209_ & ~new_n39711_;
  assign new_n39713_ = ~new_n39709_ & new_n39712_;
  assign new_n39714_ = ~new_n39209_ & ~new_n39713_;
  assign new_n39715_ = \b[38]  & ~new_n39187_;
  assign new_n39716_ = ~new_n39185_ & new_n39715_;
  assign new_n39717_ = ~new_n39200_ & ~new_n39716_;
  assign new_n39718_ = ~new_n39714_ & new_n39717_;
  assign new_n39719_ = ~new_n39200_ & ~new_n39718_;
  assign new_n39720_ = \b[39]  & ~new_n39197_;
  assign new_n39721_ = ~new_n39195_ & new_n39720_;
  assign new_n39722_ = ~new_n39199_ & ~new_n39721_;
  assign new_n39723_ = ~new_n39719_ & new_n39722_;
  assign new_n39724_ = ~new_n39199_ & ~new_n39723_;
  assign new_n39725_ = new_n11619_ & ~new_n39724_;
  assign new_n39726_ = ~new_n39188_ & ~new_n39725_;
  assign new_n39727_ = ~new_n39209_ & new_n39717_;
  assign new_n39728_ = ~new_n39713_ & new_n39727_;
  assign new_n39729_ = ~new_n39714_ & ~new_n39717_;
  assign new_n39730_ = ~new_n39728_ & ~new_n39729_;
  assign new_n39731_ = new_n11619_ & ~new_n39730_;
  assign new_n39732_ = ~new_n39724_ & new_n39731_;
  assign new_n39733_ = ~new_n39726_ & ~new_n39732_;
  assign new_n39734_ = ~new_n39198_ & ~new_n39725_;
  assign new_n39735_ = ~new_n39200_ & new_n39722_;
  assign new_n39736_ = ~new_n39718_ & new_n39735_;
  assign new_n39737_ = ~new_n39719_ & ~new_n39722_;
  assign new_n39738_ = ~new_n39736_ & ~new_n39737_;
  assign new_n39739_ = new_n39725_ & ~new_n39738_;
  assign new_n39740_ = ~new_n39734_ & ~new_n39739_;
  assign new_n39741_ = ~\b[40]  & ~new_n39740_;
  assign new_n39742_ = ~\b[39]  & ~new_n39733_;
  assign new_n39743_ = ~new_n39208_ & ~new_n39725_;
  assign new_n39744_ = ~new_n39218_ & new_n39712_;
  assign new_n39745_ = ~new_n39708_ & new_n39744_;
  assign new_n39746_ = ~new_n39709_ & ~new_n39712_;
  assign new_n39747_ = ~new_n39745_ & ~new_n39746_;
  assign new_n39748_ = new_n11619_ & ~new_n39747_;
  assign new_n39749_ = ~new_n39724_ & new_n39748_;
  assign new_n39750_ = ~new_n39743_ & ~new_n39749_;
  assign new_n39751_ = ~\b[38]  & ~new_n39750_;
  assign new_n39752_ = ~new_n39217_ & ~new_n39725_;
  assign new_n39753_ = ~new_n39227_ & new_n39707_;
  assign new_n39754_ = ~new_n39703_ & new_n39753_;
  assign new_n39755_ = ~new_n39704_ & ~new_n39707_;
  assign new_n39756_ = ~new_n39754_ & ~new_n39755_;
  assign new_n39757_ = new_n11619_ & ~new_n39756_;
  assign new_n39758_ = ~new_n39724_ & new_n39757_;
  assign new_n39759_ = ~new_n39752_ & ~new_n39758_;
  assign new_n39760_ = ~\b[37]  & ~new_n39759_;
  assign new_n39761_ = ~new_n39226_ & ~new_n39725_;
  assign new_n39762_ = ~new_n39236_ & new_n39702_;
  assign new_n39763_ = ~new_n39698_ & new_n39762_;
  assign new_n39764_ = ~new_n39699_ & ~new_n39702_;
  assign new_n39765_ = ~new_n39763_ & ~new_n39764_;
  assign new_n39766_ = new_n11619_ & ~new_n39765_;
  assign new_n39767_ = ~new_n39724_ & new_n39766_;
  assign new_n39768_ = ~new_n39761_ & ~new_n39767_;
  assign new_n39769_ = ~\b[36]  & ~new_n39768_;
  assign new_n39770_ = ~new_n39235_ & ~new_n39725_;
  assign new_n39771_ = ~new_n39245_ & new_n39697_;
  assign new_n39772_ = ~new_n39693_ & new_n39771_;
  assign new_n39773_ = ~new_n39694_ & ~new_n39697_;
  assign new_n39774_ = ~new_n39772_ & ~new_n39773_;
  assign new_n39775_ = new_n11619_ & ~new_n39774_;
  assign new_n39776_ = ~new_n39724_ & new_n39775_;
  assign new_n39777_ = ~new_n39770_ & ~new_n39776_;
  assign new_n39778_ = ~\b[35]  & ~new_n39777_;
  assign new_n39779_ = ~new_n39244_ & ~new_n39725_;
  assign new_n39780_ = ~new_n39254_ & new_n39692_;
  assign new_n39781_ = ~new_n39688_ & new_n39780_;
  assign new_n39782_ = ~new_n39689_ & ~new_n39692_;
  assign new_n39783_ = ~new_n39781_ & ~new_n39782_;
  assign new_n39784_ = new_n11619_ & ~new_n39783_;
  assign new_n39785_ = ~new_n39724_ & new_n39784_;
  assign new_n39786_ = ~new_n39779_ & ~new_n39785_;
  assign new_n39787_ = ~\b[34]  & ~new_n39786_;
  assign new_n39788_ = ~new_n39253_ & ~new_n39725_;
  assign new_n39789_ = ~new_n39263_ & new_n39687_;
  assign new_n39790_ = ~new_n39683_ & new_n39789_;
  assign new_n39791_ = ~new_n39684_ & ~new_n39687_;
  assign new_n39792_ = ~new_n39790_ & ~new_n39791_;
  assign new_n39793_ = new_n11619_ & ~new_n39792_;
  assign new_n39794_ = ~new_n39724_ & new_n39793_;
  assign new_n39795_ = ~new_n39788_ & ~new_n39794_;
  assign new_n39796_ = ~\b[33]  & ~new_n39795_;
  assign new_n39797_ = ~new_n39262_ & ~new_n39725_;
  assign new_n39798_ = ~new_n39272_ & new_n39682_;
  assign new_n39799_ = ~new_n39678_ & new_n39798_;
  assign new_n39800_ = ~new_n39679_ & ~new_n39682_;
  assign new_n39801_ = ~new_n39799_ & ~new_n39800_;
  assign new_n39802_ = new_n11619_ & ~new_n39801_;
  assign new_n39803_ = ~new_n39724_ & new_n39802_;
  assign new_n39804_ = ~new_n39797_ & ~new_n39803_;
  assign new_n39805_ = ~\b[32]  & ~new_n39804_;
  assign new_n39806_ = ~new_n39271_ & ~new_n39725_;
  assign new_n39807_ = ~new_n39281_ & new_n39677_;
  assign new_n39808_ = ~new_n39673_ & new_n39807_;
  assign new_n39809_ = ~new_n39674_ & ~new_n39677_;
  assign new_n39810_ = ~new_n39808_ & ~new_n39809_;
  assign new_n39811_ = new_n11619_ & ~new_n39810_;
  assign new_n39812_ = ~new_n39724_ & new_n39811_;
  assign new_n39813_ = ~new_n39806_ & ~new_n39812_;
  assign new_n39814_ = ~\b[31]  & ~new_n39813_;
  assign new_n39815_ = ~new_n39280_ & ~new_n39725_;
  assign new_n39816_ = ~new_n39290_ & new_n39672_;
  assign new_n39817_ = ~new_n39668_ & new_n39816_;
  assign new_n39818_ = ~new_n39669_ & ~new_n39672_;
  assign new_n39819_ = ~new_n39817_ & ~new_n39818_;
  assign new_n39820_ = new_n11619_ & ~new_n39819_;
  assign new_n39821_ = ~new_n39724_ & new_n39820_;
  assign new_n39822_ = ~new_n39815_ & ~new_n39821_;
  assign new_n39823_ = ~\b[30]  & ~new_n39822_;
  assign new_n39824_ = ~new_n39289_ & ~new_n39725_;
  assign new_n39825_ = ~new_n39299_ & new_n39667_;
  assign new_n39826_ = ~new_n39663_ & new_n39825_;
  assign new_n39827_ = ~new_n39664_ & ~new_n39667_;
  assign new_n39828_ = ~new_n39826_ & ~new_n39827_;
  assign new_n39829_ = new_n11619_ & ~new_n39828_;
  assign new_n39830_ = ~new_n39724_ & new_n39829_;
  assign new_n39831_ = ~new_n39824_ & ~new_n39830_;
  assign new_n39832_ = ~\b[29]  & ~new_n39831_;
  assign new_n39833_ = ~new_n39298_ & ~new_n39725_;
  assign new_n39834_ = ~new_n39308_ & new_n39662_;
  assign new_n39835_ = ~new_n39658_ & new_n39834_;
  assign new_n39836_ = ~new_n39659_ & ~new_n39662_;
  assign new_n39837_ = ~new_n39835_ & ~new_n39836_;
  assign new_n39838_ = new_n11619_ & ~new_n39837_;
  assign new_n39839_ = ~new_n39724_ & new_n39838_;
  assign new_n39840_ = ~new_n39833_ & ~new_n39839_;
  assign new_n39841_ = ~\b[28]  & ~new_n39840_;
  assign new_n39842_ = ~new_n39307_ & ~new_n39725_;
  assign new_n39843_ = ~new_n39317_ & new_n39657_;
  assign new_n39844_ = ~new_n39653_ & new_n39843_;
  assign new_n39845_ = ~new_n39654_ & ~new_n39657_;
  assign new_n39846_ = ~new_n39844_ & ~new_n39845_;
  assign new_n39847_ = new_n11619_ & ~new_n39846_;
  assign new_n39848_ = ~new_n39724_ & new_n39847_;
  assign new_n39849_ = ~new_n39842_ & ~new_n39848_;
  assign new_n39850_ = ~\b[27]  & ~new_n39849_;
  assign new_n39851_ = ~new_n39316_ & ~new_n39725_;
  assign new_n39852_ = ~new_n39326_ & new_n39652_;
  assign new_n39853_ = ~new_n39648_ & new_n39852_;
  assign new_n39854_ = ~new_n39649_ & ~new_n39652_;
  assign new_n39855_ = ~new_n39853_ & ~new_n39854_;
  assign new_n39856_ = new_n11619_ & ~new_n39855_;
  assign new_n39857_ = ~new_n39724_ & new_n39856_;
  assign new_n39858_ = ~new_n39851_ & ~new_n39857_;
  assign new_n39859_ = ~\b[26]  & ~new_n39858_;
  assign new_n39860_ = ~new_n39325_ & ~new_n39725_;
  assign new_n39861_ = ~new_n39335_ & new_n39647_;
  assign new_n39862_ = ~new_n39643_ & new_n39861_;
  assign new_n39863_ = ~new_n39644_ & ~new_n39647_;
  assign new_n39864_ = ~new_n39862_ & ~new_n39863_;
  assign new_n39865_ = new_n11619_ & ~new_n39864_;
  assign new_n39866_ = ~new_n39724_ & new_n39865_;
  assign new_n39867_ = ~new_n39860_ & ~new_n39866_;
  assign new_n39868_ = ~\b[25]  & ~new_n39867_;
  assign new_n39869_ = ~new_n39334_ & ~new_n39725_;
  assign new_n39870_ = ~new_n39344_ & new_n39642_;
  assign new_n39871_ = ~new_n39638_ & new_n39870_;
  assign new_n39872_ = ~new_n39639_ & ~new_n39642_;
  assign new_n39873_ = ~new_n39871_ & ~new_n39872_;
  assign new_n39874_ = new_n11619_ & ~new_n39873_;
  assign new_n39875_ = ~new_n39724_ & new_n39874_;
  assign new_n39876_ = ~new_n39869_ & ~new_n39875_;
  assign new_n39877_ = ~\b[24]  & ~new_n39876_;
  assign new_n39878_ = ~new_n39343_ & ~new_n39725_;
  assign new_n39879_ = ~new_n39353_ & new_n39637_;
  assign new_n39880_ = ~new_n39633_ & new_n39879_;
  assign new_n39881_ = ~new_n39634_ & ~new_n39637_;
  assign new_n39882_ = ~new_n39880_ & ~new_n39881_;
  assign new_n39883_ = new_n11619_ & ~new_n39882_;
  assign new_n39884_ = ~new_n39724_ & new_n39883_;
  assign new_n39885_ = ~new_n39878_ & ~new_n39884_;
  assign new_n39886_ = ~\b[23]  & ~new_n39885_;
  assign new_n39887_ = ~new_n39352_ & ~new_n39725_;
  assign new_n39888_ = ~new_n39362_ & new_n39632_;
  assign new_n39889_ = ~new_n39628_ & new_n39888_;
  assign new_n39890_ = ~new_n39629_ & ~new_n39632_;
  assign new_n39891_ = ~new_n39889_ & ~new_n39890_;
  assign new_n39892_ = new_n11619_ & ~new_n39891_;
  assign new_n39893_ = ~new_n39724_ & new_n39892_;
  assign new_n39894_ = ~new_n39887_ & ~new_n39893_;
  assign new_n39895_ = ~\b[22]  & ~new_n39894_;
  assign new_n39896_ = ~new_n39361_ & ~new_n39725_;
  assign new_n39897_ = ~new_n39371_ & new_n39627_;
  assign new_n39898_ = ~new_n39623_ & new_n39897_;
  assign new_n39899_ = ~new_n39624_ & ~new_n39627_;
  assign new_n39900_ = ~new_n39898_ & ~new_n39899_;
  assign new_n39901_ = new_n11619_ & ~new_n39900_;
  assign new_n39902_ = ~new_n39724_ & new_n39901_;
  assign new_n39903_ = ~new_n39896_ & ~new_n39902_;
  assign new_n39904_ = ~\b[21]  & ~new_n39903_;
  assign new_n39905_ = ~new_n39370_ & ~new_n39725_;
  assign new_n39906_ = ~new_n39380_ & new_n39622_;
  assign new_n39907_ = ~new_n39618_ & new_n39906_;
  assign new_n39908_ = ~new_n39619_ & ~new_n39622_;
  assign new_n39909_ = ~new_n39907_ & ~new_n39908_;
  assign new_n39910_ = new_n11619_ & ~new_n39909_;
  assign new_n39911_ = ~new_n39724_ & new_n39910_;
  assign new_n39912_ = ~new_n39905_ & ~new_n39911_;
  assign new_n39913_ = ~\b[20]  & ~new_n39912_;
  assign new_n39914_ = ~new_n39379_ & ~new_n39725_;
  assign new_n39915_ = ~new_n39389_ & new_n39617_;
  assign new_n39916_ = ~new_n39613_ & new_n39915_;
  assign new_n39917_ = ~new_n39614_ & ~new_n39617_;
  assign new_n39918_ = ~new_n39916_ & ~new_n39917_;
  assign new_n39919_ = new_n11619_ & ~new_n39918_;
  assign new_n39920_ = ~new_n39724_ & new_n39919_;
  assign new_n39921_ = ~new_n39914_ & ~new_n39920_;
  assign new_n39922_ = ~\b[19]  & ~new_n39921_;
  assign new_n39923_ = ~new_n39388_ & ~new_n39725_;
  assign new_n39924_ = ~new_n39398_ & new_n39612_;
  assign new_n39925_ = ~new_n39608_ & new_n39924_;
  assign new_n39926_ = ~new_n39609_ & ~new_n39612_;
  assign new_n39927_ = ~new_n39925_ & ~new_n39926_;
  assign new_n39928_ = new_n11619_ & ~new_n39927_;
  assign new_n39929_ = ~new_n39724_ & new_n39928_;
  assign new_n39930_ = ~new_n39923_ & ~new_n39929_;
  assign new_n39931_ = ~\b[18]  & ~new_n39930_;
  assign new_n39932_ = ~new_n39397_ & ~new_n39725_;
  assign new_n39933_ = ~new_n39407_ & new_n39607_;
  assign new_n39934_ = ~new_n39603_ & new_n39933_;
  assign new_n39935_ = ~new_n39604_ & ~new_n39607_;
  assign new_n39936_ = ~new_n39934_ & ~new_n39935_;
  assign new_n39937_ = new_n11619_ & ~new_n39936_;
  assign new_n39938_ = ~new_n39724_ & new_n39937_;
  assign new_n39939_ = ~new_n39932_ & ~new_n39938_;
  assign new_n39940_ = ~\b[17]  & ~new_n39939_;
  assign new_n39941_ = ~new_n39406_ & ~new_n39725_;
  assign new_n39942_ = ~new_n39416_ & new_n39602_;
  assign new_n39943_ = ~new_n39598_ & new_n39942_;
  assign new_n39944_ = ~new_n39599_ & ~new_n39602_;
  assign new_n39945_ = ~new_n39943_ & ~new_n39944_;
  assign new_n39946_ = new_n11619_ & ~new_n39945_;
  assign new_n39947_ = ~new_n39724_ & new_n39946_;
  assign new_n39948_ = ~new_n39941_ & ~new_n39947_;
  assign new_n39949_ = ~\b[16]  & ~new_n39948_;
  assign new_n39950_ = ~new_n39415_ & ~new_n39725_;
  assign new_n39951_ = ~new_n39425_ & new_n39597_;
  assign new_n39952_ = ~new_n39593_ & new_n39951_;
  assign new_n39953_ = ~new_n39594_ & ~new_n39597_;
  assign new_n39954_ = ~new_n39952_ & ~new_n39953_;
  assign new_n39955_ = new_n11619_ & ~new_n39954_;
  assign new_n39956_ = ~new_n39724_ & new_n39955_;
  assign new_n39957_ = ~new_n39950_ & ~new_n39956_;
  assign new_n39958_ = ~\b[15]  & ~new_n39957_;
  assign new_n39959_ = ~new_n39424_ & ~new_n39725_;
  assign new_n39960_ = ~new_n39434_ & new_n39592_;
  assign new_n39961_ = ~new_n39588_ & new_n39960_;
  assign new_n39962_ = ~new_n39589_ & ~new_n39592_;
  assign new_n39963_ = ~new_n39961_ & ~new_n39962_;
  assign new_n39964_ = new_n11619_ & ~new_n39963_;
  assign new_n39965_ = ~new_n39724_ & new_n39964_;
  assign new_n39966_ = ~new_n39959_ & ~new_n39965_;
  assign new_n39967_ = ~\b[14]  & ~new_n39966_;
  assign new_n39968_ = ~new_n39433_ & ~new_n39725_;
  assign new_n39969_ = ~new_n39443_ & new_n39587_;
  assign new_n39970_ = ~new_n39583_ & new_n39969_;
  assign new_n39971_ = ~new_n39584_ & ~new_n39587_;
  assign new_n39972_ = ~new_n39970_ & ~new_n39971_;
  assign new_n39973_ = new_n11619_ & ~new_n39972_;
  assign new_n39974_ = ~new_n39724_ & new_n39973_;
  assign new_n39975_ = ~new_n39968_ & ~new_n39974_;
  assign new_n39976_ = ~\b[13]  & ~new_n39975_;
  assign new_n39977_ = ~new_n39442_ & ~new_n39725_;
  assign new_n39978_ = ~new_n39452_ & new_n39582_;
  assign new_n39979_ = ~new_n39578_ & new_n39978_;
  assign new_n39980_ = ~new_n39579_ & ~new_n39582_;
  assign new_n39981_ = ~new_n39979_ & ~new_n39980_;
  assign new_n39982_ = new_n11619_ & ~new_n39981_;
  assign new_n39983_ = ~new_n39724_ & new_n39982_;
  assign new_n39984_ = ~new_n39977_ & ~new_n39983_;
  assign new_n39985_ = ~\b[12]  & ~new_n39984_;
  assign new_n39986_ = ~new_n39451_ & ~new_n39725_;
  assign new_n39987_ = ~new_n39461_ & new_n39577_;
  assign new_n39988_ = ~new_n39573_ & new_n39987_;
  assign new_n39989_ = ~new_n39574_ & ~new_n39577_;
  assign new_n39990_ = ~new_n39988_ & ~new_n39989_;
  assign new_n39991_ = new_n11619_ & ~new_n39990_;
  assign new_n39992_ = ~new_n39724_ & new_n39991_;
  assign new_n39993_ = ~new_n39986_ & ~new_n39992_;
  assign new_n39994_ = ~\b[11]  & ~new_n39993_;
  assign new_n39995_ = ~new_n39460_ & ~new_n39725_;
  assign new_n39996_ = ~new_n39470_ & new_n39572_;
  assign new_n39997_ = ~new_n39568_ & new_n39996_;
  assign new_n39998_ = ~new_n39569_ & ~new_n39572_;
  assign new_n39999_ = ~new_n39997_ & ~new_n39998_;
  assign new_n40000_ = new_n11619_ & ~new_n39999_;
  assign new_n40001_ = ~new_n39724_ & new_n40000_;
  assign new_n40002_ = ~new_n39995_ & ~new_n40001_;
  assign new_n40003_ = ~\b[10]  & ~new_n40002_;
  assign new_n40004_ = ~new_n39469_ & ~new_n39725_;
  assign new_n40005_ = ~new_n39479_ & new_n39567_;
  assign new_n40006_ = ~new_n39563_ & new_n40005_;
  assign new_n40007_ = ~new_n39564_ & ~new_n39567_;
  assign new_n40008_ = ~new_n40006_ & ~new_n40007_;
  assign new_n40009_ = new_n11619_ & ~new_n40008_;
  assign new_n40010_ = ~new_n39724_ & new_n40009_;
  assign new_n40011_ = ~new_n40004_ & ~new_n40010_;
  assign new_n40012_ = ~\b[9]  & ~new_n40011_;
  assign new_n40013_ = ~new_n39478_ & ~new_n39725_;
  assign new_n40014_ = ~new_n39488_ & new_n39562_;
  assign new_n40015_ = ~new_n39558_ & new_n40014_;
  assign new_n40016_ = ~new_n39559_ & ~new_n39562_;
  assign new_n40017_ = ~new_n40015_ & ~new_n40016_;
  assign new_n40018_ = new_n11619_ & ~new_n40017_;
  assign new_n40019_ = ~new_n39724_ & new_n40018_;
  assign new_n40020_ = ~new_n40013_ & ~new_n40019_;
  assign new_n40021_ = ~\b[8]  & ~new_n40020_;
  assign new_n40022_ = ~new_n39487_ & ~new_n39725_;
  assign new_n40023_ = ~new_n39497_ & new_n39557_;
  assign new_n40024_ = ~new_n39553_ & new_n40023_;
  assign new_n40025_ = ~new_n39554_ & ~new_n39557_;
  assign new_n40026_ = ~new_n40024_ & ~new_n40025_;
  assign new_n40027_ = new_n11619_ & ~new_n40026_;
  assign new_n40028_ = ~new_n39724_ & new_n40027_;
  assign new_n40029_ = ~new_n40022_ & ~new_n40028_;
  assign new_n40030_ = ~\b[7]  & ~new_n40029_;
  assign new_n40031_ = ~new_n39496_ & ~new_n39725_;
  assign new_n40032_ = ~new_n39506_ & new_n39552_;
  assign new_n40033_ = ~new_n39548_ & new_n40032_;
  assign new_n40034_ = ~new_n39549_ & ~new_n39552_;
  assign new_n40035_ = ~new_n40033_ & ~new_n40034_;
  assign new_n40036_ = new_n11619_ & ~new_n40035_;
  assign new_n40037_ = ~new_n39724_ & new_n40036_;
  assign new_n40038_ = ~new_n40031_ & ~new_n40037_;
  assign new_n40039_ = ~\b[6]  & ~new_n40038_;
  assign new_n40040_ = ~new_n39505_ & ~new_n39725_;
  assign new_n40041_ = ~new_n39515_ & new_n39547_;
  assign new_n40042_ = ~new_n39543_ & new_n40041_;
  assign new_n40043_ = ~new_n39544_ & ~new_n39547_;
  assign new_n40044_ = ~new_n40042_ & ~new_n40043_;
  assign new_n40045_ = new_n11619_ & ~new_n40044_;
  assign new_n40046_ = ~new_n39724_ & new_n40045_;
  assign new_n40047_ = ~new_n40040_ & ~new_n40046_;
  assign new_n40048_ = ~\b[5]  & ~new_n40047_;
  assign new_n40049_ = ~new_n39514_ & ~new_n39725_;
  assign new_n40050_ = ~new_n39523_ & new_n39542_;
  assign new_n40051_ = ~new_n39538_ & new_n40050_;
  assign new_n40052_ = ~new_n39539_ & ~new_n39542_;
  assign new_n40053_ = ~new_n40051_ & ~new_n40052_;
  assign new_n40054_ = new_n11619_ & ~new_n40053_;
  assign new_n40055_ = ~new_n39724_ & new_n40054_;
  assign new_n40056_ = ~new_n40049_ & ~new_n40055_;
  assign new_n40057_ = ~\b[4]  & ~new_n40056_;
  assign new_n40058_ = ~new_n39522_ & ~new_n39725_;
  assign new_n40059_ = ~new_n39533_ & new_n39537_;
  assign new_n40060_ = ~new_n39532_ & new_n40059_;
  assign new_n40061_ = ~new_n39534_ & ~new_n39537_;
  assign new_n40062_ = ~new_n40060_ & ~new_n40061_;
  assign new_n40063_ = new_n11619_ & ~new_n40062_;
  assign new_n40064_ = ~new_n39724_ & new_n40063_;
  assign new_n40065_ = ~new_n40058_ & ~new_n40064_;
  assign new_n40066_ = ~\b[3]  & ~new_n40065_;
  assign new_n40067_ = ~new_n39527_ & ~new_n39725_;
  assign new_n40068_ = new_n11425_ & ~new_n39530_;
  assign new_n40069_ = ~new_n39528_ & new_n40068_;
  assign new_n40070_ = new_n11619_ & ~new_n40069_;
  assign new_n40071_ = ~new_n39532_ & new_n40070_;
  assign new_n40072_ = ~new_n39724_ & new_n40071_;
  assign new_n40073_ = ~new_n40067_ & ~new_n40072_;
  assign new_n40074_ = ~\b[2]  & ~new_n40073_;
  assign new_n40075_ = new_n11973_ & ~new_n39724_;
  assign new_n40076_ = \a[24]  & ~new_n40075_;
  assign new_n40077_ = new_n11978_ & ~new_n39724_;
  assign new_n40078_ = ~new_n40076_ & ~new_n40077_;
  assign new_n40079_ = \b[1]  & ~new_n40078_;
  assign new_n40080_ = ~\b[1]  & ~new_n40077_;
  assign new_n40081_ = ~new_n40076_ & new_n40080_;
  assign new_n40082_ = ~new_n40079_ & ~new_n40081_;
  assign new_n40083_ = ~new_n11985_ & ~new_n40082_;
  assign new_n40084_ = ~\b[1]  & ~new_n40078_;
  assign new_n40085_ = ~new_n40083_ & ~new_n40084_;
  assign new_n40086_ = \b[2]  & ~new_n40072_;
  assign new_n40087_ = ~new_n40067_ & new_n40086_;
  assign new_n40088_ = ~new_n40074_ & ~new_n40087_;
  assign new_n40089_ = ~new_n40085_ & new_n40088_;
  assign new_n40090_ = ~new_n40074_ & ~new_n40089_;
  assign new_n40091_ = \b[3]  & ~new_n40064_;
  assign new_n40092_ = ~new_n40058_ & new_n40091_;
  assign new_n40093_ = ~new_n40066_ & ~new_n40092_;
  assign new_n40094_ = ~new_n40090_ & new_n40093_;
  assign new_n40095_ = ~new_n40066_ & ~new_n40094_;
  assign new_n40096_ = \b[4]  & ~new_n40055_;
  assign new_n40097_ = ~new_n40049_ & new_n40096_;
  assign new_n40098_ = ~new_n40057_ & ~new_n40097_;
  assign new_n40099_ = ~new_n40095_ & new_n40098_;
  assign new_n40100_ = ~new_n40057_ & ~new_n40099_;
  assign new_n40101_ = \b[5]  & ~new_n40046_;
  assign new_n40102_ = ~new_n40040_ & new_n40101_;
  assign new_n40103_ = ~new_n40048_ & ~new_n40102_;
  assign new_n40104_ = ~new_n40100_ & new_n40103_;
  assign new_n40105_ = ~new_n40048_ & ~new_n40104_;
  assign new_n40106_ = \b[6]  & ~new_n40037_;
  assign new_n40107_ = ~new_n40031_ & new_n40106_;
  assign new_n40108_ = ~new_n40039_ & ~new_n40107_;
  assign new_n40109_ = ~new_n40105_ & new_n40108_;
  assign new_n40110_ = ~new_n40039_ & ~new_n40109_;
  assign new_n40111_ = \b[7]  & ~new_n40028_;
  assign new_n40112_ = ~new_n40022_ & new_n40111_;
  assign new_n40113_ = ~new_n40030_ & ~new_n40112_;
  assign new_n40114_ = ~new_n40110_ & new_n40113_;
  assign new_n40115_ = ~new_n40030_ & ~new_n40114_;
  assign new_n40116_ = \b[8]  & ~new_n40019_;
  assign new_n40117_ = ~new_n40013_ & new_n40116_;
  assign new_n40118_ = ~new_n40021_ & ~new_n40117_;
  assign new_n40119_ = ~new_n40115_ & new_n40118_;
  assign new_n40120_ = ~new_n40021_ & ~new_n40119_;
  assign new_n40121_ = \b[9]  & ~new_n40010_;
  assign new_n40122_ = ~new_n40004_ & new_n40121_;
  assign new_n40123_ = ~new_n40012_ & ~new_n40122_;
  assign new_n40124_ = ~new_n40120_ & new_n40123_;
  assign new_n40125_ = ~new_n40012_ & ~new_n40124_;
  assign new_n40126_ = \b[10]  & ~new_n40001_;
  assign new_n40127_ = ~new_n39995_ & new_n40126_;
  assign new_n40128_ = ~new_n40003_ & ~new_n40127_;
  assign new_n40129_ = ~new_n40125_ & new_n40128_;
  assign new_n40130_ = ~new_n40003_ & ~new_n40129_;
  assign new_n40131_ = \b[11]  & ~new_n39992_;
  assign new_n40132_ = ~new_n39986_ & new_n40131_;
  assign new_n40133_ = ~new_n39994_ & ~new_n40132_;
  assign new_n40134_ = ~new_n40130_ & new_n40133_;
  assign new_n40135_ = ~new_n39994_ & ~new_n40134_;
  assign new_n40136_ = \b[12]  & ~new_n39983_;
  assign new_n40137_ = ~new_n39977_ & new_n40136_;
  assign new_n40138_ = ~new_n39985_ & ~new_n40137_;
  assign new_n40139_ = ~new_n40135_ & new_n40138_;
  assign new_n40140_ = ~new_n39985_ & ~new_n40139_;
  assign new_n40141_ = \b[13]  & ~new_n39974_;
  assign new_n40142_ = ~new_n39968_ & new_n40141_;
  assign new_n40143_ = ~new_n39976_ & ~new_n40142_;
  assign new_n40144_ = ~new_n40140_ & new_n40143_;
  assign new_n40145_ = ~new_n39976_ & ~new_n40144_;
  assign new_n40146_ = \b[14]  & ~new_n39965_;
  assign new_n40147_ = ~new_n39959_ & new_n40146_;
  assign new_n40148_ = ~new_n39967_ & ~new_n40147_;
  assign new_n40149_ = ~new_n40145_ & new_n40148_;
  assign new_n40150_ = ~new_n39967_ & ~new_n40149_;
  assign new_n40151_ = \b[15]  & ~new_n39956_;
  assign new_n40152_ = ~new_n39950_ & new_n40151_;
  assign new_n40153_ = ~new_n39958_ & ~new_n40152_;
  assign new_n40154_ = ~new_n40150_ & new_n40153_;
  assign new_n40155_ = ~new_n39958_ & ~new_n40154_;
  assign new_n40156_ = \b[16]  & ~new_n39947_;
  assign new_n40157_ = ~new_n39941_ & new_n40156_;
  assign new_n40158_ = ~new_n39949_ & ~new_n40157_;
  assign new_n40159_ = ~new_n40155_ & new_n40158_;
  assign new_n40160_ = ~new_n39949_ & ~new_n40159_;
  assign new_n40161_ = \b[17]  & ~new_n39938_;
  assign new_n40162_ = ~new_n39932_ & new_n40161_;
  assign new_n40163_ = ~new_n39940_ & ~new_n40162_;
  assign new_n40164_ = ~new_n40160_ & new_n40163_;
  assign new_n40165_ = ~new_n39940_ & ~new_n40164_;
  assign new_n40166_ = \b[18]  & ~new_n39929_;
  assign new_n40167_ = ~new_n39923_ & new_n40166_;
  assign new_n40168_ = ~new_n39931_ & ~new_n40167_;
  assign new_n40169_ = ~new_n40165_ & new_n40168_;
  assign new_n40170_ = ~new_n39931_ & ~new_n40169_;
  assign new_n40171_ = \b[19]  & ~new_n39920_;
  assign new_n40172_ = ~new_n39914_ & new_n40171_;
  assign new_n40173_ = ~new_n39922_ & ~new_n40172_;
  assign new_n40174_ = ~new_n40170_ & new_n40173_;
  assign new_n40175_ = ~new_n39922_ & ~new_n40174_;
  assign new_n40176_ = \b[20]  & ~new_n39911_;
  assign new_n40177_ = ~new_n39905_ & new_n40176_;
  assign new_n40178_ = ~new_n39913_ & ~new_n40177_;
  assign new_n40179_ = ~new_n40175_ & new_n40178_;
  assign new_n40180_ = ~new_n39913_ & ~new_n40179_;
  assign new_n40181_ = \b[21]  & ~new_n39902_;
  assign new_n40182_ = ~new_n39896_ & new_n40181_;
  assign new_n40183_ = ~new_n39904_ & ~new_n40182_;
  assign new_n40184_ = ~new_n40180_ & new_n40183_;
  assign new_n40185_ = ~new_n39904_ & ~new_n40184_;
  assign new_n40186_ = \b[22]  & ~new_n39893_;
  assign new_n40187_ = ~new_n39887_ & new_n40186_;
  assign new_n40188_ = ~new_n39895_ & ~new_n40187_;
  assign new_n40189_ = ~new_n40185_ & new_n40188_;
  assign new_n40190_ = ~new_n39895_ & ~new_n40189_;
  assign new_n40191_ = \b[23]  & ~new_n39884_;
  assign new_n40192_ = ~new_n39878_ & new_n40191_;
  assign new_n40193_ = ~new_n39886_ & ~new_n40192_;
  assign new_n40194_ = ~new_n40190_ & new_n40193_;
  assign new_n40195_ = ~new_n39886_ & ~new_n40194_;
  assign new_n40196_ = \b[24]  & ~new_n39875_;
  assign new_n40197_ = ~new_n39869_ & new_n40196_;
  assign new_n40198_ = ~new_n39877_ & ~new_n40197_;
  assign new_n40199_ = ~new_n40195_ & new_n40198_;
  assign new_n40200_ = ~new_n39877_ & ~new_n40199_;
  assign new_n40201_ = \b[25]  & ~new_n39866_;
  assign new_n40202_ = ~new_n39860_ & new_n40201_;
  assign new_n40203_ = ~new_n39868_ & ~new_n40202_;
  assign new_n40204_ = ~new_n40200_ & new_n40203_;
  assign new_n40205_ = ~new_n39868_ & ~new_n40204_;
  assign new_n40206_ = \b[26]  & ~new_n39857_;
  assign new_n40207_ = ~new_n39851_ & new_n40206_;
  assign new_n40208_ = ~new_n39859_ & ~new_n40207_;
  assign new_n40209_ = ~new_n40205_ & new_n40208_;
  assign new_n40210_ = ~new_n39859_ & ~new_n40209_;
  assign new_n40211_ = \b[27]  & ~new_n39848_;
  assign new_n40212_ = ~new_n39842_ & new_n40211_;
  assign new_n40213_ = ~new_n39850_ & ~new_n40212_;
  assign new_n40214_ = ~new_n40210_ & new_n40213_;
  assign new_n40215_ = ~new_n39850_ & ~new_n40214_;
  assign new_n40216_ = \b[28]  & ~new_n39839_;
  assign new_n40217_ = ~new_n39833_ & new_n40216_;
  assign new_n40218_ = ~new_n39841_ & ~new_n40217_;
  assign new_n40219_ = ~new_n40215_ & new_n40218_;
  assign new_n40220_ = ~new_n39841_ & ~new_n40219_;
  assign new_n40221_ = \b[29]  & ~new_n39830_;
  assign new_n40222_ = ~new_n39824_ & new_n40221_;
  assign new_n40223_ = ~new_n39832_ & ~new_n40222_;
  assign new_n40224_ = ~new_n40220_ & new_n40223_;
  assign new_n40225_ = ~new_n39832_ & ~new_n40224_;
  assign new_n40226_ = \b[30]  & ~new_n39821_;
  assign new_n40227_ = ~new_n39815_ & new_n40226_;
  assign new_n40228_ = ~new_n39823_ & ~new_n40227_;
  assign new_n40229_ = ~new_n40225_ & new_n40228_;
  assign new_n40230_ = ~new_n39823_ & ~new_n40229_;
  assign new_n40231_ = \b[31]  & ~new_n39812_;
  assign new_n40232_ = ~new_n39806_ & new_n40231_;
  assign new_n40233_ = ~new_n39814_ & ~new_n40232_;
  assign new_n40234_ = ~new_n40230_ & new_n40233_;
  assign new_n40235_ = ~new_n39814_ & ~new_n40234_;
  assign new_n40236_ = \b[32]  & ~new_n39803_;
  assign new_n40237_ = ~new_n39797_ & new_n40236_;
  assign new_n40238_ = ~new_n39805_ & ~new_n40237_;
  assign new_n40239_ = ~new_n40235_ & new_n40238_;
  assign new_n40240_ = ~new_n39805_ & ~new_n40239_;
  assign new_n40241_ = \b[33]  & ~new_n39794_;
  assign new_n40242_ = ~new_n39788_ & new_n40241_;
  assign new_n40243_ = ~new_n39796_ & ~new_n40242_;
  assign new_n40244_ = ~new_n40240_ & new_n40243_;
  assign new_n40245_ = ~new_n39796_ & ~new_n40244_;
  assign new_n40246_ = \b[34]  & ~new_n39785_;
  assign new_n40247_ = ~new_n39779_ & new_n40246_;
  assign new_n40248_ = ~new_n39787_ & ~new_n40247_;
  assign new_n40249_ = ~new_n40245_ & new_n40248_;
  assign new_n40250_ = ~new_n39787_ & ~new_n40249_;
  assign new_n40251_ = \b[35]  & ~new_n39776_;
  assign new_n40252_ = ~new_n39770_ & new_n40251_;
  assign new_n40253_ = ~new_n39778_ & ~new_n40252_;
  assign new_n40254_ = ~new_n40250_ & new_n40253_;
  assign new_n40255_ = ~new_n39778_ & ~new_n40254_;
  assign new_n40256_ = \b[36]  & ~new_n39767_;
  assign new_n40257_ = ~new_n39761_ & new_n40256_;
  assign new_n40258_ = ~new_n39769_ & ~new_n40257_;
  assign new_n40259_ = ~new_n40255_ & new_n40258_;
  assign new_n40260_ = ~new_n39769_ & ~new_n40259_;
  assign new_n40261_ = \b[37]  & ~new_n39758_;
  assign new_n40262_ = ~new_n39752_ & new_n40261_;
  assign new_n40263_ = ~new_n39760_ & ~new_n40262_;
  assign new_n40264_ = ~new_n40260_ & new_n40263_;
  assign new_n40265_ = ~new_n39760_ & ~new_n40264_;
  assign new_n40266_ = \b[38]  & ~new_n39749_;
  assign new_n40267_ = ~new_n39743_ & new_n40266_;
  assign new_n40268_ = ~new_n39751_ & ~new_n40267_;
  assign new_n40269_ = ~new_n40265_ & new_n40268_;
  assign new_n40270_ = ~new_n39751_ & ~new_n40269_;
  assign new_n40271_ = \b[39]  & ~new_n39732_;
  assign new_n40272_ = ~new_n39726_ & new_n40271_;
  assign new_n40273_ = ~new_n39742_ & ~new_n40272_;
  assign new_n40274_ = ~new_n40270_ & new_n40273_;
  assign new_n40275_ = ~new_n39742_ & ~new_n40274_;
  assign new_n40276_ = \b[40]  & ~new_n39734_;
  assign new_n40277_ = ~new_n39739_ & new_n40276_;
  assign new_n40278_ = ~new_n39741_ & ~new_n40277_;
  assign new_n40279_ = ~new_n40275_ & new_n40278_;
  assign new_n40280_ = ~new_n39741_ & ~new_n40279_;
  assign new_n40281_ = new_n12184_ & ~new_n40280_;
  assign new_n40282_ = ~new_n39733_ & ~new_n40281_;
  assign new_n40283_ = ~new_n39751_ & new_n40273_;
  assign new_n40284_ = ~new_n40269_ & new_n40283_;
  assign new_n40285_ = ~new_n40270_ & ~new_n40273_;
  assign new_n40286_ = ~new_n40284_ & ~new_n40285_;
  assign new_n40287_ = new_n12184_ & ~new_n40286_;
  assign new_n40288_ = ~new_n40280_ & new_n40287_;
  assign new_n40289_ = ~new_n40282_ & ~new_n40288_;
  assign new_n40290_ = ~\b[40]  & ~new_n40289_;
  assign new_n40291_ = ~new_n39750_ & ~new_n40281_;
  assign new_n40292_ = ~new_n39760_ & new_n40268_;
  assign new_n40293_ = ~new_n40264_ & new_n40292_;
  assign new_n40294_ = ~new_n40265_ & ~new_n40268_;
  assign new_n40295_ = ~new_n40293_ & ~new_n40294_;
  assign new_n40296_ = new_n12184_ & ~new_n40295_;
  assign new_n40297_ = ~new_n40280_ & new_n40296_;
  assign new_n40298_ = ~new_n40291_ & ~new_n40297_;
  assign new_n40299_ = ~\b[39]  & ~new_n40298_;
  assign new_n40300_ = ~new_n39759_ & ~new_n40281_;
  assign new_n40301_ = ~new_n39769_ & new_n40263_;
  assign new_n40302_ = ~new_n40259_ & new_n40301_;
  assign new_n40303_ = ~new_n40260_ & ~new_n40263_;
  assign new_n40304_ = ~new_n40302_ & ~new_n40303_;
  assign new_n40305_ = new_n12184_ & ~new_n40304_;
  assign new_n40306_ = ~new_n40280_ & new_n40305_;
  assign new_n40307_ = ~new_n40300_ & ~new_n40306_;
  assign new_n40308_ = ~\b[38]  & ~new_n40307_;
  assign new_n40309_ = ~new_n39768_ & ~new_n40281_;
  assign new_n40310_ = ~new_n39778_ & new_n40258_;
  assign new_n40311_ = ~new_n40254_ & new_n40310_;
  assign new_n40312_ = ~new_n40255_ & ~new_n40258_;
  assign new_n40313_ = ~new_n40311_ & ~new_n40312_;
  assign new_n40314_ = new_n12184_ & ~new_n40313_;
  assign new_n40315_ = ~new_n40280_ & new_n40314_;
  assign new_n40316_ = ~new_n40309_ & ~new_n40315_;
  assign new_n40317_ = ~\b[37]  & ~new_n40316_;
  assign new_n40318_ = ~new_n39777_ & ~new_n40281_;
  assign new_n40319_ = ~new_n39787_ & new_n40253_;
  assign new_n40320_ = ~new_n40249_ & new_n40319_;
  assign new_n40321_ = ~new_n40250_ & ~new_n40253_;
  assign new_n40322_ = ~new_n40320_ & ~new_n40321_;
  assign new_n40323_ = new_n12184_ & ~new_n40322_;
  assign new_n40324_ = ~new_n40280_ & new_n40323_;
  assign new_n40325_ = ~new_n40318_ & ~new_n40324_;
  assign new_n40326_ = ~\b[36]  & ~new_n40325_;
  assign new_n40327_ = ~new_n39786_ & ~new_n40281_;
  assign new_n40328_ = ~new_n39796_ & new_n40248_;
  assign new_n40329_ = ~new_n40244_ & new_n40328_;
  assign new_n40330_ = ~new_n40245_ & ~new_n40248_;
  assign new_n40331_ = ~new_n40329_ & ~new_n40330_;
  assign new_n40332_ = new_n12184_ & ~new_n40331_;
  assign new_n40333_ = ~new_n40280_ & new_n40332_;
  assign new_n40334_ = ~new_n40327_ & ~new_n40333_;
  assign new_n40335_ = ~\b[35]  & ~new_n40334_;
  assign new_n40336_ = ~new_n39795_ & ~new_n40281_;
  assign new_n40337_ = ~new_n39805_ & new_n40243_;
  assign new_n40338_ = ~new_n40239_ & new_n40337_;
  assign new_n40339_ = ~new_n40240_ & ~new_n40243_;
  assign new_n40340_ = ~new_n40338_ & ~new_n40339_;
  assign new_n40341_ = new_n12184_ & ~new_n40340_;
  assign new_n40342_ = ~new_n40280_ & new_n40341_;
  assign new_n40343_ = ~new_n40336_ & ~new_n40342_;
  assign new_n40344_ = ~\b[34]  & ~new_n40343_;
  assign new_n40345_ = ~new_n39804_ & ~new_n40281_;
  assign new_n40346_ = ~new_n39814_ & new_n40238_;
  assign new_n40347_ = ~new_n40234_ & new_n40346_;
  assign new_n40348_ = ~new_n40235_ & ~new_n40238_;
  assign new_n40349_ = ~new_n40347_ & ~new_n40348_;
  assign new_n40350_ = new_n12184_ & ~new_n40349_;
  assign new_n40351_ = ~new_n40280_ & new_n40350_;
  assign new_n40352_ = ~new_n40345_ & ~new_n40351_;
  assign new_n40353_ = ~\b[33]  & ~new_n40352_;
  assign new_n40354_ = ~new_n39813_ & ~new_n40281_;
  assign new_n40355_ = ~new_n39823_ & new_n40233_;
  assign new_n40356_ = ~new_n40229_ & new_n40355_;
  assign new_n40357_ = ~new_n40230_ & ~new_n40233_;
  assign new_n40358_ = ~new_n40356_ & ~new_n40357_;
  assign new_n40359_ = new_n12184_ & ~new_n40358_;
  assign new_n40360_ = ~new_n40280_ & new_n40359_;
  assign new_n40361_ = ~new_n40354_ & ~new_n40360_;
  assign new_n40362_ = ~\b[32]  & ~new_n40361_;
  assign new_n40363_ = ~new_n39822_ & ~new_n40281_;
  assign new_n40364_ = ~new_n39832_ & new_n40228_;
  assign new_n40365_ = ~new_n40224_ & new_n40364_;
  assign new_n40366_ = ~new_n40225_ & ~new_n40228_;
  assign new_n40367_ = ~new_n40365_ & ~new_n40366_;
  assign new_n40368_ = new_n12184_ & ~new_n40367_;
  assign new_n40369_ = ~new_n40280_ & new_n40368_;
  assign new_n40370_ = ~new_n40363_ & ~new_n40369_;
  assign new_n40371_ = ~\b[31]  & ~new_n40370_;
  assign new_n40372_ = ~new_n39831_ & ~new_n40281_;
  assign new_n40373_ = ~new_n39841_ & new_n40223_;
  assign new_n40374_ = ~new_n40219_ & new_n40373_;
  assign new_n40375_ = ~new_n40220_ & ~new_n40223_;
  assign new_n40376_ = ~new_n40374_ & ~new_n40375_;
  assign new_n40377_ = new_n12184_ & ~new_n40376_;
  assign new_n40378_ = ~new_n40280_ & new_n40377_;
  assign new_n40379_ = ~new_n40372_ & ~new_n40378_;
  assign new_n40380_ = ~\b[30]  & ~new_n40379_;
  assign new_n40381_ = ~new_n39840_ & ~new_n40281_;
  assign new_n40382_ = ~new_n39850_ & new_n40218_;
  assign new_n40383_ = ~new_n40214_ & new_n40382_;
  assign new_n40384_ = ~new_n40215_ & ~new_n40218_;
  assign new_n40385_ = ~new_n40383_ & ~new_n40384_;
  assign new_n40386_ = new_n12184_ & ~new_n40385_;
  assign new_n40387_ = ~new_n40280_ & new_n40386_;
  assign new_n40388_ = ~new_n40381_ & ~new_n40387_;
  assign new_n40389_ = ~\b[29]  & ~new_n40388_;
  assign new_n40390_ = ~new_n39849_ & ~new_n40281_;
  assign new_n40391_ = ~new_n39859_ & new_n40213_;
  assign new_n40392_ = ~new_n40209_ & new_n40391_;
  assign new_n40393_ = ~new_n40210_ & ~new_n40213_;
  assign new_n40394_ = ~new_n40392_ & ~new_n40393_;
  assign new_n40395_ = new_n12184_ & ~new_n40394_;
  assign new_n40396_ = ~new_n40280_ & new_n40395_;
  assign new_n40397_ = ~new_n40390_ & ~new_n40396_;
  assign new_n40398_ = ~\b[28]  & ~new_n40397_;
  assign new_n40399_ = ~new_n39858_ & ~new_n40281_;
  assign new_n40400_ = ~new_n39868_ & new_n40208_;
  assign new_n40401_ = ~new_n40204_ & new_n40400_;
  assign new_n40402_ = ~new_n40205_ & ~new_n40208_;
  assign new_n40403_ = ~new_n40401_ & ~new_n40402_;
  assign new_n40404_ = new_n12184_ & ~new_n40403_;
  assign new_n40405_ = ~new_n40280_ & new_n40404_;
  assign new_n40406_ = ~new_n40399_ & ~new_n40405_;
  assign new_n40407_ = ~\b[27]  & ~new_n40406_;
  assign new_n40408_ = ~new_n39867_ & ~new_n40281_;
  assign new_n40409_ = ~new_n39877_ & new_n40203_;
  assign new_n40410_ = ~new_n40199_ & new_n40409_;
  assign new_n40411_ = ~new_n40200_ & ~new_n40203_;
  assign new_n40412_ = ~new_n40410_ & ~new_n40411_;
  assign new_n40413_ = new_n12184_ & ~new_n40412_;
  assign new_n40414_ = ~new_n40280_ & new_n40413_;
  assign new_n40415_ = ~new_n40408_ & ~new_n40414_;
  assign new_n40416_ = ~\b[26]  & ~new_n40415_;
  assign new_n40417_ = ~new_n39876_ & ~new_n40281_;
  assign new_n40418_ = ~new_n39886_ & new_n40198_;
  assign new_n40419_ = ~new_n40194_ & new_n40418_;
  assign new_n40420_ = ~new_n40195_ & ~new_n40198_;
  assign new_n40421_ = ~new_n40419_ & ~new_n40420_;
  assign new_n40422_ = new_n12184_ & ~new_n40421_;
  assign new_n40423_ = ~new_n40280_ & new_n40422_;
  assign new_n40424_ = ~new_n40417_ & ~new_n40423_;
  assign new_n40425_ = ~\b[25]  & ~new_n40424_;
  assign new_n40426_ = ~new_n39885_ & ~new_n40281_;
  assign new_n40427_ = ~new_n39895_ & new_n40193_;
  assign new_n40428_ = ~new_n40189_ & new_n40427_;
  assign new_n40429_ = ~new_n40190_ & ~new_n40193_;
  assign new_n40430_ = ~new_n40428_ & ~new_n40429_;
  assign new_n40431_ = new_n12184_ & ~new_n40430_;
  assign new_n40432_ = ~new_n40280_ & new_n40431_;
  assign new_n40433_ = ~new_n40426_ & ~new_n40432_;
  assign new_n40434_ = ~\b[24]  & ~new_n40433_;
  assign new_n40435_ = ~new_n39894_ & ~new_n40281_;
  assign new_n40436_ = ~new_n39904_ & new_n40188_;
  assign new_n40437_ = ~new_n40184_ & new_n40436_;
  assign new_n40438_ = ~new_n40185_ & ~new_n40188_;
  assign new_n40439_ = ~new_n40437_ & ~new_n40438_;
  assign new_n40440_ = new_n12184_ & ~new_n40439_;
  assign new_n40441_ = ~new_n40280_ & new_n40440_;
  assign new_n40442_ = ~new_n40435_ & ~new_n40441_;
  assign new_n40443_ = ~\b[23]  & ~new_n40442_;
  assign new_n40444_ = ~new_n39903_ & ~new_n40281_;
  assign new_n40445_ = ~new_n39913_ & new_n40183_;
  assign new_n40446_ = ~new_n40179_ & new_n40445_;
  assign new_n40447_ = ~new_n40180_ & ~new_n40183_;
  assign new_n40448_ = ~new_n40446_ & ~new_n40447_;
  assign new_n40449_ = new_n12184_ & ~new_n40448_;
  assign new_n40450_ = ~new_n40280_ & new_n40449_;
  assign new_n40451_ = ~new_n40444_ & ~new_n40450_;
  assign new_n40452_ = ~\b[22]  & ~new_n40451_;
  assign new_n40453_ = ~new_n39912_ & ~new_n40281_;
  assign new_n40454_ = ~new_n39922_ & new_n40178_;
  assign new_n40455_ = ~new_n40174_ & new_n40454_;
  assign new_n40456_ = ~new_n40175_ & ~new_n40178_;
  assign new_n40457_ = ~new_n40455_ & ~new_n40456_;
  assign new_n40458_ = new_n12184_ & ~new_n40457_;
  assign new_n40459_ = ~new_n40280_ & new_n40458_;
  assign new_n40460_ = ~new_n40453_ & ~new_n40459_;
  assign new_n40461_ = ~\b[21]  & ~new_n40460_;
  assign new_n40462_ = ~new_n39921_ & ~new_n40281_;
  assign new_n40463_ = ~new_n39931_ & new_n40173_;
  assign new_n40464_ = ~new_n40169_ & new_n40463_;
  assign new_n40465_ = ~new_n40170_ & ~new_n40173_;
  assign new_n40466_ = ~new_n40464_ & ~new_n40465_;
  assign new_n40467_ = new_n12184_ & ~new_n40466_;
  assign new_n40468_ = ~new_n40280_ & new_n40467_;
  assign new_n40469_ = ~new_n40462_ & ~new_n40468_;
  assign new_n40470_ = ~\b[20]  & ~new_n40469_;
  assign new_n40471_ = ~new_n39930_ & ~new_n40281_;
  assign new_n40472_ = ~new_n39940_ & new_n40168_;
  assign new_n40473_ = ~new_n40164_ & new_n40472_;
  assign new_n40474_ = ~new_n40165_ & ~new_n40168_;
  assign new_n40475_ = ~new_n40473_ & ~new_n40474_;
  assign new_n40476_ = new_n12184_ & ~new_n40475_;
  assign new_n40477_ = ~new_n40280_ & new_n40476_;
  assign new_n40478_ = ~new_n40471_ & ~new_n40477_;
  assign new_n40479_ = ~\b[19]  & ~new_n40478_;
  assign new_n40480_ = ~new_n39939_ & ~new_n40281_;
  assign new_n40481_ = ~new_n39949_ & new_n40163_;
  assign new_n40482_ = ~new_n40159_ & new_n40481_;
  assign new_n40483_ = ~new_n40160_ & ~new_n40163_;
  assign new_n40484_ = ~new_n40482_ & ~new_n40483_;
  assign new_n40485_ = new_n12184_ & ~new_n40484_;
  assign new_n40486_ = ~new_n40280_ & new_n40485_;
  assign new_n40487_ = ~new_n40480_ & ~new_n40486_;
  assign new_n40488_ = ~\b[18]  & ~new_n40487_;
  assign new_n40489_ = ~new_n39948_ & ~new_n40281_;
  assign new_n40490_ = ~new_n39958_ & new_n40158_;
  assign new_n40491_ = ~new_n40154_ & new_n40490_;
  assign new_n40492_ = ~new_n40155_ & ~new_n40158_;
  assign new_n40493_ = ~new_n40491_ & ~new_n40492_;
  assign new_n40494_ = new_n12184_ & ~new_n40493_;
  assign new_n40495_ = ~new_n40280_ & new_n40494_;
  assign new_n40496_ = ~new_n40489_ & ~new_n40495_;
  assign new_n40497_ = ~\b[17]  & ~new_n40496_;
  assign new_n40498_ = ~new_n39957_ & ~new_n40281_;
  assign new_n40499_ = ~new_n39967_ & new_n40153_;
  assign new_n40500_ = ~new_n40149_ & new_n40499_;
  assign new_n40501_ = ~new_n40150_ & ~new_n40153_;
  assign new_n40502_ = ~new_n40500_ & ~new_n40501_;
  assign new_n40503_ = new_n12184_ & ~new_n40502_;
  assign new_n40504_ = ~new_n40280_ & new_n40503_;
  assign new_n40505_ = ~new_n40498_ & ~new_n40504_;
  assign new_n40506_ = ~\b[16]  & ~new_n40505_;
  assign new_n40507_ = ~new_n39966_ & ~new_n40281_;
  assign new_n40508_ = ~new_n39976_ & new_n40148_;
  assign new_n40509_ = ~new_n40144_ & new_n40508_;
  assign new_n40510_ = ~new_n40145_ & ~new_n40148_;
  assign new_n40511_ = ~new_n40509_ & ~new_n40510_;
  assign new_n40512_ = new_n12184_ & ~new_n40511_;
  assign new_n40513_ = ~new_n40280_ & new_n40512_;
  assign new_n40514_ = ~new_n40507_ & ~new_n40513_;
  assign new_n40515_ = ~\b[15]  & ~new_n40514_;
  assign new_n40516_ = ~new_n39975_ & ~new_n40281_;
  assign new_n40517_ = ~new_n39985_ & new_n40143_;
  assign new_n40518_ = ~new_n40139_ & new_n40517_;
  assign new_n40519_ = ~new_n40140_ & ~new_n40143_;
  assign new_n40520_ = ~new_n40518_ & ~new_n40519_;
  assign new_n40521_ = new_n12184_ & ~new_n40520_;
  assign new_n40522_ = ~new_n40280_ & new_n40521_;
  assign new_n40523_ = ~new_n40516_ & ~new_n40522_;
  assign new_n40524_ = ~\b[14]  & ~new_n40523_;
  assign new_n40525_ = ~new_n39984_ & ~new_n40281_;
  assign new_n40526_ = ~new_n39994_ & new_n40138_;
  assign new_n40527_ = ~new_n40134_ & new_n40526_;
  assign new_n40528_ = ~new_n40135_ & ~new_n40138_;
  assign new_n40529_ = ~new_n40527_ & ~new_n40528_;
  assign new_n40530_ = new_n12184_ & ~new_n40529_;
  assign new_n40531_ = ~new_n40280_ & new_n40530_;
  assign new_n40532_ = ~new_n40525_ & ~new_n40531_;
  assign new_n40533_ = ~\b[13]  & ~new_n40532_;
  assign new_n40534_ = ~new_n39993_ & ~new_n40281_;
  assign new_n40535_ = ~new_n40003_ & new_n40133_;
  assign new_n40536_ = ~new_n40129_ & new_n40535_;
  assign new_n40537_ = ~new_n40130_ & ~new_n40133_;
  assign new_n40538_ = ~new_n40536_ & ~new_n40537_;
  assign new_n40539_ = new_n12184_ & ~new_n40538_;
  assign new_n40540_ = ~new_n40280_ & new_n40539_;
  assign new_n40541_ = ~new_n40534_ & ~new_n40540_;
  assign new_n40542_ = ~\b[12]  & ~new_n40541_;
  assign new_n40543_ = ~new_n40002_ & ~new_n40281_;
  assign new_n40544_ = ~new_n40012_ & new_n40128_;
  assign new_n40545_ = ~new_n40124_ & new_n40544_;
  assign new_n40546_ = ~new_n40125_ & ~new_n40128_;
  assign new_n40547_ = ~new_n40545_ & ~new_n40546_;
  assign new_n40548_ = new_n12184_ & ~new_n40547_;
  assign new_n40549_ = ~new_n40280_ & new_n40548_;
  assign new_n40550_ = ~new_n40543_ & ~new_n40549_;
  assign new_n40551_ = ~\b[11]  & ~new_n40550_;
  assign new_n40552_ = ~new_n40011_ & ~new_n40281_;
  assign new_n40553_ = ~new_n40021_ & new_n40123_;
  assign new_n40554_ = ~new_n40119_ & new_n40553_;
  assign new_n40555_ = ~new_n40120_ & ~new_n40123_;
  assign new_n40556_ = ~new_n40554_ & ~new_n40555_;
  assign new_n40557_ = new_n12184_ & ~new_n40556_;
  assign new_n40558_ = ~new_n40280_ & new_n40557_;
  assign new_n40559_ = ~new_n40552_ & ~new_n40558_;
  assign new_n40560_ = ~\b[10]  & ~new_n40559_;
  assign new_n40561_ = ~new_n40020_ & ~new_n40281_;
  assign new_n40562_ = ~new_n40030_ & new_n40118_;
  assign new_n40563_ = ~new_n40114_ & new_n40562_;
  assign new_n40564_ = ~new_n40115_ & ~new_n40118_;
  assign new_n40565_ = ~new_n40563_ & ~new_n40564_;
  assign new_n40566_ = new_n12184_ & ~new_n40565_;
  assign new_n40567_ = ~new_n40280_ & new_n40566_;
  assign new_n40568_ = ~new_n40561_ & ~new_n40567_;
  assign new_n40569_ = ~\b[9]  & ~new_n40568_;
  assign new_n40570_ = ~new_n40029_ & ~new_n40281_;
  assign new_n40571_ = ~new_n40039_ & new_n40113_;
  assign new_n40572_ = ~new_n40109_ & new_n40571_;
  assign new_n40573_ = ~new_n40110_ & ~new_n40113_;
  assign new_n40574_ = ~new_n40572_ & ~new_n40573_;
  assign new_n40575_ = new_n12184_ & ~new_n40574_;
  assign new_n40576_ = ~new_n40280_ & new_n40575_;
  assign new_n40577_ = ~new_n40570_ & ~new_n40576_;
  assign new_n40578_ = ~\b[8]  & ~new_n40577_;
  assign new_n40579_ = ~new_n40038_ & ~new_n40281_;
  assign new_n40580_ = ~new_n40048_ & new_n40108_;
  assign new_n40581_ = ~new_n40104_ & new_n40580_;
  assign new_n40582_ = ~new_n40105_ & ~new_n40108_;
  assign new_n40583_ = ~new_n40581_ & ~new_n40582_;
  assign new_n40584_ = new_n12184_ & ~new_n40583_;
  assign new_n40585_ = ~new_n40280_ & new_n40584_;
  assign new_n40586_ = ~new_n40579_ & ~new_n40585_;
  assign new_n40587_ = ~\b[7]  & ~new_n40586_;
  assign new_n40588_ = ~new_n40047_ & ~new_n40281_;
  assign new_n40589_ = ~new_n40057_ & new_n40103_;
  assign new_n40590_ = ~new_n40099_ & new_n40589_;
  assign new_n40591_ = ~new_n40100_ & ~new_n40103_;
  assign new_n40592_ = ~new_n40590_ & ~new_n40591_;
  assign new_n40593_ = new_n12184_ & ~new_n40592_;
  assign new_n40594_ = ~new_n40280_ & new_n40593_;
  assign new_n40595_ = ~new_n40588_ & ~new_n40594_;
  assign new_n40596_ = ~\b[6]  & ~new_n40595_;
  assign new_n40597_ = ~new_n40056_ & ~new_n40281_;
  assign new_n40598_ = ~new_n40066_ & new_n40098_;
  assign new_n40599_ = ~new_n40094_ & new_n40598_;
  assign new_n40600_ = ~new_n40095_ & ~new_n40098_;
  assign new_n40601_ = ~new_n40599_ & ~new_n40600_;
  assign new_n40602_ = new_n12184_ & ~new_n40601_;
  assign new_n40603_ = ~new_n40280_ & new_n40602_;
  assign new_n40604_ = ~new_n40597_ & ~new_n40603_;
  assign new_n40605_ = ~\b[5]  & ~new_n40604_;
  assign new_n40606_ = ~new_n40065_ & ~new_n40281_;
  assign new_n40607_ = ~new_n40074_ & new_n40093_;
  assign new_n40608_ = ~new_n40089_ & new_n40607_;
  assign new_n40609_ = ~new_n40090_ & ~new_n40093_;
  assign new_n40610_ = ~new_n40608_ & ~new_n40609_;
  assign new_n40611_ = new_n12184_ & ~new_n40610_;
  assign new_n40612_ = ~new_n40280_ & new_n40611_;
  assign new_n40613_ = ~new_n40606_ & ~new_n40612_;
  assign new_n40614_ = ~\b[4]  & ~new_n40613_;
  assign new_n40615_ = ~new_n40073_ & ~new_n40281_;
  assign new_n40616_ = ~new_n40084_ & new_n40088_;
  assign new_n40617_ = ~new_n40083_ & new_n40616_;
  assign new_n40618_ = ~new_n40085_ & ~new_n40088_;
  assign new_n40619_ = ~new_n40617_ & ~new_n40618_;
  assign new_n40620_ = new_n12184_ & ~new_n40619_;
  assign new_n40621_ = ~new_n40280_ & new_n40620_;
  assign new_n40622_ = ~new_n40615_ & ~new_n40621_;
  assign new_n40623_ = ~\b[3]  & ~new_n40622_;
  assign new_n40624_ = ~new_n40078_ & ~new_n40281_;
  assign new_n40625_ = new_n11985_ & ~new_n40081_;
  assign new_n40626_ = ~new_n40079_ & new_n40625_;
  assign new_n40627_ = new_n12184_ & ~new_n40626_;
  assign new_n40628_ = ~new_n40083_ & new_n40627_;
  assign new_n40629_ = ~new_n40280_ & new_n40628_;
  assign new_n40630_ = ~new_n40624_ & ~new_n40629_;
  assign new_n40631_ = ~\b[2]  & ~new_n40630_;
  assign new_n40632_ = new_n12539_ & ~new_n40280_;
  assign new_n40633_ = \a[23]  & ~new_n40632_;
  assign new_n40634_ = new_n12544_ & ~new_n40280_;
  assign new_n40635_ = ~new_n40633_ & ~new_n40634_;
  assign new_n40636_ = \b[1]  & ~new_n40635_;
  assign new_n40637_ = ~\b[1]  & ~new_n40634_;
  assign new_n40638_ = ~new_n40633_ & new_n40637_;
  assign new_n40639_ = ~new_n40636_ & ~new_n40638_;
  assign new_n40640_ = ~new_n12551_ & ~new_n40639_;
  assign new_n40641_ = ~\b[1]  & ~new_n40635_;
  assign new_n40642_ = ~new_n40640_ & ~new_n40641_;
  assign new_n40643_ = \b[2]  & ~new_n40629_;
  assign new_n40644_ = ~new_n40624_ & new_n40643_;
  assign new_n40645_ = ~new_n40631_ & ~new_n40644_;
  assign new_n40646_ = ~new_n40642_ & new_n40645_;
  assign new_n40647_ = ~new_n40631_ & ~new_n40646_;
  assign new_n40648_ = \b[3]  & ~new_n40621_;
  assign new_n40649_ = ~new_n40615_ & new_n40648_;
  assign new_n40650_ = ~new_n40623_ & ~new_n40649_;
  assign new_n40651_ = ~new_n40647_ & new_n40650_;
  assign new_n40652_ = ~new_n40623_ & ~new_n40651_;
  assign new_n40653_ = \b[4]  & ~new_n40612_;
  assign new_n40654_ = ~new_n40606_ & new_n40653_;
  assign new_n40655_ = ~new_n40614_ & ~new_n40654_;
  assign new_n40656_ = ~new_n40652_ & new_n40655_;
  assign new_n40657_ = ~new_n40614_ & ~new_n40656_;
  assign new_n40658_ = \b[5]  & ~new_n40603_;
  assign new_n40659_ = ~new_n40597_ & new_n40658_;
  assign new_n40660_ = ~new_n40605_ & ~new_n40659_;
  assign new_n40661_ = ~new_n40657_ & new_n40660_;
  assign new_n40662_ = ~new_n40605_ & ~new_n40661_;
  assign new_n40663_ = \b[6]  & ~new_n40594_;
  assign new_n40664_ = ~new_n40588_ & new_n40663_;
  assign new_n40665_ = ~new_n40596_ & ~new_n40664_;
  assign new_n40666_ = ~new_n40662_ & new_n40665_;
  assign new_n40667_ = ~new_n40596_ & ~new_n40666_;
  assign new_n40668_ = \b[7]  & ~new_n40585_;
  assign new_n40669_ = ~new_n40579_ & new_n40668_;
  assign new_n40670_ = ~new_n40587_ & ~new_n40669_;
  assign new_n40671_ = ~new_n40667_ & new_n40670_;
  assign new_n40672_ = ~new_n40587_ & ~new_n40671_;
  assign new_n40673_ = \b[8]  & ~new_n40576_;
  assign new_n40674_ = ~new_n40570_ & new_n40673_;
  assign new_n40675_ = ~new_n40578_ & ~new_n40674_;
  assign new_n40676_ = ~new_n40672_ & new_n40675_;
  assign new_n40677_ = ~new_n40578_ & ~new_n40676_;
  assign new_n40678_ = \b[9]  & ~new_n40567_;
  assign new_n40679_ = ~new_n40561_ & new_n40678_;
  assign new_n40680_ = ~new_n40569_ & ~new_n40679_;
  assign new_n40681_ = ~new_n40677_ & new_n40680_;
  assign new_n40682_ = ~new_n40569_ & ~new_n40681_;
  assign new_n40683_ = \b[10]  & ~new_n40558_;
  assign new_n40684_ = ~new_n40552_ & new_n40683_;
  assign new_n40685_ = ~new_n40560_ & ~new_n40684_;
  assign new_n40686_ = ~new_n40682_ & new_n40685_;
  assign new_n40687_ = ~new_n40560_ & ~new_n40686_;
  assign new_n40688_ = \b[11]  & ~new_n40549_;
  assign new_n40689_ = ~new_n40543_ & new_n40688_;
  assign new_n40690_ = ~new_n40551_ & ~new_n40689_;
  assign new_n40691_ = ~new_n40687_ & new_n40690_;
  assign new_n40692_ = ~new_n40551_ & ~new_n40691_;
  assign new_n40693_ = \b[12]  & ~new_n40540_;
  assign new_n40694_ = ~new_n40534_ & new_n40693_;
  assign new_n40695_ = ~new_n40542_ & ~new_n40694_;
  assign new_n40696_ = ~new_n40692_ & new_n40695_;
  assign new_n40697_ = ~new_n40542_ & ~new_n40696_;
  assign new_n40698_ = \b[13]  & ~new_n40531_;
  assign new_n40699_ = ~new_n40525_ & new_n40698_;
  assign new_n40700_ = ~new_n40533_ & ~new_n40699_;
  assign new_n40701_ = ~new_n40697_ & new_n40700_;
  assign new_n40702_ = ~new_n40533_ & ~new_n40701_;
  assign new_n40703_ = \b[14]  & ~new_n40522_;
  assign new_n40704_ = ~new_n40516_ & new_n40703_;
  assign new_n40705_ = ~new_n40524_ & ~new_n40704_;
  assign new_n40706_ = ~new_n40702_ & new_n40705_;
  assign new_n40707_ = ~new_n40524_ & ~new_n40706_;
  assign new_n40708_ = \b[15]  & ~new_n40513_;
  assign new_n40709_ = ~new_n40507_ & new_n40708_;
  assign new_n40710_ = ~new_n40515_ & ~new_n40709_;
  assign new_n40711_ = ~new_n40707_ & new_n40710_;
  assign new_n40712_ = ~new_n40515_ & ~new_n40711_;
  assign new_n40713_ = \b[16]  & ~new_n40504_;
  assign new_n40714_ = ~new_n40498_ & new_n40713_;
  assign new_n40715_ = ~new_n40506_ & ~new_n40714_;
  assign new_n40716_ = ~new_n40712_ & new_n40715_;
  assign new_n40717_ = ~new_n40506_ & ~new_n40716_;
  assign new_n40718_ = \b[17]  & ~new_n40495_;
  assign new_n40719_ = ~new_n40489_ & new_n40718_;
  assign new_n40720_ = ~new_n40497_ & ~new_n40719_;
  assign new_n40721_ = ~new_n40717_ & new_n40720_;
  assign new_n40722_ = ~new_n40497_ & ~new_n40721_;
  assign new_n40723_ = \b[18]  & ~new_n40486_;
  assign new_n40724_ = ~new_n40480_ & new_n40723_;
  assign new_n40725_ = ~new_n40488_ & ~new_n40724_;
  assign new_n40726_ = ~new_n40722_ & new_n40725_;
  assign new_n40727_ = ~new_n40488_ & ~new_n40726_;
  assign new_n40728_ = \b[19]  & ~new_n40477_;
  assign new_n40729_ = ~new_n40471_ & new_n40728_;
  assign new_n40730_ = ~new_n40479_ & ~new_n40729_;
  assign new_n40731_ = ~new_n40727_ & new_n40730_;
  assign new_n40732_ = ~new_n40479_ & ~new_n40731_;
  assign new_n40733_ = \b[20]  & ~new_n40468_;
  assign new_n40734_ = ~new_n40462_ & new_n40733_;
  assign new_n40735_ = ~new_n40470_ & ~new_n40734_;
  assign new_n40736_ = ~new_n40732_ & new_n40735_;
  assign new_n40737_ = ~new_n40470_ & ~new_n40736_;
  assign new_n40738_ = \b[21]  & ~new_n40459_;
  assign new_n40739_ = ~new_n40453_ & new_n40738_;
  assign new_n40740_ = ~new_n40461_ & ~new_n40739_;
  assign new_n40741_ = ~new_n40737_ & new_n40740_;
  assign new_n40742_ = ~new_n40461_ & ~new_n40741_;
  assign new_n40743_ = \b[22]  & ~new_n40450_;
  assign new_n40744_ = ~new_n40444_ & new_n40743_;
  assign new_n40745_ = ~new_n40452_ & ~new_n40744_;
  assign new_n40746_ = ~new_n40742_ & new_n40745_;
  assign new_n40747_ = ~new_n40452_ & ~new_n40746_;
  assign new_n40748_ = \b[23]  & ~new_n40441_;
  assign new_n40749_ = ~new_n40435_ & new_n40748_;
  assign new_n40750_ = ~new_n40443_ & ~new_n40749_;
  assign new_n40751_ = ~new_n40747_ & new_n40750_;
  assign new_n40752_ = ~new_n40443_ & ~new_n40751_;
  assign new_n40753_ = \b[24]  & ~new_n40432_;
  assign new_n40754_ = ~new_n40426_ & new_n40753_;
  assign new_n40755_ = ~new_n40434_ & ~new_n40754_;
  assign new_n40756_ = ~new_n40752_ & new_n40755_;
  assign new_n40757_ = ~new_n40434_ & ~new_n40756_;
  assign new_n40758_ = \b[25]  & ~new_n40423_;
  assign new_n40759_ = ~new_n40417_ & new_n40758_;
  assign new_n40760_ = ~new_n40425_ & ~new_n40759_;
  assign new_n40761_ = ~new_n40757_ & new_n40760_;
  assign new_n40762_ = ~new_n40425_ & ~new_n40761_;
  assign new_n40763_ = \b[26]  & ~new_n40414_;
  assign new_n40764_ = ~new_n40408_ & new_n40763_;
  assign new_n40765_ = ~new_n40416_ & ~new_n40764_;
  assign new_n40766_ = ~new_n40762_ & new_n40765_;
  assign new_n40767_ = ~new_n40416_ & ~new_n40766_;
  assign new_n40768_ = \b[27]  & ~new_n40405_;
  assign new_n40769_ = ~new_n40399_ & new_n40768_;
  assign new_n40770_ = ~new_n40407_ & ~new_n40769_;
  assign new_n40771_ = ~new_n40767_ & new_n40770_;
  assign new_n40772_ = ~new_n40407_ & ~new_n40771_;
  assign new_n40773_ = \b[28]  & ~new_n40396_;
  assign new_n40774_ = ~new_n40390_ & new_n40773_;
  assign new_n40775_ = ~new_n40398_ & ~new_n40774_;
  assign new_n40776_ = ~new_n40772_ & new_n40775_;
  assign new_n40777_ = ~new_n40398_ & ~new_n40776_;
  assign new_n40778_ = \b[29]  & ~new_n40387_;
  assign new_n40779_ = ~new_n40381_ & new_n40778_;
  assign new_n40780_ = ~new_n40389_ & ~new_n40779_;
  assign new_n40781_ = ~new_n40777_ & new_n40780_;
  assign new_n40782_ = ~new_n40389_ & ~new_n40781_;
  assign new_n40783_ = \b[30]  & ~new_n40378_;
  assign new_n40784_ = ~new_n40372_ & new_n40783_;
  assign new_n40785_ = ~new_n40380_ & ~new_n40784_;
  assign new_n40786_ = ~new_n40782_ & new_n40785_;
  assign new_n40787_ = ~new_n40380_ & ~new_n40786_;
  assign new_n40788_ = \b[31]  & ~new_n40369_;
  assign new_n40789_ = ~new_n40363_ & new_n40788_;
  assign new_n40790_ = ~new_n40371_ & ~new_n40789_;
  assign new_n40791_ = ~new_n40787_ & new_n40790_;
  assign new_n40792_ = ~new_n40371_ & ~new_n40791_;
  assign new_n40793_ = \b[32]  & ~new_n40360_;
  assign new_n40794_ = ~new_n40354_ & new_n40793_;
  assign new_n40795_ = ~new_n40362_ & ~new_n40794_;
  assign new_n40796_ = ~new_n40792_ & new_n40795_;
  assign new_n40797_ = ~new_n40362_ & ~new_n40796_;
  assign new_n40798_ = \b[33]  & ~new_n40351_;
  assign new_n40799_ = ~new_n40345_ & new_n40798_;
  assign new_n40800_ = ~new_n40353_ & ~new_n40799_;
  assign new_n40801_ = ~new_n40797_ & new_n40800_;
  assign new_n40802_ = ~new_n40353_ & ~new_n40801_;
  assign new_n40803_ = \b[34]  & ~new_n40342_;
  assign new_n40804_ = ~new_n40336_ & new_n40803_;
  assign new_n40805_ = ~new_n40344_ & ~new_n40804_;
  assign new_n40806_ = ~new_n40802_ & new_n40805_;
  assign new_n40807_ = ~new_n40344_ & ~new_n40806_;
  assign new_n40808_ = \b[35]  & ~new_n40333_;
  assign new_n40809_ = ~new_n40327_ & new_n40808_;
  assign new_n40810_ = ~new_n40335_ & ~new_n40809_;
  assign new_n40811_ = ~new_n40807_ & new_n40810_;
  assign new_n40812_ = ~new_n40335_ & ~new_n40811_;
  assign new_n40813_ = \b[36]  & ~new_n40324_;
  assign new_n40814_ = ~new_n40318_ & new_n40813_;
  assign new_n40815_ = ~new_n40326_ & ~new_n40814_;
  assign new_n40816_ = ~new_n40812_ & new_n40815_;
  assign new_n40817_ = ~new_n40326_ & ~new_n40816_;
  assign new_n40818_ = \b[37]  & ~new_n40315_;
  assign new_n40819_ = ~new_n40309_ & new_n40818_;
  assign new_n40820_ = ~new_n40317_ & ~new_n40819_;
  assign new_n40821_ = ~new_n40817_ & new_n40820_;
  assign new_n40822_ = ~new_n40317_ & ~new_n40821_;
  assign new_n40823_ = \b[38]  & ~new_n40306_;
  assign new_n40824_ = ~new_n40300_ & new_n40823_;
  assign new_n40825_ = ~new_n40308_ & ~new_n40824_;
  assign new_n40826_ = ~new_n40822_ & new_n40825_;
  assign new_n40827_ = ~new_n40308_ & ~new_n40826_;
  assign new_n40828_ = \b[39]  & ~new_n40297_;
  assign new_n40829_ = ~new_n40291_ & new_n40828_;
  assign new_n40830_ = ~new_n40299_ & ~new_n40829_;
  assign new_n40831_ = ~new_n40827_ & new_n40830_;
  assign new_n40832_ = ~new_n40299_ & ~new_n40831_;
  assign new_n40833_ = \b[40]  & ~new_n40288_;
  assign new_n40834_ = ~new_n40282_ & new_n40833_;
  assign new_n40835_ = ~new_n40290_ & ~new_n40834_;
  assign new_n40836_ = ~new_n40832_ & new_n40835_;
  assign new_n40837_ = ~new_n40290_ & ~new_n40836_;
  assign new_n40838_ = ~new_n39740_ & ~new_n40281_;
  assign new_n40839_ = ~new_n39742_ & new_n40278_;
  assign new_n40840_ = ~new_n40274_ & new_n40839_;
  assign new_n40841_ = ~new_n40275_ & ~new_n40278_;
  assign new_n40842_ = ~new_n40840_ & ~new_n40841_;
  assign new_n40843_ = new_n40281_ & ~new_n40842_;
  assign new_n40844_ = ~new_n40838_ & ~new_n40843_;
  assign new_n40845_ = ~\b[41]  & ~new_n40844_;
  assign new_n40846_ = \b[41]  & ~new_n40838_;
  assign new_n40847_ = ~new_n40843_ & new_n40846_;
  assign new_n40848_ = new_n12761_ & ~new_n40847_;
  assign new_n40849_ = ~new_n40845_ & new_n40848_;
  assign new_n40850_ = ~new_n40837_ & new_n40849_;
  assign new_n40851_ = new_n12184_ & ~new_n40844_;
  assign new_n40852_ = ~new_n40850_ & ~new_n40851_;
  assign new_n40853_ = ~new_n40299_ & new_n40835_;
  assign new_n40854_ = ~new_n40831_ & new_n40853_;
  assign new_n40855_ = ~new_n40832_ & ~new_n40835_;
  assign new_n40856_ = ~new_n40854_ & ~new_n40855_;
  assign new_n40857_ = ~new_n40852_ & ~new_n40856_;
  assign new_n40858_ = ~new_n40289_ & ~new_n40851_;
  assign new_n40859_ = ~new_n40850_ & new_n40858_;
  assign new_n40860_ = ~new_n40857_ & ~new_n40859_;
  assign new_n40861_ = ~new_n40290_ & ~new_n40847_;
  assign new_n40862_ = ~new_n40845_ & new_n40861_;
  assign new_n40863_ = ~new_n40836_ & new_n40862_;
  assign new_n40864_ = ~new_n40845_ & ~new_n40847_;
  assign new_n40865_ = ~new_n40837_ & ~new_n40864_;
  assign new_n40866_ = ~new_n40863_ & ~new_n40865_;
  assign new_n40867_ = ~new_n40852_ & ~new_n40866_;
  assign new_n40868_ = ~new_n40844_ & ~new_n40851_;
  assign new_n40869_ = ~new_n40850_ & new_n40868_;
  assign new_n40870_ = ~new_n40867_ & ~new_n40869_;
  assign new_n40871_ = ~\b[42]  & ~new_n40870_;
  assign new_n40872_ = ~\b[41]  & ~new_n40860_;
  assign new_n40873_ = ~new_n40308_ & new_n40830_;
  assign new_n40874_ = ~new_n40826_ & new_n40873_;
  assign new_n40875_ = ~new_n40827_ & ~new_n40830_;
  assign new_n40876_ = ~new_n40874_ & ~new_n40875_;
  assign new_n40877_ = ~new_n40852_ & ~new_n40876_;
  assign new_n40878_ = ~new_n40298_ & ~new_n40851_;
  assign new_n40879_ = ~new_n40850_ & new_n40878_;
  assign new_n40880_ = ~new_n40877_ & ~new_n40879_;
  assign new_n40881_ = ~\b[40]  & ~new_n40880_;
  assign new_n40882_ = ~new_n40317_ & new_n40825_;
  assign new_n40883_ = ~new_n40821_ & new_n40882_;
  assign new_n40884_ = ~new_n40822_ & ~new_n40825_;
  assign new_n40885_ = ~new_n40883_ & ~new_n40884_;
  assign new_n40886_ = ~new_n40852_ & ~new_n40885_;
  assign new_n40887_ = ~new_n40307_ & ~new_n40851_;
  assign new_n40888_ = ~new_n40850_ & new_n40887_;
  assign new_n40889_ = ~new_n40886_ & ~new_n40888_;
  assign new_n40890_ = ~\b[39]  & ~new_n40889_;
  assign new_n40891_ = ~new_n40326_ & new_n40820_;
  assign new_n40892_ = ~new_n40816_ & new_n40891_;
  assign new_n40893_ = ~new_n40817_ & ~new_n40820_;
  assign new_n40894_ = ~new_n40892_ & ~new_n40893_;
  assign new_n40895_ = ~new_n40852_ & ~new_n40894_;
  assign new_n40896_ = ~new_n40316_ & ~new_n40851_;
  assign new_n40897_ = ~new_n40850_ & new_n40896_;
  assign new_n40898_ = ~new_n40895_ & ~new_n40897_;
  assign new_n40899_ = ~\b[38]  & ~new_n40898_;
  assign new_n40900_ = ~new_n40335_ & new_n40815_;
  assign new_n40901_ = ~new_n40811_ & new_n40900_;
  assign new_n40902_ = ~new_n40812_ & ~new_n40815_;
  assign new_n40903_ = ~new_n40901_ & ~new_n40902_;
  assign new_n40904_ = ~new_n40852_ & ~new_n40903_;
  assign new_n40905_ = ~new_n40325_ & ~new_n40851_;
  assign new_n40906_ = ~new_n40850_ & new_n40905_;
  assign new_n40907_ = ~new_n40904_ & ~new_n40906_;
  assign new_n40908_ = ~\b[37]  & ~new_n40907_;
  assign new_n40909_ = ~new_n40344_ & new_n40810_;
  assign new_n40910_ = ~new_n40806_ & new_n40909_;
  assign new_n40911_ = ~new_n40807_ & ~new_n40810_;
  assign new_n40912_ = ~new_n40910_ & ~new_n40911_;
  assign new_n40913_ = ~new_n40852_ & ~new_n40912_;
  assign new_n40914_ = ~new_n40334_ & ~new_n40851_;
  assign new_n40915_ = ~new_n40850_ & new_n40914_;
  assign new_n40916_ = ~new_n40913_ & ~new_n40915_;
  assign new_n40917_ = ~\b[36]  & ~new_n40916_;
  assign new_n40918_ = ~new_n40353_ & new_n40805_;
  assign new_n40919_ = ~new_n40801_ & new_n40918_;
  assign new_n40920_ = ~new_n40802_ & ~new_n40805_;
  assign new_n40921_ = ~new_n40919_ & ~new_n40920_;
  assign new_n40922_ = ~new_n40852_ & ~new_n40921_;
  assign new_n40923_ = ~new_n40343_ & ~new_n40851_;
  assign new_n40924_ = ~new_n40850_ & new_n40923_;
  assign new_n40925_ = ~new_n40922_ & ~new_n40924_;
  assign new_n40926_ = ~\b[35]  & ~new_n40925_;
  assign new_n40927_ = ~new_n40362_ & new_n40800_;
  assign new_n40928_ = ~new_n40796_ & new_n40927_;
  assign new_n40929_ = ~new_n40797_ & ~new_n40800_;
  assign new_n40930_ = ~new_n40928_ & ~new_n40929_;
  assign new_n40931_ = ~new_n40852_ & ~new_n40930_;
  assign new_n40932_ = ~new_n40352_ & ~new_n40851_;
  assign new_n40933_ = ~new_n40850_ & new_n40932_;
  assign new_n40934_ = ~new_n40931_ & ~new_n40933_;
  assign new_n40935_ = ~\b[34]  & ~new_n40934_;
  assign new_n40936_ = ~new_n40371_ & new_n40795_;
  assign new_n40937_ = ~new_n40791_ & new_n40936_;
  assign new_n40938_ = ~new_n40792_ & ~new_n40795_;
  assign new_n40939_ = ~new_n40937_ & ~new_n40938_;
  assign new_n40940_ = ~new_n40852_ & ~new_n40939_;
  assign new_n40941_ = ~new_n40361_ & ~new_n40851_;
  assign new_n40942_ = ~new_n40850_ & new_n40941_;
  assign new_n40943_ = ~new_n40940_ & ~new_n40942_;
  assign new_n40944_ = ~\b[33]  & ~new_n40943_;
  assign new_n40945_ = ~new_n40380_ & new_n40790_;
  assign new_n40946_ = ~new_n40786_ & new_n40945_;
  assign new_n40947_ = ~new_n40787_ & ~new_n40790_;
  assign new_n40948_ = ~new_n40946_ & ~new_n40947_;
  assign new_n40949_ = ~new_n40852_ & ~new_n40948_;
  assign new_n40950_ = ~new_n40370_ & ~new_n40851_;
  assign new_n40951_ = ~new_n40850_ & new_n40950_;
  assign new_n40952_ = ~new_n40949_ & ~new_n40951_;
  assign new_n40953_ = ~\b[32]  & ~new_n40952_;
  assign new_n40954_ = ~new_n40389_ & new_n40785_;
  assign new_n40955_ = ~new_n40781_ & new_n40954_;
  assign new_n40956_ = ~new_n40782_ & ~new_n40785_;
  assign new_n40957_ = ~new_n40955_ & ~new_n40956_;
  assign new_n40958_ = ~new_n40852_ & ~new_n40957_;
  assign new_n40959_ = ~new_n40379_ & ~new_n40851_;
  assign new_n40960_ = ~new_n40850_ & new_n40959_;
  assign new_n40961_ = ~new_n40958_ & ~new_n40960_;
  assign new_n40962_ = ~\b[31]  & ~new_n40961_;
  assign new_n40963_ = ~new_n40398_ & new_n40780_;
  assign new_n40964_ = ~new_n40776_ & new_n40963_;
  assign new_n40965_ = ~new_n40777_ & ~new_n40780_;
  assign new_n40966_ = ~new_n40964_ & ~new_n40965_;
  assign new_n40967_ = ~new_n40852_ & ~new_n40966_;
  assign new_n40968_ = ~new_n40388_ & ~new_n40851_;
  assign new_n40969_ = ~new_n40850_ & new_n40968_;
  assign new_n40970_ = ~new_n40967_ & ~new_n40969_;
  assign new_n40971_ = ~\b[30]  & ~new_n40970_;
  assign new_n40972_ = ~new_n40407_ & new_n40775_;
  assign new_n40973_ = ~new_n40771_ & new_n40972_;
  assign new_n40974_ = ~new_n40772_ & ~new_n40775_;
  assign new_n40975_ = ~new_n40973_ & ~new_n40974_;
  assign new_n40976_ = ~new_n40852_ & ~new_n40975_;
  assign new_n40977_ = ~new_n40397_ & ~new_n40851_;
  assign new_n40978_ = ~new_n40850_ & new_n40977_;
  assign new_n40979_ = ~new_n40976_ & ~new_n40978_;
  assign new_n40980_ = ~\b[29]  & ~new_n40979_;
  assign new_n40981_ = ~new_n40416_ & new_n40770_;
  assign new_n40982_ = ~new_n40766_ & new_n40981_;
  assign new_n40983_ = ~new_n40767_ & ~new_n40770_;
  assign new_n40984_ = ~new_n40982_ & ~new_n40983_;
  assign new_n40985_ = ~new_n40852_ & ~new_n40984_;
  assign new_n40986_ = ~new_n40406_ & ~new_n40851_;
  assign new_n40987_ = ~new_n40850_ & new_n40986_;
  assign new_n40988_ = ~new_n40985_ & ~new_n40987_;
  assign new_n40989_ = ~\b[28]  & ~new_n40988_;
  assign new_n40990_ = ~new_n40425_ & new_n40765_;
  assign new_n40991_ = ~new_n40761_ & new_n40990_;
  assign new_n40992_ = ~new_n40762_ & ~new_n40765_;
  assign new_n40993_ = ~new_n40991_ & ~new_n40992_;
  assign new_n40994_ = ~new_n40852_ & ~new_n40993_;
  assign new_n40995_ = ~new_n40415_ & ~new_n40851_;
  assign new_n40996_ = ~new_n40850_ & new_n40995_;
  assign new_n40997_ = ~new_n40994_ & ~new_n40996_;
  assign new_n40998_ = ~\b[27]  & ~new_n40997_;
  assign new_n40999_ = ~new_n40434_ & new_n40760_;
  assign new_n41000_ = ~new_n40756_ & new_n40999_;
  assign new_n41001_ = ~new_n40757_ & ~new_n40760_;
  assign new_n41002_ = ~new_n41000_ & ~new_n41001_;
  assign new_n41003_ = ~new_n40852_ & ~new_n41002_;
  assign new_n41004_ = ~new_n40424_ & ~new_n40851_;
  assign new_n41005_ = ~new_n40850_ & new_n41004_;
  assign new_n41006_ = ~new_n41003_ & ~new_n41005_;
  assign new_n41007_ = ~\b[26]  & ~new_n41006_;
  assign new_n41008_ = ~new_n40443_ & new_n40755_;
  assign new_n41009_ = ~new_n40751_ & new_n41008_;
  assign new_n41010_ = ~new_n40752_ & ~new_n40755_;
  assign new_n41011_ = ~new_n41009_ & ~new_n41010_;
  assign new_n41012_ = ~new_n40852_ & ~new_n41011_;
  assign new_n41013_ = ~new_n40433_ & ~new_n40851_;
  assign new_n41014_ = ~new_n40850_ & new_n41013_;
  assign new_n41015_ = ~new_n41012_ & ~new_n41014_;
  assign new_n41016_ = ~\b[25]  & ~new_n41015_;
  assign new_n41017_ = ~new_n40452_ & new_n40750_;
  assign new_n41018_ = ~new_n40746_ & new_n41017_;
  assign new_n41019_ = ~new_n40747_ & ~new_n40750_;
  assign new_n41020_ = ~new_n41018_ & ~new_n41019_;
  assign new_n41021_ = ~new_n40852_ & ~new_n41020_;
  assign new_n41022_ = ~new_n40442_ & ~new_n40851_;
  assign new_n41023_ = ~new_n40850_ & new_n41022_;
  assign new_n41024_ = ~new_n41021_ & ~new_n41023_;
  assign new_n41025_ = ~\b[24]  & ~new_n41024_;
  assign new_n41026_ = ~new_n40461_ & new_n40745_;
  assign new_n41027_ = ~new_n40741_ & new_n41026_;
  assign new_n41028_ = ~new_n40742_ & ~new_n40745_;
  assign new_n41029_ = ~new_n41027_ & ~new_n41028_;
  assign new_n41030_ = ~new_n40852_ & ~new_n41029_;
  assign new_n41031_ = ~new_n40451_ & ~new_n40851_;
  assign new_n41032_ = ~new_n40850_ & new_n41031_;
  assign new_n41033_ = ~new_n41030_ & ~new_n41032_;
  assign new_n41034_ = ~\b[23]  & ~new_n41033_;
  assign new_n41035_ = ~new_n40470_ & new_n40740_;
  assign new_n41036_ = ~new_n40736_ & new_n41035_;
  assign new_n41037_ = ~new_n40737_ & ~new_n40740_;
  assign new_n41038_ = ~new_n41036_ & ~new_n41037_;
  assign new_n41039_ = ~new_n40852_ & ~new_n41038_;
  assign new_n41040_ = ~new_n40460_ & ~new_n40851_;
  assign new_n41041_ = ~new_n40850_ & new_n41040_;
  assign new_n41042_ = ~new_n41039_ & ~new_n41041_;
  assign new_n41043_ = ~\b[22]  & ~new_n41042_;
  assign new_n41044_ = ~new_n40479_ & new_n40735_;
  assign new_n41045_ = ~new_n40731_ & new_n41044_;
  assign new_n41046_ = ~new_n40732_ & ~new_n40735_;
  assign new_n41047_ = ~new_n41045_ & ~new_n41046_;
  assign new_n41048_ = ~new_n40852_ & ~new_n41047_;
  assign new_n41049_ = ~new_n40469_ & ~new_n40851_;
  assign new_n41050_ = ~new_n40850_ & new_n41049_;
  assign new_n41051_ = ~new_n41048_ & ~new_n41050_;
  assign new_n41052_ = ~\b[21]  & ~new_n41051_;
  assign new_n41053_ = ~new_n40488_ & new_n40730_;
  assign new_n41054_ = ~new_n40726_ & new_n41053_;
  assign new_n41055_ = ~new_n40727_ & ~new_n40730_;
  assign new_n41056_ = ~new_n41054_ & ~new_n41055_;
  assign new_n41057_ = ~new_n40852_ & ~new_n41056_;
  assign new_n41058_ = ~new_n40478_ & ~new_n40851_;
  assign new_n41059_ = ~new_n40850_ & new_n41058_;
  assign new_n41060_ = ~new_n41057_ & ~new_n41059_;
  assign new_n41061_ = ~\b[20]  & ~new_n41060_;
  assign new_n41062_ = ~new_n40497_ & new_n40725_;
  assign new_n41063_ = ~new_n40721_ & new_n41062_;
  assign new_n41064_ = ~new_n40722_ & ~new_n40725_;
  assign new_n41065_ = ~new_n41063_ & ~new_n41064_;
  assign new_n41066_ = ~new_n40852_ & ~new_n41065_;
  assign new_n41067_ = ~new_n40487_ & ~new_n40851_;
  assign new_n41068_ = ~new_n40850_ & new_n41067_;
  assign new_n41069_ = ~new_n41066_ & ~new_n41068_;
  assign new_n41070_ = ~\b[19]  & ~new_n41069_;
  assign new_n41071_ = ~new_n40506_ & new_n40720_;
  assign new_n41072_ = ~new_n40716_ & new_n41071_;
  assign new_n41073_ = ~new_n40717_ & ~new_n40720_;
  assign new_n41074_ = ~new_n41072_ & ~new_n41073_;
  assign new_n41075_ = ~new_n40852_ & ~new_n41074_;
  assign new_n41076_ = ~new_n40496_ & ~new_n40851_;
  assign new_n41077_ = ~new_n40850_ & new_n41076_;
  assign new_n41078_ = ~new_n41075_ & ~new_n41077_;
  assign new_n41079_ = ~\b[18]  & ~new_n41078_;
  assign new_n41080_ = ~new_n40515_ & new_n40715_;
  assign new_n41081_ = ~new_n40711_ & new_n41080_;
  assign new_n41082_ = ~new_n40712_ & ~new_n40715_;
  assign new_n41083_ = ~new_n41081_ & ~new_n41082_;
  assign new_n41084_ = ~new_n40852_ & ~new_n41083_;
  assign new_n41085_ = ~new_n40505_ & ~new_n40851_;
  assign new_n41086_ = ~new_n40850_ & new_n41085_;
  assign new_n41087_ = ~new_n41084_ & ~new_n41086_;
  assign new_n41088_ = ~\b[17]  & ~new_n41087_;
  assign new_n41089_ = ~new_n40524_ & new_n40710_;
  assign new_n41090_ = ~new_n40706_ & new_n41089_;
  assign new_n41091_ = ~new_n40707_ & ~new_n40710_;
  assign new_n41092_ = ~new_n41090_ & ~new_n41091_;
  assign new_n41093_ = ~new_n40852_ & ~new_n41092_;
  assign new_n41094_ = ~new_n40514_ & ~new_n40851_;
  assign new_n41095_ = ~new_n40850_ & new_n41094_;
  assign new_n41096_ = ~new_n41093_ & ~new_n41095_;
  assign new_n41097_ = ~\b[16]  & ~new_n41096_;
  assign new_n41098_ = ~new_n40533_ & new_n40705_;
  assign new_n41099_ = ~new_n40701_ & new_n41098_;
  assign new_n41100_ = ~new_n40702_ & ~new_n40705_;
  assign new_n41101_ = ~new_n41099_ & ~new_n41100_;
  assign new_n41102_ = ~new_n40852_ & ~new_n41101_;
  assign new_n41103_ = ~new_n40523_ & ~new_n40851_;
  assign new_n41104_ = ~new_n40850_ & new_n41103_;
  assign new_n41105_ = ~new_n41102_ & ~new_n41104_;
  assign new_n41106_ = ~\b[15]  & ~new_n41105_;
  assign new_n41107_ = ~new_n40542_ & new_n40700_;
  assign new_n41108_ = ~new_n40696_ & new_n41107_;
  assign new_n41109_ = ~new_n40697_ & ~new_n40700_;
  assign new_n41110_ = ~new_n41108_ & ~new_n41109_;
  assign new_n41111_ = ~new_n40852_ & ~new_n41110_;
  assign new_n41112_ = ~new_n40532_ & ~new_n40851_;
  assign new_n41113_ = ~new_n40850_ & new_n41112_;
  assign new_n41114_ = ~new_n41111_ & ~new_n41113_;
  assign new_n41115_ = ~\b[14]  & ~new_n41114_;
  assign new_n41116_ = ~new_n40551_ & new_n40695_;
  assign new_n41117_ = ~new_n40691_ & new_n41116_;
  assign new_n41118_ = ~new_n40692_ & ~new_n40695_;
  assign new_n41119_ = ~new_n41117_ & ~new_n41118_;
  assign new_n41120_ = ~new_n40852_ & ~new_n41119_;
  assign new_n41121_ = ~new_n40541_ & ~new_n40851_;
  assign new_n41122_ = ~new_n40850_ & new_n41121_;
  assign new_n41123_ = ~new_n41120_ & ~new_n41122_;
  assign new_n41124_ = ~\b[13]  & ~new_n41123_;
  assign new_n41125_ = ~new_n40560_ & new_n40690_;
  assign new_n41126_ = ~new_n40686_ & new_n41125_;
  assign new_n41127_ = ~new_n40687_ & ~new_n40690_;
  assign new_n41128_ = ~new_n41126_ & ~new_n41127_;
  assign new_n41129_ = ~new_n40852_ & ~new_n41128_;
  assign new_n41130_ = ~new_n40550_ & ~new_n40851_;
  assign new_n41131_ = ~new_n40850_ & new_n41130_;
  assign new_n41132_ = ~new_n41129_ & ~new_n41131_;
  assign new_n41133_ = ~\b[12]  & ~new_n41132_;
  assign new_n41134_ = ~new_n40569_ & new_n40685_;
  assign new_n41135_ = ~new_n40681_ & new_n41134_;
  assign new_n41136_ = ~new_n40682_ & ~new_n40685_;
  assign new_n41137_ = ~new_n41135_ & ~new_n41136_;
  assign new_n41138_ = ~new_n40852_ & ~new_n41137_;
  assign new_n41139_ = ~new_n40559_ & ~new_n40851_;
  assign new_n41140_ = ~new_n40850_ & new_n41139_;
  assign new_n41141_ = ~new_n41138_ & ~new_n41140_;
  assign new_n41142_ = ~\b[11]  & ~new_n41141_;
  assign new_n41143_ = ~new_n40578_ & new_n40680_;
  assign new_n41144_ = ~new_n40676_ & new_n41143_;
  assign new_n41145_ = ~new_n40677_ & ~new_n40680_;
  assign new_n41146_ = ~new_n41144_ & ~new_n41145_;
  assign new_n41147_ = ~new_n40852_ & ~new_n41146_;
  assign new_n41148_ = ~new_n40568_ & ~new_n40851_;
  assign new_n41149_ = ~new_n40850_ & new_n41148_;
  assign new_n41150_ = ~new_n41147_ & ~new_n41149_;
  assign new_n41151_ = ~\b[10]  & ~new_n41150_;
  assign new_n41152_ = ~new_n40587_ & new_n40675_;
  assign new_n41153_ = ~new_n40671_ & new_n41152_;
  assign new_n41154_ = ~new_n40672_ & ~new_n40675_;
  assign new_n41155_ = ~new_n41153_ & ~new_n41154_;
  assign new_n41156_ = ~new_n40852_ & ~new_n41155_;
  assign new_n41157_ = ~new_n40577_ & ~new_n40851_;
  assign new_n41158_ = ~new_n40850_ & new_n41157_;
  assign new_n41159_ = ~new_n41156_ & ~new_n41158_;
  assign new_n41160_ = ~\b[9]  & ~new_n41159_;
  assign new_n41161_ = ~new_n40596_ & new_n40670_;
  assign new_n41162_ = ~new_n40666_ & new_n41161_;
  assign new_n41163_ = ~new_n40667_ & ~new_n40670_;
  assign new_n41164_ = ~new_n41162_ & ~new_n41163_;
  assign new_n41165_ = ~new_n40852_ & ~new_n41164_;
  assign new_n41166_ = ~new_n40586_ & ~new_n40851_;
  assign new_n41167_ = ~new_n40850_ & new_n41166_;
  assign new_n41168_ = ~new_n41165_ & ~new_n41167_;
  assign new_n41169_ = ~\b[8]  & ~new_n41168_;
  assign new_n41170_ = ~new_n40605_ & new_n40665_;
  assign new_n41171_ = ~new_n40661_ & new_n41170_;
  assign new_n41172_ = ~new_n40662_ & ~new_n40665_;
  assign new_n41173_ = ~new_n41171_ & ~new_n41172_;
  assign new_n41174_ = ~new_n40852_ & ~new_n41173_;
  assign new_n41175_ = ~new_n40595_ & ~new_n40851_;
  assign new_n41176_ = ~new_n40850_ & new_n41175_;
  assign new_n41177_ = ~new_n41174_ & ~new_n41176_;
  assign new_n41178_ = ~\b[7]  & ~new_n41177_;
  assign new_n41179_ = ~new_n40614_ & new_n40660_;
  assign new_n41180_ = ~new_n40656_ & new_n41179_;
  assign new_n41181_ = ~new_n40657_ & ~new_n40660_;
  assign new_n41182_ = ~new_n41180_ & ~new_n41181_;
  assign new_n41183_ = ~new_n40852_ & ~new_n41182_;
  assign new_n41184_ = ~new_n40604_ & ~new_n40851_;
  assign new_n41185_ = ~new_n40850_ & new_n41184_;
  assign new_n41186_ = ~new_n41183_ & ~new_n41185_;
  assign new_n41187_ = ~\b[6]  & ~new_n41186_;
  assign new_n41188_ = ~new_n40623_ & new_n40655_;
  assign new_n41189_ = ~new_n40651_ & new_n41188_;
  assign new_n41190_ = ~new_n40652_ & ~new_n40655_;
  assign new_n41191_ = ~new_n41189_ & ~new_n41190_;
  assign new_n41192_ = ~new_n40852_ & ~new_n41191_;
  assign new_n41193_ = ~new_n40613_ & ~new_n40851_;
  assign new_n41194_ = ~new_n40850_ & new_n41193_;
  assign new_n41195_ = ~new_n41192_ & ~new_n41194_;
  assign new_n41196_ = ~\b[5]  & ~new_n41195_;
  assign new_n41197_ = ~new_n40631_ & new_n40650_;
  assign new_n41198_ = ~new_n40646_ & new_n41197_;
  assign new_n41199_ = ~new_n40647_ & ~new_n40650_;
  assign new_n41200_ = ~new_n41198_ & ~new_n41199_;
  assign new_n41201_ = ~new_n40852_ & ~new_n41200_;
  assign new_n41202_ = ~new_n40622_ & ~new_n40851_;
  assign new_n41203_ = ~new_n40850_ & new_n41202_;
  assign new_n41204_ = ~new_n41201_ & ~new_n41203_;
  assign new_n41205_ = ~\b[4]  & ~new_n41204_;
  assign new_n41206_ = ~new_n40641_ & new_n40645_;
  assign new_n41207_ = ~new_n40640_ & new_n41206_;
  assign new_n41208_ = ~new_n40642_ & ~new_n40645_;
  assign new_n41209_ = ~new_n41207_ & ~new_n41208_;
  assign new_n41210_ = ~new_n40852_ & ~new_n41209_;
  assign new_n41211_ = ~new_n40630_ & ~new_n40851_;
  assign new_n41212_ = ~new_n40850_ & new_n41211_;
  assign new_n41213_ = ~new_n41210_ & ~new_n41212_;
  assign new_n41214_ = ~\b[3]  & ~new_n41213_;
  assign new_n41215_ = new_n12551_ & ~new_n40638_;
  assign new_n41216_ = ~new_n40636_ & new_n41215_;
  assign new_n41217_ = ~new_n40640_ & ~new_n41216_;
  assign new_n41218_ = ~new_n40852_ & new_n41217_;
  assign new_n41219_ = ~new_n40635_ & ~new_n40851_;
  assign new_n41220_ = ~new_n40850_ & new_n41219_;
  assign new_n41221_ = ~new_n41218_ & ~new_n41220_;
  assign new_n41222_ = ~\b[2]  & ~new_n41221_;
  assign new_n41223_ = \b[0]  & ~new_n40852_;
  assign new_n41224_ = \a[22]  & ~new_n41223_;
  assign new_n41225_ = new_n12551_ & ~new_n40852_;
  assign new_n41226_ = ~new_n41224_ & ~new_n41225_;
  assign new_n41227_ = \b[1]  & ~new_n41226_;
  assign new_n41228_ = ~\b[1]  & ~new_n41225_;
  assign new_n41229_ = ~new_n41224_ & new_n41228_;
  assign new_n41230_ = ~new_n41227_ & ~new_n41229_;
  assign new_n41231_ = ~new_n13145_ & ~new_n41230_;
  assign new_n41232_ = ~\b[1]  & ~new_n41226_;
  assign new_n41233_ = ~new_n41231_ & ~new_n41232_;
  assign new_n41234_ = \b[2]  & ~new_n41220_;
  assign new_n41235_ = ~new_n41218_ & new_n41234_;
  assign new_n41236_ = ~new_n41222_ & ~new_n41235_;
  assign new_n41237_ = ~new_n41233_ & new_n41236_;
  assign new_n41238_ = ~new_n41222_ & ~new_n41237_;
  assign new_n41239_ = \b[3]  & ~new_n41212_;
  assign new_n41240_ = ~new_n41210_ & new_n41239_;
  assign new_n41241_ = ~new_n41214_ & ~new_n41240_;
  assign new_n41242_ = ~new_n41238_ & new_n41241_;
  assign new_n41243_ = ~new_n41214_ & ~new_n41242_;
  assign new_n41244_ = \b[4]  & ~new_n41203_;
  assign new_n41245_ = ~new_n41201_ & new_n41244_;
  assign new_n41246_ = ~new_n41205_ & ~new_n41245_;
  assign new_n41247_ = ~new_n41243_ & new_n41246_;
  assign new_n41248_ = ~new_n41205_ & ~new_n41247_;
  assign new_n41249_ = \b[5]  & ~new_n41194_;
  assign new_n41250_ = ~new_n41192_ & new_n41249_;
  assign new_n41251_ = ~new_n41196_ & ~new_n41250_;
  assign new_n41252_ = ~new_n41248_ & new_n41251_;
  assign new_n41253_ = ~new_n41196_ & ~new_n41252_;
  assign new_n41254_ = \b[6]  & ~new_n41185_;
  assign new_n41255_ = ~new_n41183_ & new_n41254_;
  assign new_n41256_ = ~new_n41187_ & ~new_n41255_;
  assign new_n41257_ = ~new_n41253_ & new_n41256_;
  assign new_n41258_ = ~new_n41187_ & ~new_n41257_;
  assign new_n41259_ = \b[7]  & ~new_n41176_;
  assign new_n41260_ = ~new_n41174_ & new_n41259_;
  assign new_n41261_ = ~new_n41178_ & ~new_n41260_;
  assign new_n41262_ = ~new_n41258_ & new_n41261_;
  assign new_n41263_ = ~new_n41178_ & ~new_n41262_;
  assign new_n41264_ = \b[8]  & ~new_n41167_;
  assign new_n41265_ = ~new_n41165_ & new_n41264_;
  assign new_n41266_ = ~new_n41169_ & ~new_n41265_;
  assign new_n41267_ = ~new_n41263_ & new_n41266_;
  assign new_n41268_ = ~new_n41169_ & ~new_n41267_;
  assign new_n41269_ = \b[9]  & ~new_n41158_;
  assign new_n41270_ = ~new_n41156_ & new_n41269_;
  assign new_n41271_ = ~new_n41160_ & ~new_n41270_;
  assign new_n41272_ = ~new_n41268_ & new_n41271_;
  assign new_n41273_ = ~new_n41160_ & ~new_n41272_;
  assign new_n41274_ = \b[10]  & ~new_n41149_;
  assign new_n41275_ = ~new_n41147_ & new_n41274_;
  assign new_n41276_ = ~new_n41151_ & ~new_n41275_;
  assign new_n41277_ = ~new_n41273_ & new_n41276_;
  assign new_n41278_ = ~new_n41151_ & ~new_n41277_;
  assign new_n41279_ = \b[11]  & ~new_n41140_;
  assign new_n41280_ = ~new_n41138_ & new_n41279_;
  assign new_n41281_ = ~new_n41142_ & ~new_n41280_;
  assign new_n41282_ = ~new_n41278_ & new_n41281_;
  assign new_n41283_ = ~new_n41142_ & ~new_n41282_;
  assign new_n41284_ = \b[12]  & ~new_n41131_;
  assign new_n41285_ = ~new_n41129_ & new_n41284_;
  assign new_n41286_ = ~new_n41133_ & ~new_n41285_;
  assign new_n41287_ = ~new_n41283_ & new_n41286_;
  assign new_n41288_ = ~new_n41133_ & ~new_n41287_;
  assign new_n41289_ = \b[13]  & ~new_n41122_;
  assign new_n41290_ = ~new_n41120_ & new_n41289_;
  assign new_n41291_ = ~new_n41124_ & ~new_n41290_;
  assign new_n41292_ = ~new_n41288_ & new_n41291_;
  assign new_n41293_ = ~new_n41124_ & ~new_n41292_;
  assign new_n41294_ = \b[14]  & ~new_n41113_;
  assign new_n41295_ = ~new_n41111_ & new_n41294_;
  assign new_n41296_ = ~new_n41115_ & ~new_n41295_;
  assign new_n41297_ = ~new_n41293_ & new_n41296_;
  assign new_n41298_ = ~new_n41115_ & ~new_n41297_;
  assign new_n41299_ = \b[15]  & ~new_n41104_;
  assign new_n41300_ = ~new_n41102_ & new_n41299_;
  assign new_n41301_ = ~new_n41106_ & ~new_n41300_;
  assign new_n41302_ = ~new_n41298_ & new_n41301_;
  assign new_n41303_ = ~new_n41106_ & ~new_n41302_;
  assign new_n41304_ = \b[16]  & ~new_n41095_;
  assign new_n41305_ = ~new_n41093_ & new_n41304_;
  assign new_n41306_ = ~new_n41097_ & ~new_n41305_;
  assign new_n41307_ = ~new_n41303_ & new_n41306_;
  assign new_n41308_ = ~new_n41097_ & ~new_n41307_;
  assign new_n41309_ = \b[17]  & ~new_n41086_;
  assign new_n41310_ = ~new_n41084_ & new_n41309_;
  assign new_n41311_ = ~new_n41088_ & ~new_n41310_;
  assign new_n41312_ = ~new_n41308_ & new_n41311_;
  assign new_n41313_ = ~new_n41088_ & ~new_n41312_;
  assign new_n41314_ = \b[18]  & ~new_n41077_;
  assign new_n41315_ = ~new_n41075_ & new_n41314_;
  assign new_n41316_ = ~new_n41079_ & ~new_n41315_;
  assign new_n41317_ = ~new_n41313_ & new_n41316_;
  assign new_n41318_ = ~new_n41079_ & ~new_n41317_;
  assign new_n41319_ = \b[19]  & ~new_n41068_;
  assign new_n41320_ = ~new_n41066_ & new_n41319_;
  assign new_n41321_ = ~new_n41070_ & ~new_n41320_;
  assign new_n41322_ = ~new_n41318_ & new_n41321_;
  assign new_n41323_ = ~new_n41070_ & ~new_n41322_;
  assign new_n41324_ = \b[20]  & ~new_n41059_;
  assign new_n41325_ = ~new_n41057_ & new_n41324_;
  assign new_n41326_ = ~new_n41061_ & ~new_n41325_;
  assign new_n41327_ = ~new_n41323_ & new_n41326_;
  assign new_n41328_ = ~new_n41061_ & ~new_n41327_;
  assign new_n41329_ = \b[21]  & ~new_n41050_;
  assign new_n41330_ = ~new_n41048_ & new_n41329_;
  assign new_n41331_ = ~new_n41052_ & ~new_n41330_;
  assign new_n41332_ = ~new_n41328_ & new_n41331_;
  assign new_n41333_ = ~new_n41052_ & ~new_n41332_;
  assign new_n41334_ = \b[22]  & ~new_n41041_;
  assign new_n41335_ = ~new_n41039_ & new_n41334_;
  assign new_n41336_ = ~new_n41043_ & ~new_n41335_;
  assign new_n41337_ = ~new_n41333_ & new_n41336_;
  assign new_n41338_ = ~new_n41043_ & ~new_n41337_;
  assign new_n41339_ = \b[23]  & ~new_n41032_;
  assign new_n41340_ = ~new_n41030_ & new_n41339_;
  assign new_n41341_ = ~new_n41034_ & ~new_n41340_;
  assign new_n41342_ = ~new_n41338_ & new_n41341_;
  assign new_n41343_ = ~new_n41034_ & ~new_n41342_;
  assign new_n41344_ = \b[24]  & ~new_n41023_;
  assign new_n41345_ = ~new_n41021_ & new_n41344_;
  assign new_n41346_ = ~new_n41025_ & ~new_n41345_;
  assign new_n41347_ = ~new_n41343_ & new_n41346_;
  assign new_n41348_ = ~new_n41025_ & ~new_n41347_;
  assign new_n41349_ = \b[25]  & ~new_n41014_;
  assign new_n41350_ = ~new_n41012_ & new_n41349_;
  assign new_n41351_ = ~new_n41016_ & ~new_n41350_;
  assign new_n41352_ = ~new_n41348_ & new_n41351_;
  assign new_n41353_ = ~new_n41016_ & ~new_n41352_;
  assign new_n41354_ = \b[26]  & ~new_n41005_;
  assign new_n41355_ = ~new_n41003_ & new_n41354_;
  assign new_n41356_ = ~new_n41007_ & ~new_n41355_;
  assign new_n41357_ = ~new_n41353_ & new_n41356_;
  assign new_n41358_ = ~new_n41007_ & ~new_n41357_;
  assign new_n41359_ = \b[27]  & ~new_n40996_;
  assign new_n41360_ = ~new_n40994_ & new_n41359_;
  assign new_n41361_ = ~new_n40998_ & ~new_n41360_;
  assign new_n41362_ = ~new_n41358_ & new_n41361_;
  assign new_n41363_ = ~new_n40998_ & ~new_n41362_;
  assign new_n41364_ = \b[28]  & ~new_n40987_;
  assign new_n41365_ = ~new_n40985_ & new_n41364_;
  assign new_n41366_ = ~new_n40989_ & ~new_n41365_;
  assign new_n41367_ = ~new_n41363_ & new_n41366_;
  assign new_n41368_ = ~new_n40989_ & ~new_n41367_;
  assign new_n41369_ = \b[29]  & ~new_n40978_;
  assign new_n41370_ = ~new_n40976_ & new_n41369_;
  assign new_n41371_ = ~new_n40980_ & ~new_n41370_;
  assign new_n41372_ = ~new_n41368_ & new_n41371_;
  assign new_n41373_ = ~new_n40980_ & ~new_n41372_;
  assign new_n41374_ = \b[30]  & ~new_n40969_;
  assign new_n41375_ = ~new_n40967_ & new_n41374_;
  assign new_n41376_ = ~new_n40971_ & ~new_n41375_;
  assign new_n41377_ = ~new_n41373_ & new_n41376_;
  assign new_n41378_ = ~new_n40971_ & ~new_n41377_;
  assign new_n41379_ = \b[31]  & ~new_n40960_;
  assign new_n41380_ = ~new_n40958_ & new_n41379_;
  assign new_n41381_ = ~new_n40962_ & ~new_n41380_;
  assign new_n41382_ = ~new_n41378_ & new_n41381_;
  assign new_n41383_ = ~new_n40962_ & ~new_n41382_;
  assign new_n41384_ = \b[32]  & ~new_n40951_;
  assign new_n41385_ = ~new_n40949_ & new_n41384_;
  assign new_n41386_ = ~new_n40953_ & ~new_n41385_;
  assign new_n41387_ = ~new_n41383_ & new_n41386_;
  assign new_n41388_ = ~new_n40953_ & ~new_n41387_;
  assign new_n41389_ = \b[33]  & ~new_n40942_;
  assign new_n41390_ = ~new_n40940_ & new_n41389_;
  assign new_n41391_ = ~new_n40944_ & ~new_n41390_;
  assign new_n41392_ = ~new_n41388_ & new_n41391_;
  assign new_n41393_ = ~new_n40944_ & ~new_n41392_;
  assign new_n41394_ = \b[34]  & ~new_n40933_;
  assign new_n41395_ = ~new_n40931_ & new_n41394_;
  assign new_n41396_ = ~new_n40935_ & ~new_n41395_;
  assign new_n41397_ = ~new_n41393_ & new_n41396_;
  assign new_n41398_ = ~new_n40935_ & ~new_n41397_;
  assign new_n41399_ = \b[35]  & ~new_n40924_;
  assign new_n41400_ = ~new_n40922_ & new_n41399_;
  assign new_n41401_ = ~new_n40926_ & ~new_n41400_;
  assign new_n41402_ = ~new_n41398_ & new_n41401_;
  assign new_n41403_ = ~new_n40926_ & ~new_n41402_;
  assign new_n41404_ = \b[36]  & ~new_n40915_;
  assign new_n41405_ = ~new_n40913_ & new_n41404_;
  assign new_n41406_ = ~new_n40917_ & ~new_n41405_;
  assign new_n41407_ = ~new_n41403_ & new_n41406_;
  assign new_n41408_ = ~new_n40917_ & ~new_n41407_;
  assign new_n41409_ = \b[37]  & ~new_n40906_;
  assign new_n41410_ = ~new_n40904_ & new_n41409_;
  assign new_n41411_ = ~new_n40908_ & ~new_n41410_;
  assign new_n41412_ = ~new_n41408_ & new_n41411_;
  assign new_n41413_ = ~new_n40908_ & ~new_n41412_;
  assign new_n41414_ = \b[38]  & ~new_n40897_;
  assign new_n41415_ = ~new_n40895_ & new_n41414_;
  assign new_n41416_ = ~new_n40899_ & ~new_n41415_;
  assign new_n41417_ = ~new_n41413_ & new_n41416_;
  assign new_n41418_ = ~new_n40899_ & ~new_n41417_;
  assign new_n41419_ = \b[39]  & ~new_n40888_;
  assign new_n41420_ = ~new_n40886_ & new_n41419_;
  assign new_n41421_ = ~new_n40890_ & ~new_n41420_;
  assign new_n41422_ = ~new_n41418_ & new_n41421_;
  assign new_n41423_ = ~new_n40890_ & ~new_n41422_;
  assign new_n41424_ = \b[40]  & ~new_n40879_;
  assign new_n41425_ = ~new_n40877_ & new_n41424_;
  assign new_n41426_ = ~new_n40881_ & ~new_n41425_;
  assign new_n41427_ = ~new_n41423_ & new_n41426_;
  assign new_n41428_ = ~new_n40881_ & ~new_n41427_;
  assign new_n41429_ = \b[41]  & ~new_n40859_;
  assign new_n41430_ = ~new_n40857_ & new_n41429_;
  assign new_n41431_ = ~new_n40872_ & ~new_n41430_;
  assign new_n41432_ = ~new_n41428_ & new_n41431_;
  assign new_n41433_ = ~new_n40872_ & ~new_n41432_;
  assign new_n41434_ = \b[42]  & ~new_n40869_;
  assign new_n41435_ = ~new_n40867_ & new_n41434_;
  assign new_n41436_ = ~new_n40871_ & ~new_n41435_;
  assign new_n41437_ = ~new_n41433_ & new_n41436_;
  assign new_n41438_ = ~new_n40871_ & ~new_n41437_;
  assign new_n41439_ = new_n13355_ & ~new_n41438_;
  assign new_n41440_ = ~new_n40860_ & ~new_n41439_;
  assign new_n41441_ = ~new_n40881_ & new_n41431_;
  assign new_n41442_ = ~new_n41427_ & new_n41441_;
  assign new_n41443_ = ~new_n41428_ & ~new_n41431_;
  assign new_n41444_ = ~new_n41442_ & ~new_n41443_;
  assign new_n41445_ = new_n13355_ & ~new_n41444_;
  assign new_n41446_ = ~new_n41438_ & new_n41445_;
  assign new_n41447_ = ~new_n41440_ & ~new_n41446_;
  assign new_n41448_ = ~\b[42]  & ~new_n41447_;
  assign new_n41449_ = ~new_n40880_ & ~new_n41439_;
  assign new_n41450_ = ~new_n40890_ & new_n41426_;
  assign new_n41451_ = ~new_n41422_ & new_n41450_;
  assign new_n41452_ = ~new_n41423_ & ~new_n41426_;
  assign new_n41453_ = ~new_n41451_ & ~new_n41452_;
  assign new_n41454_ = new_n13355_ & ~new_n41453_;
  assign new_n41455_ = ~new_n41438_ & new_n41454_;
  assign new_n41456_ = ~new_n41449_ & ~new_n41455_;
  assign new_n41457_ = ~\b[41]  & ~new_n41456_;
  assign new_n41458_ = ~new_n40889_ & ~new_n41439_;
  assign new_n41459_ = ~new_n40899_ & new_n41421_;
  assign new_n41460_ = ~new_n41417_ & new_n41459_;
  assign new_n41461_ = ~new_n41418_ & ~new_n41421_;
  assign new_n41462_ = ~new_n41460_ & ~new_n41461_;
  assign new_n41463_ = new_n13355_ & ~new_n41462_;
  assign new_n41464_ = ~new_n41438_ & new_n41463_;
  assign new_n41465_ = ~new_n41458_ & ~new_n41464_;
  assign new_n41466_ = ~\b[40]  & ~new_n41465_;
  assign new_n41467_ = ~new_n40898_ & ~new_n41439_;
  assign new_n41468_ = ~new_n40908_ & new_n41416_;
  assign new_n41469_ = ~new_n41412_ & new_n41468_;
  assign new_n41470_ = ~new_n41413_ & ~new_n41416_;
  assign new_n41471_ = ~new_n41469_ & ~new_n41470_;
  assign new_n41472_ = new_n13355_ & ~new_n41471_;
  assign new_n41473_ = ~new_n41438_ & new_n41472_;
  assign new_n41474_ = ~new_n41467_ & ~new_n41473_;
  assign new_n41475_ = ~\b[39]  & ~new_n41474_;
  assign new_n41476_ = ~new_n40907_ & ~new_n41439_;
  assign new_n41477_ = ~new_n40917_ & new_n41411_;
  assign new_n41478_ = ~new_n41407_ & new_n41477_;
  assign new_n41479_ = ~new_n41408_ & ~new_n41411_;
  assign new_n41480_ = ~new_n41478_ & ~new_n41479_;
  assign new_n41481_ = new_n13355_ & ~new_n41480_;
  assign new_n41482_ = ~new_n41438_ & new_n41481_;
  assign new_n41483_ = ~new_n41476_ & ~new_n41482_;
  assign new_n41484_ = ~\b[38]  & ~new_n41483_;
  assign new_n41485_ = ~new_n40916_ & ~new_n41439_;
  assign new_n41486_ = ~new_n40926_ & new_n41406_;
  assign new_n41487_ = ~new_n41402_ & new_n41486_;
  assign new_n41488_ = ~new_n41403_ & ~new_n41406_;
  assign new_n41489_ = ~new_n41487_ & ~new_n41488_;
  assign new_n41490_ = new_n13355_ & ~new_n41489_;
  assign new_n41491_ = ~new_n41438_ & new_n41490_;
  assign new_n41492_ = ~new_n41485_ & ~new_n41491_;
  assign new_n41493_ = ~\b[37]  & ~new_n41492_;
  assign new_n41494_ = ~new_n40925_ & ~new_n41439_;
  assign new_n41495_ = ~new_n40935_ & new_n41401_;
  assign new_n41496_ = ~new_n41397_ & new_n41495_;
  assign new_n41497_ = ~new_n41398_ & ~new_n41401_;
  assign new_n41498_ = ~new_n41496_ & ~new_n41497_;
  assign new_n41499_ = new_n13355_ & ~new_n41498_;
  assign new_n41500_ = ~new_n41438_ & new_n41499_;
  assign new_n41501_ = ~new_n41494_ & ~new_n41500_;
  assign new_n41502_ = ~\b[36]  & ~new_n41501_;
  assign new_n41503_ = ~new_n40934_ & ~new_n41439_;
  assign new_n41504_ = ~new_n40944_ & new_n41396_;
  assign new_n41505_ = ~new_n41392_ & new_n41504_;
  assign new_n41506_ = ~new_n41393_ & ~new_n41396_;
  assign new_n41507_ = ~new_n41505_ & ~new_n41506_;
  assign new_n41508_ = new_n13355_ & ~new_n41507_;
  assign new_n41509_ = ~new_n41438_ & new_n41508_;
  assign new_n41510_ = ~new_n41503_ & ~new_n41509_;
  assign new_n41511_ = ~\b[35]  & ~new_n41510_;
  assign new_n41512_ = ~new_n40943_ & ~new_n41439_;
  assign new_n41513_ = ~new_n40953_ & new_n41391_;
  assign new_n41514_ = ~new_n41387_ & new_n41513_;
  assign new_n41515_ = ~new_n41388_ & ~new_n41391_;
  assign new_n41516_ = ~new_n41514_ & ~new_n41515_;
  assign new_n41517_ = new_n13355_ & ~new_n41516_;
  assign new_n41518_ = ~new_n41438_ & new_n41517_;
  assign new_n41519_ = ~new_n41512_ & ~new_n41518_;
  assign new_n41520_ = ~\b[34]  & ~new_n41519_;
  assign new_n41521_ = ~new_n40952_ & ~new_n41439_;
  assign new_n41522_ = ~new_n40962_ & new_n41386_;
  assign new_n41523_ = ~new_n41382_ & new_n41522_;
  assign new_n41524_ = ~new_n41383_ & ~new_n41386_;
  assign new_n41525_ = ~new_n41523_ & ~new_n41524_;
  assign new_n41526_ = new_n13355_ & ~new_n41525_;
  assign new_n41527_ = ~new_n41438_ & new_n41526_;
  assign new_n41528_ = ~new_n41521_ & ~new_n41527_;
  assign new_n41529_ = ~\b[33]  & ~new_n41528_;
  assign new_n41530_ = ~new_n40961_ & ~new_n41439_;
  assign new_n41531_ = ~new_n40971_ & new_n41381_;
  assign new_n41532_ = ~new_n41377_ & new_n41531_;
  assign new_n41533_ = ~new_n41378_ & ~new_n41381_;
  assign new_n41534_ = ~new_n41532_ & ~new_n41533_;
  assign new_n41535_ = new_n13355_ & ~new_n41534_;
  assign new_n41536_ = ~new_n41438_ & new_n41535_;
  assign new_n41537_ = ~new_n41530_ & ~new_n41536_;
  assign new_n41538_ = ~\b[32]  & ~new_n41537_;
  assign new_n41539_ = ~new_n40970_ & ~new_n41439_;
  assign new_n41540_ = ~new_n40980_ & new_n41376_;
  assign new_n41541_ = ~new_n41372_ & new_n41540_;
  assign new_n41542_ = ~new_n41373_ & ~new_n41376_;
  assign new_n41543_ = ~new_n41541_ & ~new_n41542_;
  assign new_n41544_ = new_n13355_ & ~new_n41543_;
  assign new_n41545_ = ~new_n41438_ & new_n41544_;
  assign new_n41546_ = ~new_n41539_ & ~new_n41545_;
  assign new_n41547_ = ~\b[31]  & ~new_n41546_;
  assign new_n41548_ = ~new_n40979_ & ~new_n41439_;
  assign new_n41549_ = ~new_n40989_ & new_n41371_;
  assign new_n41550_ = ~new_n41367_ & new_n41549_;
  assign new_n41551_ = ~new_n41368_ & ~new_n41371_;
  assign new_n41552_ = ~new_n41550_ & ~new_n41551_;
  assign new_n41553_ = new_n13355_ & ~new_n41552_;
  assign new_n41554_ = ~new_n41438_ & new_n41553_;
  assign new_n41555_ = ~new_n41548_ & ~new_n41554_;
  assign new_n41556_ = ~\b[30]  & ~new_n41555_;
  assign new_n41557_ = ~new_n40988_ & ~new_n41439_;
  assign new_n41558_ = ~new_n40998_ & new_n41366_;
  assign new_n41559_ = ~new_n41362_ & new_n41558_;
  assign new_n41560_ = ~new_n41363_ & ~new_n41366_;
  assign new_n41561_ = ~new_n41559_ & ~new_n41560_;
  assign new_n41562_ = new_n13355_ & ~new_n41561_;
  assign new_n41563_ = ~new_n41438_ & new_n41562_;
  assign new_n41564_ = ~new_n41557_ & ~new_n41563_;
  assign new_n41565_ = ~\b[29]  & ~new_n41564_;
  assign new_n41566_ = ~new_n40997_ & ~new_n41439_;
  assign new_n41567_ = ~new_n41007_ & new_n41361_;
  assign new_n41568_ = ~new_n41357_ & new_n41567_;
  assign new_n41569_ = ~new_n41358_ & ~new_n41361_;
  assign new_n41570_ = ~new_n41568_ & ~new_n41569_;
  assign new_n41571_ = new_n13355_ & ~new_n41570_;
  assign new_n41572_ = ~new_n41438_ & new_n41571_;
  assign new_n41573_ = ~new_n41566_ & ~new_n41572_;
  assign new_n41574_ = ~\b[28]  & ~new_n41573_;
  assign new_n41575_ = ~new_n41006_ & ~new_n41439_;
  assign new_n41576_ = ~new_n41016_ & new_n41356_;
  assign new_n41577_ = ~new_n41352_ & new_n41576_;
  assign new_n41578_ = ~new_n41353_ & ~new_n41356_;
  assign new_n41579_ = ~new_n41577_ & ~new_n41578_;
  assign new_n41580_ = new_n13355_ & ~new_n41579_;
  assign new_n41581_ = ~new_n41438_ & new_n41580_;
  assign new_n41582_ = ~new_n41575_ & ~new_n41581_;
  assign new_n41583_ = ~\b[27]  & ~new_n41582_;
  assign new_n41584_ = ~new_n41015_ & ~new_n41439_;
  assign new_n41585_ = ~new_n41025_ & new_n41351_;
  assign new_n41586_ = ~new_n41347_ & new_n41585_;
  assign new_n41587_ = ~new_n41348_ & ~new_n41351_;
  assign new_n41588_ = ~new_n41586_ & ~new_n41587_;
  assign new_n41589_ = new_n13355_ & ~new_n41588_;
  assign new_n41590_ = ~new_n41438_ & new_n41589_;
  assign new_n41591_ = ~new_n41584_ & ~new_n41590_;
  assign new_n41592_ = ~\b[26]  & ~new_n41591_;
  assign new_n41593_ = ~new_n41024_ & ~new_n41439_;
  assign new_n41594_ = ~new_n41034_ & new_n41346_;
  assign new_n41595_ = ~new_n41342_ & new_n41594_;
  assign new_n41596_ = ~new_n41343_ & ~new_n41346_;
  assign new_n41597_ = ~new_n41595_ & ~new_n41596_;
  assign new_n41598_ = new_n13355_ & ~new_n41597_;
  assign new_n41599_ = ~new_n41438_ & new_n41598_;
  assign new_n41600_ = ~new_n41593_ & ~new_n41599_;
  assign new_n41601_ = ~\b[25]  & ~new_n41600_;
  assign new_n41602_ = ~new_n41033_ & ~new_n41439_;
  assign new_n41603_ = ~new_n41043_ & new_n41341_;
  assign new_n41604_ = ~new_n41337_ & new_n41603_;
  assign new_n41605_ = ~new_n41338_ & ~new_n41341_;
  assign new_n41606_ = ~new_n41604_ & ~new_n41605_;
  assign new_n41607_ = new_n13355_ & ~new_n41606_;
  assign new_n41608_ = ~new_n41438_ & new_n41607_;
  assign new_n41609_ = ~new_n41602_ & ~new_n41608_;
  assign new_n41610_ = ~\b[24]  & ~new_n41609_;
  assign new_n41611_ = ~new_n41042_ & ~new_n41439_;
  assign new_n41612_ = ~new_n41052_ & new_n41336_;
  assign new_n41613_ = ~new_n41332_ & new_n41612_;
  assign new_n41614_ = ~new_n41333_ & ~new_n41336_;
  assign new_n41615_ = ~new_n41613_ & ~new_n41614_;
  assign new_n41616_ = new_n13355_ & ~new_n41615_;
  assign new_n41617_ = ~new_n41438_ & new_n41616_;
  assign new_n41618_ = ~new_n41611_ & ~new_n41617_;
  assign new_n41619_ = ~\b[23]  & ~new_n41618_;
  assign new_n41620_ = ~new_n41051_ & ~new_n41439_;
  assign new_n41621_ = ~new_n41061_ & new_n41331_;
  assign new_n41622_ = ~new_n41327_ & new_n41621_;
  assign new_n41623_ = ~new_n41328_ & ~new_n41331_;
  assign new_n41624_ = ~new_n41622_ & ~new_n41623_;
  assign new_n41625_ = new_n13355_ & ~new_n41624_;
  assign new_n41626_ = ~new_n41438_ & new_n41625_;
  assign new_n41627_ = ~new_n41620_ & ~new_n41626_;
  assign new_n41628_ = ~\b[22]  & ~new_n41627_;
  assign new_n41629_ = ~new_n41060_ & ~new_n41439_;
  assign new_n41630_ = ~new_n41070_ & new_n41326_;
  assign new_n41631_ = ~new_n41322_ & new_n41630_;
  assign new_n41632_ = ~new_n41323_ & ~new_n41326_;
  assign new_n41633_ = ~new_n41631_ & ~new_n41632_;
  assign new_n41634_ = new_n13355_ & ~new_n41633_;
  assign new_n41635_ = ~new_n41438_ & new_n41634_;
  assign new_n41636_ = ~new_n41629_ & ~new_n41635_;
  assign new_n41637_ = ~\b[21]  & ~new_n41636_;
  assign new_n41638_ = ~new_n41069_ & ~new_n41439_;
  assign new_n41639_ = ~new_n41079_ & new_n41321_;
  assign new_n41640_ = ~new_n41317_ & new_n41639_;
  assign new_n41641_ = ~new_n41318_ & ~new_n41321_;
  assign new_n41642_ = ~new_n41640_ & ~new_n41641_;
  assign new_n41643_ = new_n13355_ & ~new_n41642_;
  assign new_n41644_ = ~new_n41438_ & new_n41643_;
  assign new_n41645_ = ~new_n41638_ & ~new_n41644_;
  assign new_n41646_ = ~\b[20]  & ~new_n41645_;
  assign new_n41647_ = ~new_n41078_ & ~new_n41439_;
  assign new_n41648_ = ~new_n41088_ & new_n41316_;
  assign new_n41649_ = ~new_n41312_ & new_n41648_;
  assign new_n41650_ = ~new_n41313_ & ~new_n41316_;
  assign new_n41651_ = ~new_n41649_ & ~new_n41650_;
  assign new_n41652_ = new_n13355_ & ~new_n41651_;
  assign new_n41653_ = ~new_n41438_ & new_n41652_;
  assign new_n41654_ = ~new_n41647_ & ~new_n41653_;
  assign new_n41655_ = ~\b[19]  & ~new_n41654_;
  assign new_n41656_ = ~new_n41087_ & ~new_n41439_;
  assign new_n41657_ = ~new_n41097_ & new_n41311_;
  assign new_n41658_ = ~new_n41307_ & new_n41657_;
  assign new_n41659_ = ~new_n41308_ & ~new_n41311_;
  assign new_n41660_ = ~new_n41658_ & ~new_n41659_;
  assign new_n41661_ = new_n13355_ & ~new_n41660_;
  assign new_n41662_ = ~new_n41438_ & new_n41661_;
  assign new_n41663_ = ~new_n41656_ & ~new_n41662_;
  assign new_n41664_ = ~\b[18]  & ~new_n41663_;
  assign new_n41665_ = ~new_n41096_ & ~new_n41439_;
  assign new_n41666_ = ~new_n41106_ & new_n41306_;
  assign new_n41667_ = ~new_n41302_ & new_n41666_;
  assign new_n41668_ = ~new_n41303_ & ~new_n41306_;
  assign new_n41669_ = ~new_n41667_ & ~new_n41668_;
  assign new_n41670_ = new_n13355_ & ~new_n41669_;
  assign new_n41671_ = ~new_n41438_ & new_n41670_;
  assign new_n41672_ = ~new_n41665_ & ~new_n41671_;
  assign new_n41673_ = ~\b[17]  & ~new_n41672_;
  assign new_n41674_ = ~new_n41105_ & ~new_n41439_;
  assign new_n41675_ = ~new_n41115_ & new_n41301_;
  assign new_n41676_ = ~new_n41297_ & new_n41675_;
  assign new_n41677_ = ~new_n41298_ & ~new_n41301_;
  assign new_n41678_ = ~new_n41676_ & ~new_n41677_;
  assign new_n41679_ = new_n13355_ & ~new_n41678_;
  assign new_n41680_ = ~new_n41438_ & new_n41679_;
  assign new_n41681_ = ~new_n41674_ & ~new_n41680_;
  assign new_n41682_ = ~\b[16]  & ~new_n41681_;
  assign new_n41683_ = ~new_n41114_ & ~new_n41439_;
  assign new_n41684_ = ~new_n41124_ & new_n41296_;
  assign new_n41685_ = ~new_n41292_ & new_n41684_;
  assign new_n41686_ = ~new_n41293_ & ~new_n41296_;
  assign new_n41687_ = ~new_n41685_ & ~new_n41686_;
  assign new_n41688_ = new_n13355_ & ~new_n41687_;
  assign new_n41689_ = ~new_n41438_ & new_n41688_;
  assign new_n41690_ = ~new_n41683_ & ~new_n41689_;
  assign new_n41691_ = ~\b[15]  & ~new_n41690_;
  assign new_n41692_ = ~new_n41123_ & ~new_n41439_;
  assign new_n41693_ = ~new_n41133_ & new_n41291_;
  assign new_n41694_ = ~new_n41287_ & new_n41693_;
  assign new_n41695_ = ~new_n41288_ & ~new_n41291_;
  assign new_n41696_ = ~new_n41694_ & ~new_n41695_;
  assign new_n41697_ = new_n13355_ & ~new_n41696_;
  assign new_n41698_ = ~new_n41438_ & new_n41697_;
  assign new_n41699_ = ~new_n41692_ & ~new_n41698_;
  assign new_n41700_ = ~\b[14]  & ~new_n41699_;
  assign new_n41701_ = ~new_n41132_ & ~new_n41439_;
  assign new_n41702_ = ~new_n41142_ & new_n41286_;
  assign new_n41703_ = ~new_n41282_ & new_n41702_;
  assign new_n41704_ = ~new_n41283_ & ~new_n41286_;
  assign new_n41705_ = ~new_n41703_ & ~new_n41704_;
  assign new_n41706_ = new_n13355_ & ~new_n41705_;
  assign new_n41707_ = ~new_n41438_ & new_n41706_;
  assign new_n41708_ = ~new_n41701_ & ~new_n41707_;
  assign new_n41709_ = ~\b[13]  & ~new_n41708_;
  assign new_n41710_ = ~new_n41141_ & ~new_n41439_;
  assign new_n41711_ = ~new_n41151_ & new_n41281_;
  assign new_n41712_ = ~new_n41277_ & new_n41711_;
  assign new_n41713_ = ~new_n41278_ & ~new_n41281_;
  assign new_n41714_ = ~new_n41712_ & ~new_n41713_;
  assign new_n41715_ = new_n13355_ & ~new_n41714_;
  assign new_n41716_ = ~new_n41438_ & new_n41715_;
  assign new_n41717_ = ~new_n41710_ & ~new_n41716_;
  assign new_n41718_ = ~\b[12]  & ~new_n41717_;
  assign new_n41719_ = ~new_n41150_ & ~new_n41439_;
  assign new_n41720_ = ~new_n41160_ & new_n41276_;
  assign new_n41721_ = ~new_n41272_ & new_n41720_;
  assign new_n41722_ = ~new_n41273_ & ~new_n41276_;
  assign new_n41723_ = ~new_n41721_ & ~new_n41722_;
  assign new_n41724_ = new_n13355_ & ~new_n41723_;
  assign new_n41725_ = ~new_n41438_ & new_n41724_;
  assign new_n41726_ = ~new_n41719_ & ~new_n41725_;
  assign new_n41727_ = ~\b[11]  & ~new_n41726_;
  assign new_n41728_ = ~new_n41159_ & ~new_n41439_;
  assign new_n41729_ = ~new_n41169_ & new_n41271_;
  assign new_n41730_ = ~new_n41267_ & new_n41729_;
  assign new_n41731_ = ~new_n41268_ & ~new_n41271_;
  assign new_n41732_ = ~new_n41730_ & ~new_n41731_;
  assign new_n41733_ = new_n13355_ & ~new_n41732_;
  assign new_n41734_ = ~new_n41438_ & new_n41733_;
  assign new_n41735_ = ~new_n41728_ & ~new_n41734_;
  assign new_n41736_ = ~\b[10]  & ~new_n41735_;
  assign new_n41737_ = ~new_n41168_ & ~new_n41439_;
  assign new_n41738_ = ~new_n41178_ & new_n41266_;
  assign new_n41739_ = ~new_n41262_ & new_n41738_;
  assign new_n41740_ = ~new_n41263_ & ~new_n41266_;
  assign new_n41741_ = ~new_n41739_ & ~new_n41740_;
  assign new_n41742_ = new_n13355_ & ~new_n41741_;
  assign new_n41743_ = ~new_n41438_ & new_n41742_;
  assign new_n41744_ = ~new_n41737_ & ~new_n41743_;
  assign new_n41745_ = ~\b[9]  & ~new_n41744_;
  assign new_n41746_ = ~new_n41177_ & ~new_n41439_;
  assign new_n41747_ = ~new_n41187_ & new_n41261_;
  assign new_n41748_ = ~new_n41257_ & new_n41747_;
  assign new_n41749_ = ~new_n41258_ & ~new_n41261_;
  assign new_n41750_ = ~new_n41748_ & ~new_n41749_;
  assign new_n41751_ = new_n13355_ & ~new_n41750_;
  assign new_n41752_ = ~new_n41438_ & new_n41751_;
  assign new_n41753_ = ~new_n41746_ & ~new_n41752_;
  assign new_n41754_ = ~\b[8]  & ~new_n41753_;
  assign new_n41755_ = ~new_n41186_ & ~new_n41439_;
  assign new_n41756_ = ~new_n41196_ & new_n41256_;
  assign new_n41757_ = ~new_n41252_ & new_n41756_;
  assign new_n41758_ = ~new_n41253_ & ~new_n41256_;
  assign new_n41759_ = ~new_n41757_ & ~new_n41758_;
  assign new_n41760_ = new_n13355_ & ~new_n41759_;
  assign new_n41761_ = ~new_n41438_ & new_n41760_;
  assign new_n41762_ = ~new_n41755_ & ~new_n41761_;
  assign new_n41763_ = ~\b[7]  & ~new_n41762_;
  assign new_n41764_ = ~new_n41195_ & ~new_n41439_;
  assign new_n41765_ = ~new_n41205_ & new_n41251_;
  assign new_n41766_ = ~new_n41247_ & new_n41765_;
  assign new_n41767_ = ~new_n41248_ & ~new_n41251_;
  assign new_n41768_ = ~new_n41766_ & ~new_n41767_;
  assign new_n41769_ = new_n13355_ & ~new_n41768_;
  assign new_n41770_ = ~new_n41438_ & new_n41769_;
  assign new_n41771_ = ~new_n41764_ & ~new_n41770_;
  assign new_n41772_ = ~\b[6]  & ~new_n41771_;
  assign new_n41773_ = ~new_n41204_ & ~new_n41439_;
  assign new_n41774_ = ~new_n41214_ & new_n41246_;
  assign new_n41775_ = ~new_n41242_ & new_n41774_;
  assign new_n41776_ = ~new_n41243_ & ~new_n41246_;
  assign new_n41777_ = ~new_n41775_ & ~new_n41776_;
  assign new_n41778_ = new_n13355_ & ~new_n41777_;
  assign new_n41779_ = ~new_n41438_ & new_n41778_;
  assign new_n41780_ = ~new_n41773_ & ~new_n41779_;
  assign new_n41781_ = ~\b[5]  & ~new_n41780_;
  assign new_n41782_ = ~new_n41213_ & ~new_n41439_;
  assign new_n41783_ = ~new_n41222_ & new_n41241_;
  assign new_n41784_ = ~new_n41237_ & new_n41783_;
  assign new_n41785_ = ~new_n41238_ & ~new_n41241_;
  assign new_n41786_ = ~new_n41784_ & ~new_n41785_;
  assign new_n41787_ = new_n13355_ & ~new_n41786_;
  assign new_n41788_ = ~new_n41438_ & new_n41787_;
  assign new_n41789_ = ~new_n41782_ & ~new_n41788_;
  assign new_n41790_ = ~\b[4]  & ~new_n41789_;
  assign new_n41791_ = ~new_n41221_ & ~new_n41439_;
  assign new_n41792_ = ~new_n41232_ & new_n41236_;
  assign new_n41793_ = ~new_n41231_ & new_n41792_;
  assign new_n41794_ = ~new_n41233_ & ~new_n41236_;
  assign new_n41795_ = ~new_n41793_ & ~new_n41794_;
  assign new_n41796_ = new_n13355_ & ~new_n41795_;
  assign new_n41797_ = ~new_n41438_ & new_n41796_;
  assign new_n41798_ = ~new_n41791_ & ~new_n41797_;
  assign new_n41799_ = ~\b[3]  & ~new_n41798_;
  assign new_n41800_ = ~new_n41226_ & ~new_n41439_;
  assign new_n41801_ = new_n13145_ & ~new_n41229_;
  assign new_n41802_ = ~new_n41227_ & new_n41801_;
  assign new_n41803_ = new_n13355_ & ~new_n41802_;
  assign new_n41804_ = ~new_n41231_ & new_n41803_;
  assign new_n41805_ = ~new_n41438_ & new_n41804_;
  assign new_n41806_ = ~new_n41800_ & ~new_n41805_;
  assign new_n41807_ = ~\b[2]  & ~new_n41806_;
  assign new_n41808_ = new_n13727_ & ~new_n41438_;
  assign new_n41809_ = \a[21]  & ~new_n41808_;
  assign new_n41810_ = new_n13732_ & ~new_n41438_;
  assign new_n41811_ = ~new_n41809_ & ~new_n41810_;
  assign new_n41812_ = \b[1]  & ~new_n41811_;
  assign new_n41813_ = ~\b[1]  & ~new_n41810_;
  assign new_n41814_ = ~new_n41809_ & new_n41813_;
  assign new_n41815_ = ~new_n41812_ & ~new_n41814_;
  assign new_n41816_ = ~new_n13739_ & ~new_n41815_;
  assign new_n41817_ = ~\b[1]  & ~new_n41811_;
  assign new_n41818_ = ~new_n41816_ & ~new_n41817_;
  assign new_n41819_ = \b[2]  & ~new_n41805_;
  assign new_n41820_ = ~new_n41800_ & new_n41819_;
  assign new_n41821_ = ~new_n41807_ & ~new_n41820_;
  assign new_n41822_ = ~new_n41818_ & new_n41821_;
  assign new_n41823_ = ~new_n41807_ & ~new_n41822_;
  assign new_n41824_ = \b[3]  & ~new_n41797_;
  assign new_n41825_ = ~new_n41791_ & new_n41824_;
  assign new_n41826_ = ~new_n41799_ & ~new_n41825_;
  assign new_n41827_ = ~new_n41823_ & new_n41826_;
  assign new_n41828_ = ~new_n41799_ & ~new_n41827_;
  assign new_n41829_ = \b[4]  & ~new_n41788_;
  assign new_n41830_ = ~new_n41782_ & new_n41829_;
  assign new_n41831_ = ~new_n41790_ & ~new_n41830_;
  assign new_n41832_ = ~new_n41828_ & new_n41831_;
  assign new_n41833_ = ~new_n41790_ & ~new_n41832_;
  assign new_n41834_ = \b[5]  & ~new_n41779_;
  assign new_n41835_ = ~new_n41773_ & new_n41834_;
  assign new_n41836_ = ~new_n41781_ & ~new_n41835_;
  assign new_n41837_ = ~new_n41833_ & new_n41836_;
  assign new_n41838_ = ~new_n41781_ & ~new_n41837_;
  assign new_n41839_ = \b[6]  & ~new_n41770_;
  assign new_n41840_ = ~new_n41764_ & new_n41839_;
  assign new_n41841_ = ~new_n41772_ & ~new_n41840_;
  assign new_n41842_ = ~new_n41838_ & new_n41841_;
  assign new_n41843_ = ~new_n41772_ & ~new_n41842_;
  assign new_n41844_ = \b[7]  & ~new_n41761_;
  assign new_n41845_ = ~new_n41755_ & new_n41844_;
  assign new_n41846_ = ~new_n41763_ & ~new_n41845_;
  assign new_n41847_ = ~new_n41843_ & new_n41846_;
  assign new_n41848_ = ~new_n41763_ & ~new_n41847_;
  assign new_n41849_ = \b[8]  & ~new_n41752_;
  assign new_n41850_ = ~new_n41746_ & new_n41849_;
  assign new_n41851_ = ~new_n41754_ & ~new_n41850_;
  assign new_n41852_ = ~new_n41848_ & new_n41851_;
  assign new_n41853_ = ~new_n41754_ & ~new_n41852_;
  assign new_n41854_ = \b[9]  & ~new_n41743_;
  assign new_n41855_ = ~new_n41737_ & new_n41854_;
  assign new_n41856_ = ~new_n41745_ & ~new_n41855_;
  assign new_n41857_ = ~new_n41853_ & new_n41856_;
  assign new_n41858_ = ~new_n41745_ & ~new_n41857_;
  assign new_n41859_ = \b[10]  & ~new_n41734_;
  assign new_n41860_ = ~new_n41728_ & new_n41859_;
  assign new_n41861_ = ~new_n41736_ & ~new_n41860_;
  assign new_n41862_ = ~new_n41858_ & new_n41861_;
  assign new_n41863_ = ~new_n41736_ & ~new_n41862_;
  assign new_n41864_ = \b[11]  & ~new_n41725_;
  assign new_n41865_ = ~new_n41719_ & new_n41864_;
  assign new_n41866_ = ~new_n41727_ & ~new_n41865_;
  assign new_n41867_ = ~new_n41863_ & new_n41866_;
  assign new_n41868_ = ~new_n41727_ & ~new_n41867_;
  assign new_n41869_ = \b[12]  & ~new_n41716_;
  assign new_n41870_ = ~new_n41710_ & new_n41869_;
  assign new_n41871_ = ~new_n41718_ & ~new_n41870_;
  assign new_n41872_ = ~new_n41868_ & new_n41871_;
  assign new_n41873_ = ~new_n41718_ & ~new_n41872_;
  assign new_n41874_ = \b[13]  & ~new_n41707_;
  assign new_n41875_ = ~new_n41701_ & new_n41874_;
  assign new_n41876_ = ~new_n41709_ & ~new_n41875_;
  assign new_n41877_ = ~new_n41873_ & new_n41876_;
  assign new_n41878_ = ~new_n41709_ & ~new_n41877_;
  assign new_n41879_ = \b[14]  & ~new_n41698_;
  assign new_n41880_ = ~new_n41692_ & new_n41879_;
  assign new_n41881_ = ~new_n41700_ & ~new_n41880_;
  assign new_n41882_ = ~new_n41878_ & new_n41881_;
  assign new_n41883_ = ~new_n41700_ & ~new_n41882_;
  assign new_n41884_ = \b[15]  & ~new_n41689_;
  assign new_n41885_ = ~new_n41683_ & new_n41884_;
  assign new_n41886_ = ~new_n41691_ & ~new_n41885_;
  assign new_n41887_ = ~new_n41883_ & new_n41886_;
  assign new_n41888_ = ~new_n41691_ & ~new_n41887_;
  assign new_n41889_ = \b[16]  & ~new_n41680_;
  assign new_n41890_ = ~new_n41674_ & new_n41889_;
  assign new_n41891_ = ~new_n41682_ & ~new_n41890_;
  assign new_n41892_ = ~new_n41888_ & new_n41891_;
  assign new_n41893_ = ~new_n41682_ & ~new_n41892_;
  assign new_n41894_ = \b[17]  & ~new_n41671_;
  assign new_n41895_ = ~new_n41665_ & new_n41894_;
  assign new_n41896_ = ~new_n41673_ & ~new_n41895_;
  assign new_n41897_ = ~new_n41893_ & new_n41896_;
  assign new_n41898_ = ~new_n41673_ & ~new_n41897_;
  assign new_n41899_ = \b[18]  & ~new_n41662_;
  assign new_n41900_ = ~new_n41656_ & new_n41899_;
  assign new_n41901_ = ~new_n41664_ & ~new_n41900_;
  assign new_n41902_ = ~new_n41898_ & new_n41901_;
  assign new_n41903_ = ~new_n41664_ & ~new_n41902_;
  assign new_n41904_ = \b[19]  & ~new_n41653_;
  assign new_n41905_ = ~new_n41647_ & new_n41904_;
  assign new_n41906_ = ~new_n41655_ & ~new_n41905_;
  assign new_n41907_ = ~new_n41903_ & new_n41906_;
  assign new_n41908_ = ~new_n41655_ & ~new_n41907_;
  assign new_n41909_ = \b[20]  & ~new_n41644_;
  assign new_n41910_ = ~new_n41638_ & new_n41909_;
  assign new_n41911_ = ~new_n41646_ & ~new_n41910_;
  assign new_n41912_ = ~new_n41908_ & new_n41911_;
  assign new_n41913_ = ~new_n41646_ & ~new_n41912_;
  assign new_n41914_ = \b[21]  & ~new_n41635_;
  assign new_n41915_ = ~new_n41629_ & new_n41914_;
  assign new_n41916_ = ~new_n41637_ & ~new_n41915_;
  assign new_n41917_ = ~new_n41913_ & new_n41916_;
  assign new_n41918_ = ~new_n41637_ & ~new_n41917_;
  assign new_n41919_ = \b[22]  & ~new_n41626_;
  assign new_n41920_ = ~new_n41620_ & new_n41919_;
  assign new_n41921_ = ~new_n41628_ & ~new_n41920_;
  assign new_n41922_ = ~new_n41918_ & new_n41921_;
  assign new_n41923_ = ~new_n41628_ & ~new_n41922_;
  assign new_n41924_ = \b[23]  & ~new_n41617_;
  assign new_n41925_ = ~new_n41611_ & new_n41924_;
  assign new_n41926_ = ~new_n41619_ & ~new_n41925_;
  assign new_n41927_ = ~new_n41923_ & new_n41926_;
  assign new_n41928_ = ~new_n41619_ & ~new_n41927_;
  assign new_n41929_ = \b[24]  & ~new_n41608_;
  assign new_n41930_ = ~new_n41602_ & new_n41929_;
  assign new_n41931_ = ~new_n41610_ & ~new_n41930_;
  assign new_n41932_ = ~new_n41928_ & new_n41931_;
  assign new_n41933_ = ~new_n41610_ & ~new_n41932_;
  assign new_n41934_ = \b[25]  & ~new_n41599_;
  assign new_n41935_ = ~new_n41593_ & new_n41934_;
  assign new_n41936_ = ~new_n41601_ & ~new_n41935_;
  assign new_n41937_ = ~new_n41933_ & new_n41936_;
  assign new_n41938_ = ~new_n41601_ & ~new_n41937_;
  assign new_n41939_ = \b[26]  & ~new_n41590_;
  assign new_n41940_ = ~new_n41584_ & new_n41939_;
  assign new_n41941_ = ~new_n41592_ & ~new_n41940_;
  assign new_n41942_ = ~new_n41938_ & new_n41941_;
  assign new_n41943_ = ~new_n41592_ & ~new_n41942_;
  assign new_n41944_ = \b[27]  & ~new_n41581_;
  assign new_n41945_ = ~new_n41575_ & new_n41944_;
  assign new_n41946_ = ~new_n41583_ & ~new_n41945_;
  assign new_n41947_ = ~new_n41943_ & new_n41946_;
  assign new_n41948_ = ~new_n41583_ & ~new_n41947_;
  assign new_n41949_ = \b[28]  & ~new_n41572_;
  assign new_n41950_ = ~new_n41566_ & new_n41949_;
  assign new_n41951_ = ~new_n41574_ & ~new_n41950_;
  assign new_n41952_ = ~new_n41948_ & new_n41951_;
  assign new_n41953_ = ~new_n41574_ & ~new_n41952_;
  assign new_n41954_ = \b[29]  & ~new_n41563_;
  assign new_n41955_ = ~new_n41557_ & new_n41954_;
  assign new_n41956_ = ~new_n41565_ & ~new_n41955_;
  assign new_n41957_ = ~new_n41953_ & new_n41956_;
  assign new_n41958_ = ~new_n41565_ & ~new_n41957_;
  assign new_n41959_ = \b[30]  & ~new_n41554_;
  assign new_n41960_ = ~new_n41548_ & new_n41959_;
  assign new_n41961_ = ~new_n41556_ & ~new_n41960_;
  assign new_n41962_ = ~new_n41958_ & new_n41961_;
  assign new_n41963_ = ~new_n41556_ & ~new_n41962_;
  assign new_n41964_ = \b[31]  & ~new_n41545_;
  assign new_n41965_ = ~new_n41539_ & new_n41964_;
  assign new_n41966_ = ~new_n41547_ & ~new_n41965_;
  assign new_n41967_ = ~new_n41963_ & new_n41966_;
  assign new_n41968_ = ~new_n41547_ & ~new_n41967_;
  assign new_n41969_ = \b[32]  & ~new_n41536_;
  assign new_n41970_ = ~new_n41530_ & new_n41969_;
  assign new_n41971_ = ~new_n41538_ & ~new_n41970_;
  assign new_n41972_ = ~new_n41968_ & new_n41971_;
  assign new_n41973_ = ~new_n41538_ & ~new_n41972_;
  assign new_n41974_ = \b[33]  & ~new_n41527_;
  assign new_n41975_ = ~new_n41521_ & new_n41974_;
  assign new_n41976_ = ~new_n41529_ & ~new_n41975_;
  assign new_n41977_ = ~new_n41973_ & new_n41976_;
  assign new_n41978_ = ~new_n41529_ & ~new_n41977_;
  assign new_n41979_ = \b[34]  & ~new_n41518_;
  assign new_n41980_ = ~new_n41512_ & new_n41979_;
  assign new_n41981_ = ~new_n41520_ & ~new_n41980_;
  assign new_n41982_ = ~new_n41978_ & new_n41981_;
  assign new_n41983_ = ~new_n41520_ & ~new_n41982_;
  assign new_n41984_ = \b[35]  & ~new_n41509_;
  assign new_n41985_ = ~new_n41503_ & new_n41984_;
  assign new_n41986_ = ~new_n41511_ & ~new_n41985_;
  assign new_n41987_ = ~new_n41983_ & new_n41986_;
  assign new_n41988_ = ~new_n41511_ & ~new_n41987_;
  assign new_n41989_ = \b[36]  & ~new_n41500_;
  assign new_n41990_ = ~new_n41494_ & new_n41989_;
  assign new_n41991_ = ~new_n41502_ & ~new_n41990_;
  assign new_n41992_ = ~new_n41988_ & new_n41991_;
  assign new_n41993_ = ~new_n41502_ & ~new_n41992_;
  assign new_n41994_ = \b[37]  & ~new_n41491_;
  assign new_n41995_ = ~new_n41485_ & new_n41994_;
  assign new_n41996_ = ~new_n41493_ & ~new_n41995_;
  assign new_n41997_ = ~new_n41993_ & new_n41996_;
  assign new_n41998_ = ~new_n41493_ & ~new_n41997_;
  assign new_n41999_ = \b[38]  & ~new_n41482_;
  assign new_n42000_ = ~new_n41476_ & new_n41999_;
  assign new_n42001_ = ~new_n41484_ & ~new_n42000_;
  assign new_n42002_ = ~new_n41998_ & new_n42001_;
  assign new_n42003_ = ~new_n41484_ & ~new_n42002_;
  assign new_n42004_ = \b[39]  & ~new_n41473_;
  assign new_n42005_ = ~new_n41467_ & new_n42004_;
  assign new_n42006_ = ~new_n41475_ & ~new_n42005_;
  assign new_n42007_ = ~new_n42003_ & new_n42006_;
  assign new_n42008_ = ~new_n41475_ & ~new_n42007_;
  assign new_n42009_ = \b[40]  & ~new_n41464_;
  assign new_n42010_ = ~new_n41458_ & new_n42009_;
  assign new_n42011_ = ~new_n41466_ & ~new_n42010_;
  assign new_n42012_ = ~new_n42008_ & new_n42011_;
  assign new_n42013_ = ~new_n41466_ & ~new_n42012_;
  assign new_n42014_ = \b[41]  & ~new_n41455_;
  assign new_n42015_ = ~new_n41449_ & new_n42014_;
  assign new_n42016_ = ~new_n41457_ & ~new_n42015_;
  assign new_n42017_ = ~new_n42013_ & new_n42016_;
  assign new_n42018_ = ~new_n41457_ & ~new_n42017_;
  assign new_n42019_ = \b[42]  & ~new_n41446_;
  assign new_n42020_ = ~new_n41440_ & new_n42019_;
  assign new_n42021_ = ~new_n41448_ & ~new_n42020_;
  assign new_n42022_ = ~new_n42018_ & new_n42021_;
  assign new_n42023_ = ~new_n41448_ & ~new_n42022_;
  assign new_n42024_ = ~new_n40870_ & ~new_n41439_;
  assign new_n42025_ = ~new_n40872_ & new_n41436_;
  assign new_n42026_ = ~new_n41432_ & new_n42025_;
  assign new_n42027_ = ~new_n41433_ & ~new_n41436_;
  assign new_n42028_ = ~new_n42026_ & ~new_n42027_;
  assign new_n42029_ = new_n41439_ & ~new_n42028_;
  assign new_n42030_ = ~new_n42024_ & ~new_n42029_;
  assign new_n42031_ = ~\b[43]  & ~new_n42030_;
  assign new_n42032_ = \b[43]  & ~new_n42024_;
  assign new_n42033_ = ~new_n42029_ & new_n42032_;
  assign new_n42034_ = new_n13958_ & ~new_n42033_;
  assign new_n42035_ = ~new_n42031_ & new_n42034_;
  assign new_n42036_ = ~new_n42023_ & new_n42035_;
  assign new_n42037_ = new_n13355_ & ~new_n42030_;
  assign new_n42038_ = ~new_n42036_ & ~new_n42037_;
  assign new_n42039_ = ~new_n41457_ & new_n42021_;
  assign new_n42040_ = ~new_n42017_ & new_n42039_;
  assign new_n42041_ = ~new_n42018_ & ~new_n42021_;
  assign new_n42042_ = ~new_n42040_ & ~new_n42041_;
  assign new_n42043_ = ~new_n42038_ & ~new_n42042_;
  assign new_n42044_ = ~new_n41447_ & ~new_n42037_;
  assign new_n42045_ = ~new_n42036_ & new_n42044_;
  assign new_n42046_ = ~new_n42043_ & ~new_n42045_;
  assign new_n42047_ = ~\b[43]  & ~new_n42046_;
  assign new_n42048_ = ~new_n41466_ & new_n42016_;
  assign new_n42049_ = ~new_n42012_ & new_n42048_;
  assign new_n42050_ = ~new_n42013_ & ~new_n42016_;
  assign new_n42051_ = ~new_n42049_ & ~new_n42050_;
  assign new_n42052_ = ~new_n42038_ & ~new_n42051_;
  assign new_n42053_ = ~new_n41456_ & ~new_n42037_;
  assign new_n42054_ = ~new_n42036_ & new_n42053_;
  assign new_n42055_ = ~new_n42052_ & ~new_n42054_;
  assign new_n42056_ = ~\b[42]  & ~new_n42055_;
  assign new_n42057_ = ~new_n41475_ & new_n42011_;
  assign new_n42058_ = ~new_n42007_ & new_n42057_;
  assign new_n42059_ = ~new_n42008_ & ~new_n42011_;
  assign new_n42060_ = ~new_n42058_ & ~new_n42059_;
  assign new_n42061_ = ~new_n42038_ & ~new_n42060_;
  assign new_n42062_ = ~new_n41465_ & ~new_n42037_;
  assign new_n42063_ = ~new_n42036_ & new_n42062_;
  assign new_n42064_ = ~new_n42061_ & ~new_n42063_;
  assign new_n42065_ = ~\b[41]  & ~new_n42064_;
  assign new_n42066_ = ~new_n41484_ & new_n42006_;
  assign new_n42067_ = ~new_n42002_ & new_n42066_;
  assign new_n42068_ = ~new_n42003_ & ~new_n42006_;
  assign new_n42069_ = ~new_n42067_ & ~new_n42068_;
  assign new_n42070_ = ~new_n42038_ & ~new_n42069_;
  assign new_n42071_ = ~new_n41474_ & ~new_n42037_;
  assign new_n42072_ = ~new_n42036_ & new_n42071_;
  assign new_n42073_ = ~new_n42070_ & ~new_n42072_;
  assign new_n42074_ = ~\b[40]  & ~new_n42073_;
  assign new_n42075_ = ~new_n41493_ & new_n42001_;
  assign new_n42076_ = ~new_n41997_ & new_n42075_;
  assign new_n42077_ = ~new_n41998_ & ~new_n42001_;
  assign new_n42078_ = ~new_n42076_ & ~new_n42077_;
  assign new_n42079_ = ~new_n42038_ & ~new_n42078_;
  assign new_n42080_ = ~new_n41483_ & ~new_n42037_;
  assign new_n42081_ = ~new_n42036_ & new_n42080_;
  assign new_n42082_ = ~new_n42079_ & ~new_n42081_;
  assign new_n42083_ = ~\b[39]  & ~new_n42082_;
  assign new_n42084_ = ~new_n41502_ & new_n41996_;
  assign new_n42085_ = ~new_n41992_ & new_n42084_;
  assign new_n42086_ = ~new_n41993_ & ~new_n41996_;
  assign new_n42087_ = ~new_n42085_ & ~new_n42086_;
  assign new_n42088_ = ~new_n42038_ & ~new_n42087_;
  assign new_n42089_ = ~new_n41492_ & ~new_n42037_;
  assign new_n42090_ = ~new_n42036_ & new_n42089_;
  assign new_n42091_ = ~new_n42088_ & ~new_n42090_;
  assign new_n42092_ = ~\b[38]  & ~new_n42091_;
  assign new_n42093_ = ~new_n41511_ & new_n41991_;
  assign new_n42094_ = ~new_n41987_ & new_n42093_;
  assign new_n42095_ = ~new_n41988_ & ~new_n41991_;
  assign new_n42096_ = ~new_n42094_ & ~new_n42095_;
  assign new_n42097_ = ~new_n42038_ & ~new_n42096_;
  assign new_n42098_ = ~new_n41501_ & ~new_n42037_;
  assign new_n42099_ = ~new_n42036_ & new_n42098_;
  assign new_n42100_ = ~new_n42097_ & ~new_n42099_;
  assign new_n42101_ = ~\b[37]  & ~new_n42100_;
  assign new_n42102_ = ~new_n41520_ & new_n41986_;
  assign new_n42103_ = ~new_n41982_ & new_n42102_;
  assign new_n42104_ = ~new_n41983_ & ~new_n41986_;
  assign new_n42105_ = ~new_n42103_ & ~new_n42104_;
  assign new_n42106_ = ~new_n42038_ & ~new_n42105_;
  assign new_n42107_ = ~new_n41510_ & ~new_n42037_;
  assign new_n42108_ = ~new_n42036_ & new_n42107_;
  assign new_n42109_ = ~new_n42106_ & ~new_n42108_;
  assign new_n42110_ = ~\b[36]  & ~new_n42109_;
  assign new_n42111_ = ~new_n41529_ & new_n41981_;
  assign new_n42112_ = ~new_n41977_ & new_n42111_;
  assign new_n42113_ = ~new_n41978_ & ~new_n41981_;
  assign new_n42114_ = ~new_n42112_ & ~new_n42113_;
  assign new_n42115_ = ~new_n42038_ & ~new_n42114_;
  assign new_n42116_ = ~new_n41519_ & ~new_n42037_;
  assign new_n42117_ = ~new_n42036_ & new_n42116_;
  assign new_n42118_ = ~new_n42115_ & ~new_n42117_;
  assign new_n42119_ = ~\b[35]  & ~new_n42118_;
  assign new_n42120_ = ~new_n41538_ & new_n41976_;
  assign new_n42121_ = ~new_n41972_ & new_n42120_;
  assign new_n42122_ = ~new_n41973_ & ~new_n41976_;
  assign new_n42123_ = ~new_n42121_ & ~new_n42122_;
  assign new_n42124_ = ~new_n42038_ & ~new_n42123_;
  assign new_n42125_ = ~new_n41528_ & ~new_n42037_;
  assign new_n42126_ = ~new_n42036_ & new_n42125_;
  assign new_n42127_ = ~new_n42124_ & ~new_n42126_;
  assign new_n42128_ = ~\b[34]  & ~new_n42127_;
  assign new_n42129_ = ~new_n41547_ & new_n41971_;
  assign new_n42130_ = ~new_n41967_ & new_n42129_;
  assign new_n42131_ = ~new_n41968_ & ~new_n41971_;
  assign new_n42132_ = ~new_n42130_ & ~new_n42131_;
  assign new_n42133_ = ~new_n42038_ & ~new_n42132_;
  assign new_n42134_ = ~new_n41537_ & ~new_n42037_;
  assign new_n42135_ = ~new_n42036_ & new_n42134_;
  assign new_n42136_ = ~new_n42133_ & ~new_n42135_;
  assign new_n42137_ = ~\b[33]  & ~new_n42136_;
  assign new_n42138_ = ~new_n41556_ & new_n41966_;
  assign new_n42139_ = ~new_n41962_ & new_n42138_;
  assign new_n42140_ = ~new_n41963_ & ~new_n41966_;
  assign new_n42141_ = ~new_n42139_ & ~new_n42140_;
  assign new_n42142_ = ~new_n42038_ & ~new_n42141_;
  assign new_n42143_ = ~new_n41546_ & ~new_n42037_;
  assign new_n42144_ = ~new_n42036_ & new_n42143_;
  assign new_n42145_ = ~new_n42142_ & ~new_n42144_;
  assign new_n42146_ = ~\b[32]  & ~new_n42145_;
  assign new_n42147_ = ~new_n41565_ & new_n41961_;
  assign new_n42148_ = ~new_n41957_ & new_n42147_;
  assign new_n42149_ = ~new_n41958_ & ~new_n41961_;
  assign new_n42150_ = ~new_n42148_ & ~new_n42149_;
  assign new_n42151_ = ~new_n42038_ & ~new_n42150_;
  assign new_n42152_ = ~new_n41555_ & ~new_n42037_;
  assign new_n42153_ = ~new_n42036_ & new_n42152_;
  assign new_n42154_ = ~new_n42151_ & ~new_n42153_;
  assign new_n42155_ = ~\b[31]  & ~new_n42154_;
  assign new_n42156_ = ~new_n41574_ & new_n41956_;
  assign new_n42157_ = ~new_n41952_ & new_n42156_;
  assign new_n42158_ = ~new_n41953_ & ~new_n41956_;
  assign new_n42159_ = ~new_n42157_ & ~new_n42158_;
  assign new_n42160_ = ~new_n42038_ & ~new_n42159_;
  assign new_n42161_ = ~new_n41564_ & ~new_n42037_;
  assign new_n42162_ = ~new_n42036_ & new_n42161_;
  assign new_n42163_ = ~new_n42160_ & ~new_n42162_;
  assign new_n42164_ = ~\b[30]  & ~new_n42163_;
  assign new_n42165_ = ~new_n41583_ & new_n41951_;
  assign new_n42166_ = ~new_n41947_ & new_n42165_;
  assign new_n42167_ = ~new_n41948_ & ~new_n41951_;
  assign new_n42168_ = ~new_n42166_ & ~new_n42167_;
  assign new_n42169_ = ~new_n42038_ & ~new_n42168_;
  assign new_n42170_ = ~new_n41573_ & ~new_n42037_;
  assign new_n42171_ = ~new_n42036_ & new_n42170_;
  assign new_n42172_ = ~new_n42169_ & ~new_n42171_;
  assign new_n42173_ = ~\b[29]  & ~new_n42172_;
  assign new_n42174_ = ~new_n41592_ & new_n41946_;
  assign new_n42175_ = ~new_n41942_ & new_n42174_;
  assign new_n42176_ = ~new_n41943_ & ~new_n41946_;
  assign new_n42177_ = ~new_n42175_ & ~new_n42176_;
  assign new_n42178_ = ~new_n42038_ & ~new_n42177_;
  assign new_n42179_ = ~new_n41582_ & ~new_n42037_;
  assign new_n42180_ = ~new_n42036_ & new_n42179_;
  assign new_n42181_ = ~new_n42178_ & ~new_n42180_;
  assign new_n42182_ = ~\b[28]  & ~new_n42181_;
  assign new_n42183_ = ~new_n41601_ & new_n41941_;
  assign new_n42184_ = ~new_n41937_ & new_n42183_;
  assign new_n42185_ = ~new_n41938_ & ~new_n41941_;
  assign new_n42186_ = ~new_n42184_ & ~new_n42185_;
  assign new_n42187_ = ~new_n42038_ & ~new_n42186_;
  assign new_n42188_ = ~new_n41591_ & ~new_n42037_;
  assign new_n42189_ = ~new_n42036_ & new_n42188_;
  assign new_n42190_ = ~new_n42187_ & ~new_n42189_;
  assign new_n42191_ = ~\b[27]  & ~new_n42190_;
  assign new_n42192_ = ~new_n41610_ & new_n41936_;
  assign new_n42193_ = ~new_n41932_ & new_n42192_;
  assign new_n42194_ = ~new_n41933_ & ~new_n41936_;
  assign new_n42195_ = ~new_n42193_ & ~new_n42194_;
  assign new_n42196_ = ~new_n42038_ & ~new_n42195_;
  assign new_n42197_ = ~new_n41600_ & ~new_n42037_;
  assign new_n42198_ = ~new_n42036_ & new_n42197_;
  assign new_n42199_ = ~new_n42196_ & ~new_n42198_;
  assign new_n42200_ = ~\b[26]  & ~new_n42199_;
  assign new_n42201_ = ~new_n41619_ & new_n41931_;
  assign new_n42202_ = ~new_n41927_ & new_n42201_;
  assign new_n42203_ = ~new_n41928_ & ~new_n41931_;
  assign new_n42204_ = ~new_n42202_ & ~new_n42203_;
  assign new_n42205_ = ~new_n42038_ & ~new_n42204_;
  assign new_n42206_ = ~new_n41609_ & ~new_n42037_;
  assign new_n42207_ = ~new_n42036_ & new_n42206_;
  assign new_n42208_ = ~new_n42205_ & ~new_n42207_;
  assign new_n42209_ = ~\b[25]  & ~new_n42208_;
  assign new_n42210_ = ~new_n41628_ & new_n41926_;
  assign new_n42211_ = ~new_n41922_ & new_n42210_;
  assign new_n42212_ = ~new_n41923_ & ~new_n41926_;
  assign new_n42213_ = ~new_n42211_ & ~new_n42212_;
  assign new_n42214_ = ~new_n42038_ & ~new_n42213_;
  assign new_n42215_ = ~new_n41618_ & ~new_n42037_;
  assign new_n42216_ = ~new_n42036_ & new_n42215_;
  assign new_n42217_ = ~new_n42214_ & ~new_n42216_;
  assign new_n42218_ = ~\b[24]  & ~new_n42217_;
  assign new_n42219_ = ~new_n41637_ & new_n41921_;
  assign new_n42220_ = ~new_n41917_ & new_n42219_;
  assign new_n42221_ = ~new_n41918_ & ~new_n41921_;
  assign new_n42222_ = ~new_n42220_ & ~new_n42221_;
  assign new_n42223_ = ~new_n42038_ & ~new_n42222_;
  assign new_n42224_ = ~new_n41627_ & ~new_n42037_;
  assign new_n42225_ = ~new_n42036_ & new_n42224_;
  assign new_n42226_ = ~new_n42223_ & ~new_n42225_;
  assign new_n42227_ = ~\b[23]  & ~new_n42226_;
  assign new_n42228_ = ~new_n41646_ & new_n41916_;
  assign new_n42229_ = ~new_n41912_ & new_n42228_;
  assign new_n42230_ = ~new_n41913_ & ~new_n41916_;
  assign new_n42231_ = ~new_n42229_ & ~new_n42230_;
  assign new_n42232_ = ~new_n42038_ & ~new_n42231_;
  assign new_n42233_ = ~new_n41636_ & ~new_n42037_;
  assign new_n42234_ = ~new_n42036_ & new_n42233_;
  assign new_n42235_ = ~new_n42232_ & ~new_n42234_;
  assign new_n42236_ = ~\b[22]  & ~new_n42235_;
  assign new_n42237_ = ~new_n41655_ & new_n41911_;
  assign new_n42238_ = ~new_n41907_ & new_n42237_;
  assign new_n42239_ = ~new_n41908_ & ~new_n41911_;
  assign new_n42240_ = ~new_n42238_ & ~new_n42239_;
  assign new_n42241_ = ~new_n42038_ & ~new_n42240_;
  assign new_n42242_ = ~new_n41645_ & ~new_n42037_;
  assign new_n42243_ = ~new_n42036_ & new_n42242_;
  assign new_n42244_ = ~new_n42241_ & ~new_n42243_;
  assign new_n42245_ = ~\b[21]  & ~new_n42244_;
  assign new_n42246_ = ~new_n41664_ & new_n41906_;
  assign new_n42247_ = ~new_n41902_ & new_n42246_;
  assign new_n42248_ = ~new_n41903_ & ~new_n41906_;
  assign new_n42249_ = ~new_n42247_ & ~new_n42248_;
  assign new_n42250_ = ~new_n42038_ & ~new_n42249_;
  assign new_n42251_ = ~new_n41654_ & ~new_n42037_;
  assign new_n42252_ = ~new_n42036_ & new_n42251_;
  assign new_n42253_ = ~new_n42250_ & ~new_n42252_;
  assign new_n42254_ = ~\b[20]  & ~new_n42253_;
  assign new_n42255_ = ~new_n41673_ & new_n41901_;
  assign new_n42256_ = ~new_n41897_ & new_n42255_;
  assign new_n42257_ = ~new_n41898_ & ~new_n41901_;
  assign new_n42258_ = ~new_n42256_ & ~new_n42257_;
  assign new_n42259_ = ~new_n42038_ & ~new_n42258_;
  assign new_n42260_ = ~new_n41663_ & ~new_n42037_;
  assign new_n42261_ = ~new_n42036_ & new_n42260_;
  assign new_n42262_ = ~new_n42259_ & ~new_n42261_;
  assign new_n42263_ = ~\b[19]  & ~new_n42262_;
  assign new_n42264_ = ~new_n41682_ & new_n41896_;
  assign new_n42265_ = ~new_n41892_ & new_n42264_;
  assign new_n42266_ = ~new_n41893_ & ~new_n41896_;
  assign new_n42267_ = ~new_n42265_ & ~new_n42266_;
  assign new_n42268_ = ~new_n42038_ & ~new_n42267_;
  assign new_n42269_ = ~new_n41672_ & ~new_n42037_;
  assign new_n42270_ = ~new_n42036_ & new_n42269_;
  assign new_n42271_ = ~new_n42268_ & ~new_n42270_;
  assign new_n42272_ = ~\b[18]  & ~new_n42271_;
  assign new_n42273_ = ~new_n41691_ & new_n41891_;
  assign new_n42274_ = ~new_n41887_ & new_n42273_;
  assign new_n42275_ = ~new_n41888_ & ~new_n41891_;
  assign new_n42276_ = ~new_n42274_ & ~new_n42275_;
  assign new_n42277_ = ~new_n42038_ & ~new_n42276_;
  assign new_n42278_ = ~new_n41681_ & ~new_n42037_;
  assign new_n42279_ = ~new_n42036_ & new_n42278_;
  assign new_n42280_ = ~new_n42277_ & ~new_n42279_;
  assign new_n42281_ = ~\b[17]  & ~new_n42280_;
  assign new_n42282_ = ~new_n41700_ & new_n41886_;
  assign new_n42283_ = ~new_n41882_ & new_n42282_;
  assign new_n42284_ = ~new_n41883_ & ~new_n41886_;
  assign new_n42285_ = ~new_n42283_ & ~new_n42284_;
  assign new_n42286_ = ~new_n42038_ & ~new_n42285_;
  assign new_n42287_ = ~new_n41690_ & ~new_n42037_;
  assign new_n42288_ = ~new_n42036_ & new_n42287_;
  assign new_n42289_ = ~new_n42286_ & ~new_n42288_;
  assign new_n42290_ = ~\b[16]  & ~new_n42289_;
  assign new_n42291_ = ~new_n41709_ & new_n41881_;
  assign new_n42292_ = ~new_n41877_ & new_n42291_;
  assign new_n42293_ = ~new_n41878_ & ~new_n41881_;
  assign new_n42294_ = ~new_n42292_ & ~new_n42293_;
  assign new_n42295_ = ~new_n42038_ & ~new_n42294_;
  assign new_n42296_ = ~new_n41699_ & ~new_n42037_;
  assign new_n42297_ = ~new_n42036_ & new_n42296_;
  assign new_n42298_ = ~new_n42295_ & ~new_n42297_;
  assign new_n42299_ = ~\b[15]  & ~new_n42298_;
  assign new_n42300_ = ~new_n41718_ & new_n41876_;
  assign new_n42301_ = ~new_n41872_ & new_n42300_;
  assign new_n42302_ = ~new_n41873_ & ~new_n41876_;
  assign new_n42303_ = ~new_n42301_ & ~new_n42302_;
  assign new_n42304_ = ~new_n42038_ & ~new_n42303_;
  assign new_n42305_ = ~new_n41708_ & ~new_n42037_;
  assign new_n42306_ = ~new_n42036_ & new_n42305_;
  assign new_n42307_ = ~new_n42304_ & ~new_n42306_;
  assign new_n42308_ = ~\b[14]  & ~new_n42307_;
  assign new_n42309_ = ~new_n41727_ & new_n41871_;
  assign new_n42310_ = ~new_n41867_ & new_n42309_;
  assign new_n42311_ = ~new_n41868_ & ~new_n41871_;
  assign new_n42312_ = ~new_n42310_ & ~new_n42311_;
  assign new_n42313_ = ~new_n42038_ & ~new_n42312_;
  assign new_n42314_ = ~new_n41717_ & ~new_n42037_;
  assign new_n42315_ = ~new_n42036_ & new_n42314_;
  assign new_n42316_ = ~new_n42313_ & ~new_n42315_;
  assign new_n42317_ = ~\b[13]  & ~new_n42316_;
  assign new_n42318_ = ~new_n41736_ & new_n41866_;
  assign new_n42319_ = ~new_n41862_ & new_n42318_;
  assign new_n42320_ = ~new_n41863_ & ~new_n41866_;
  assign new_n42321_ = ~new_n42319_ & ~new_n42320_;
  assign new_n42322_ = ~new_n42038_ & ~new_n42321_;
  assign new_n42323_ = ~new_n41726_ & ~new_n42037_;
  assign new_n42324_ = ~new_n42036_ & new_n42323_;
  assign new_n42325_ = ~new_n42322_ & ~new_n42324_;
  assign new_n42326_ = ~\b[12]  & ~new_n42325_;
  assign new_n42327_ = ~new_n41745_ & new_n41861_;
  assign new_n42328_ = ~new_n41857_ & new_n42327_;
  assign new_n42329_ = ~new_n41858_ & ~new_n41861_;
  assign new_n42330_ = ~new_n42328_ & ~new_n42329_;
  assign new_n42331_ = ~new_n42038_ & ~new_n42330_;
  assign new_n42332_ = ~new_n41735_ & ~new_n42037_;
  assign new_n42333_ = ~new_n42036_ & new_n42332_;
  assign new_n42334_ = ~new_n42331_ & ~new_n42333_;
  assign new_n42335_ = ~\b[11]  & ~new_n42334_;
  assign new_n42336_ = ~new_n41754_ & new_n41856_;
  assign new_n42337_ = ~new_n41852_ & new_n42336_;
  assign new_n42338_ = ~new_n41853_ & ~new_n41856_;
  assign new_n42339_ = ~new_n42337_ & ~new_n42338_;
  assign new_n42340_ = ~new_n42038_ & ~new_n42339_;
  assign new_n42341_ = ~new_n41744_ & ~new_n42037_;
  assign new_n42342_ = ~new_n42036_ & new_n42341_;
  assign new_n42343_ = ~new_n42340_ & ~new_n42342_;
  assign new_n42344_ = ~\b[10]  & ~new_n42343_;
  assign new_n42345_ = ~new_n41763_ & new_n41851_;
  assign new_n42346_ = ~new_n41847_ & new_n42345_;
  assign new_n42347_ = ~new_n41848_ & ~new_n41851_;
  assign new_n42348_ = ~new_n42346_ & ~new_n42347_;
  assign new_n42349_ = ~new_n42038_ & ~new_n42348_;
  assign new_n42350_ = ~new_n41753_ & ~new_n42037_;
  assign new_n42351_ = ~new_n42036_ & new_n42350_;
  assign new_n42352_ = ~new_n42349_ & ~new_n42351_;
  assign new_n42353_ = ~\b[9]  & ~new_n42352_;
  assign new_n42354_ = ~new_n41772_ & new_n41846_;
  assign new_n42355_ = ~new_n41842_ & new_n42354_;
  assign new_n42356_ = ~new_n41843_ & ~new_n41846_;
  assign new_n42357_ = ~new_n42355_ & ~new_n42356_;
  assign new_n42358_ = ~new_n42038_ & ~new_n42357_;
  assign new_n42359_ = ~new_n41762_ & ~new_n42037_;
  assign new_n42360_ = ~new_n42036_ & new_n42359_;
  assign new_n42361_ = ~new_n42358_ & ~new_n42360_;
  assign new_n42362_ = ~\b[8]  & ~new_n42361_;
  assign new_n42363_ = ~new_n41781_ & new_n41841_;
  assign new_n42364_ = ~new_n41837_ & new_n42363_;
  assign new_n42365_ = ~new_n41838_ & ~new_n41841_;
  assign new_n42366_ = ~new_n42364_ & ~new_n42365_;
  assign new_n42367_ = ~new_n42038_ & ~new_n42366_;
  assign new_n42368_ = ~new_n41771_ & ~new_n42037_;
  assign new_n42369_ = ~new_n42036_ & new_n42368_;
  assign new_n42370_ = ~new_n42367_ & ~new_n42369_;
  assign new_n42371_ = ~\b[7]  & ~new_n42370_;
  assign new_n42372_ = ~new_n41790_ & new_n41836_;
  assign new_n42373_ = ~new_n41832_ & new_n42372_;
  assign new_n42374_ = ~new_n41833_ & ~new_n41836_;
  assign new_n42375_ = ~new_n42373_ & ~new_n42374_;
  assign new_n42376_ = ~new_n42038_ & ~new_n42375_;
  assign new_n42377_ = ~new_n41780_ & ~new_n42037_;
  assign new_n42378_ = ~new_n42036_ & new_n42377_;
  assign new_n42379_ = ~new_n42376_ & ~new_n42378_;
  assign new_n42380_ = ~\b[6]  & ~new_n42379_;
  assign new_n42381_ = ~new_n41799_ & new_n41831_;
  assign new_n42382_ = ~new_n41827_ & new_n42381_;
  assign new_n42383_ = ~new_n41828_ & ~new_n41831_;
  assign new_n42384_ = ~new_n42382_ & ~new_n42383_;
  assign new_n42385_ = ~new_n42038_ & ~new_n42384_;
  assign new_n42386_ = ~new_n41789_ & ~new_n42037_;
  assign new_n42387_ = ~new_n42036_ & new_n42386_;
  assign new_n42388_ = ~new_n42385_ & ~new_n42387_;
  assign new_n42389_ = ~\b[5]  & ~new_n42388_;
  assign new_n42390_ = ~new_n41807_ & new_n41826_;
  assign new_n42391_ = ~new_n41822_ & new_n42390_;
  assign new_n42392_ = ~new_n41823_ & ~new_n41826_;
  assign new_n42393_ = ~new_n42391_ & ~new_n42392_;
  assign new_n42394_ = ~new_n42038_ & ~new_n42393_;
  assign new_n42395_ = ~new_n41798_ & ~new_n42037_;
  assign new_n42396_ = ~new_n42036_ & new_n42395_;
  assign new_n42397_ = ~new_n42394_ & ~new_n42396_;
  assign new_n42398_ = ~\b[4]  & ~new_n42397_;
  assign new_n42399_ = ~new_n41817_ & new_n41821_;
  assign new_n42400_ = ~new_n41816_ & new_n42399_;
  assign new_n42401_ = ~new_n41818_ & ~new_n41821_;
  assign new_n42402_ = ~new_n42400_ & ~new_n42401_;
  assign new_n42403_ = ~new_n42038_ & ~new_n42402_;
  assign new_n42404_ = ~new_n41806_ & ~new_n42037_;
  assign new_n42405_ = ~new_n42036_ & new_n42404_;
  assign new_n42406_ = ~new_n42403_ & ~new_n42405_;
  assign new_n42407_ = ~\b[3]  & ~new_n42406_;
  assign new_n42408_ = new_n13739_ & ~new_n41814_;
  assign new_n42409_ = ~new_n41812_ & new_n42408_;
  assign new_n42410_ = ~new_n41816_ & ~new_n42409_;
  assign new_n42411_ = ~new_n42038_ & new_n42410_;
  assign new_n42412_ = ~new_n41811_ & ~new_n42037_;
  assign new_n42413_ = ~new_n42036_ & new_n42412_;
  assign new_n42414_ = ~new_n42411_ & ~new_n42413_;
  assign new_n42415_ = ~\b[2]  & ~new_n42414_;
  assign new_n42416_ = \b[0]  & ~new_n42038_;
  assign new_n42417_ = \a[20]  & ~new_n42416_;
  assign new_n42418_ = new_n13739_ & ~new_n42038_;
  assign new_n42419_ = ~new_n42417_ & ~new_n42418_;
  assign new_n42420_ = \b[1]  & ~new_n42419_;
  assign new_n42421_ = ~\b[1]  & ~new_n42418_;
  assign new_n42422_ = ~new_n42417_ & new_n42421_;
  assign new_n42423_ = ~new_n42420_ & ~new_n42422_;
  assign new_n42424_ = ~new_n14349_ & ~new_n42423_;
  assign new_n42425_ = ~\b[1]  & ~new_n42419_;
  assign new_n42426_ = ~new_n42424_ & ~new_n42425_;
  assign new_n42427_ = \b[2]  & ~new_n42413_;
  assign new_n42428_ = ~new_n42411_ & new_n42427_;
  assign new_n42429_ = ~new_n42415_ & ~new_n42428_;
  assign new_n42430_ = ~new_n42426_ & new_n42429_;
  assign new_n42431_ = ~new_n42415_ & ~new_n42430_;
  assign new_n42432_ = \b[3]  & ~new_n42405_;
  assign new_n42433_ = ~new_n42403_ & new_n42432_;
  assign new_n42434_ = ~new_n42407_ & ~new_n42433_;
  assign new_n42435_ = ~new_n42431_ & new_n42434_;
  assign new_n42436_ = ~new_n42407_ & ~new_n42435_;
  assign new_n42437_ = \b[4]  & ~new_n42396_;
  assign new_n42438_ = ~new_n42394_ & new_n42437_;
  assign new_n42439_ = ~new_n42398_ & ~new_n42438_;
  assign new_n42440_ = ~new_n42436_ & new_n42439_;
  assign new_n42441_ = ~new_n42398_ & ~new_n42440_;
  assign new_n42442_ = \b[5]  & ~new_n42387_;
  assign new_n42443_ = ~new_n42385_ & new_n42442_;
  assign new_n42444_ = ~new_n42389_ & ~new_n42443_;
  assign new_n42445_ = ~new_n42441_ & new_n42444_;
  assign new_n42446_ = ~new_n42389_ & ~new_n42445_;
  assign new_n42447_ = \b[6]  & ~new_n42378_;
  assign new_n42448_ = ~new_n42376_ & new_n42447_;
  assign new_n42449_ = ~new_n42380_ & ~new_n42448_;
  assign new_n42450_ = ~new_n42446_ & new_n42449_;
  assign new_n42451_ = ~new_n42380_ & ~new_n42450_;
  assign new_n42452_ = \b[7]  & ~new_n42369_;
  assign new_n42453_ = ~new_n42367_ & new_n42452_;
  assign new_n42454_ = ~new_n42371_ & ~new_n42453_;
  assign new_n42455_ = ~new_n42451_ & new_n42454_;
  assign new_n42456_ = ~new_n42371_ & ~new_n42455_;
  assign new_n42457_ = \b[8]  & ~new_n42360_;
  assign new_n42458_ = ~new_n42358_ & new_n42457_;
  assign new_n42459_ = ~new_n42362_ & ~new_n42458_;
  assign new_n42460_ = ~new_n42456_ & new_n42459_;
  assign new_n42461_ = ~new_n42362_ & ~new_n42460_;
  assign new_n42462_ = \b[9]  & ~new_n42351_;
  assign new_n42463_ = ~new_n42349_ & new_n42462_;
  assign new_n42464_ = ~new_n42353_ & ~new_n42463_;
  assign new_n42465_ = ~new_n42461_ & new_n42464_;
  assign new_n42466_ = ~new_n42353_ & ~new_n42465_;
  assign new_n42467_ = \b[10]  & ~new_n42342_;
  assign new_n42468_ = ~new_n42340_ & new_n42467_;
  assign new_n42469_ = ~new_n42344_ & ~new_n42468_;
  assign new_n42470_ = ~new_n42466_ & new_n42469_;
  assign new_n42471_ = ~new_n42344_ & ~new_n42470_;
  assign new_n42472_ = \b[11]  & ~new_n42333_;
  assign new_n42473_ = ~new_n42331_ & new_n42472_;
  assign new_n42474_ = ~new_n42335_ & ~new_n42473_;
  assign new_n42475_ = ~new_n42471_ & new_n42474_;
  assign new_n42476_ = ~new_n42335_ & ~new_n42475_;
  assign new_n42477_ = \b[12]  & ~new_n42324_;
  assign new_n42478_ = ~new_n42322_ & new_n42477_;
  assign new_n42479_ = ~new_n42326_ & ~new_n42478_;
  assign new_n42480_ = ~new_n42476_ & new_n42479_;
  assign new_n42481_ = ~new_n42326_ & ~new_n42480_;
  assign new_n42482_ = \b[13]  & ~new_n42315_;
  assign new_n42483_ = ~new_n42313_ & new_n42482_;
  assign new_n42484_ = ~new_n42317_ & ~new_n42483_;
  assign new_n42485_ = ~new_n42481_ & new_n42484_;
  assign new_n42486_ = ~new_n42317_ & ~new_n42485_;
  assign new_n42487_ = \b[14]  & ~new_n42306_;
  assign new_n42488_ = ~new_n42304_ & new_n42487_;
  assign new_n42489_ = ~new_n42308_ & ~new_n42488_;
  assign new_n42490_ = ~new_n42486_ & new_n42489_;
  assign new_n42491_ = ~new_n42308_ & ~new_n42490_;
  assign new_n42492_ = \b[15]  & ~new_n42297_;
  assign new_n42493_ = ~new_n42295_ & new_n42492_;
  assign new_n42494_ = ~new_n42299_ & ~new_n42493_;
  assign new_n42495_ = ~new_n42491_ & new_n42494_;
  assign new_n42496_ = ~new_n42299_ & ~new_n42495_;
  assign new_n42497_ = \b[16]  & ~new_n42288_;
  assign new_n42498_ = ~new_n42286_ & new_n42497_;
  assign new_n42499_ = ~new_n42290_ & ~new_n42498_;
  assign new_n42500_ = ~new_n42496_ & new_n42499_;
  assign new_n42501_ = ~new_n42290_ & ~new_n42500_;
  assign new_n42502_ = \b[17]  & ~new_n42279_;
  assign new_n42503_ = ~new_n42277_ & new_n42502_;
  assign new_n42504_ = ~new_n42281_ & ~new_n42503_;
  assign new_n42505_ = ~new_n42501_ & new_n42504_;
  assign new_n42506_ = ~new_n42281_ & ~new_n42505_;
  assign new_n42507_ = \b[18]  & ~new_n42270_;
  assign new_n42508_ = ~new_n42268_ & new_n42507_;
  assign new_n42509_ = ~new_n42272_ & ~new_n42508_;
  assign new_n42510_ = ~new_n42506_ & new_n42509_;
  assign new_n42511_ = ~new_n42272_ & ~new_n42510_;
  assign new_n42512_ = \b[19]  & ~new_n42261_;
  assign new_n42513_ = ~new_n42259_ & new_n42512_;
  assign new_n42514_ = ~new_n42263_ & ~new_n42513_;
  assign new_n42515_ = ~new_n42511_ & new_n42514_;
  assign new_n42516_ = ~new_n42263_ & ~new_n42515_;
  assign new_n42517_ = \b[20]  & ~new_n42252_;
  assign new_n42518_ = ~new_n42250_ & new_n42517_;
  assign new_n42519_ = ~new_n42254_ & ~new_n42518_;
  assign new_n42520_ = ~new_n42516_ & new_n42519_;
  assign new_n42521_ = ~new_n42254_ & ~new_n42520_;
  assign new_n42522_ = \b[21]  & ~new_n42243_;
  assign new_n42523_ = ~new_n42241_ & new_n42522_;
  assign new_n42524_ = ~new_n42245_ & ~new_n42523_;
  assign new_n42525_ = ~new_n42521_ & new_n42524_;
  assign new_n42526_ = ~new_n42245_ & ~new_n42525_;
  assign new_n42527_ = \b[22]  & ~new_n42234_;
  assign new_n42528_ = ~new_n42232_ & new_n42527_;
  assign new_n42529_ = ~new_n42236_ & ~new_n42528_;
  assign new_n42530_ = ~new_n42526_ & new_n42529_;
  assign new_n42531_ = ~new_n42236_ & ~new_n42530_;
  assign new_n42532_ = \b[23]  & ~new_n42225_;
  assign new_n42533_ = ~new_n42223_ & new_n42532_;
  assign new_n42534_ = ~new_n42227_ & ~new_n42533_;
  assign new_n42535_ = ~new_n42531_ & new_n42534_;
  assign new_n42536_ = ~new_n42227_ & ~new_n42535_;
  assign new_n42537_ = \b[24]  & ~new_n42216_;
  assign new_n42538_ = ~new_n42214_ & new_n42537_;
  assign new_n42539_ = ~new_n42218_ & ~new_n42538_;
  assign new_n42540_ = ~new_n42536_ & new_n42539_;
  assign new_n42541_ = ~new_n42218_ & ~new_n42540_;
  assign new_n42542_ = \b[25]  & ~new_n42207_;
  assign new_n42543_ = ~new_n42205_ & new_n42542_;
  assign new_n42544_ = ~new_n42209_ & ~new_n42543_;
  assign new_n42545_ = ~new_n42541_ & new_n42544_;
  assign new_n42546_ = ~new_n42209_ & ~new_n42545_;
  assign new_n42547_ = \b[26]  & ~new_n42198_;
  assign new_n42548_ = ~new_n42196_ & new_n42547_;
  assign new_n42549_ = ~new_n42200_ & ~new_n42548_;
  assign new_n42550_ = ~new_n42546_ & new_n42549_;
  assign new_n42551_ = ~new_n42200_ & ~new_n42550_;
  assign new_n42552_ = \b[27]  & ~new_n42189_;
  assign new_n42553_ = ~new_n42187_ & new_n42552_;
  assign new_n42554_ = ~new_n42191_ & ~new_n42553_;
  assign new_n42555_ = ~new_n42551_ & new_n42554_;
  assign new_n42556_ = ~new_n42191_ & ~new_n42555_;
  assign new_n42557_ = \b[28]  & ~new_n42180_;
  assign new_n42558_ = ~new_n42178_ & new_n42557_;
  assign new_n42559_ = ~new_n42182_ & ~new_n42558_;
  assign new_n42560_ = ~new_n42556_ & new_n42559_;
  assign new_n42561_ = ~new_n42182_ & ~new_n42560_;
  assign new_n42562_ = \b[29]  & ~new_n42171_;
  assign new_n42563_ = ~new_n42169_ & new_n42562_;
  assign new_n42564_ = ~new_n42173_ & ~new_n42563_;
  assign new_n42565_ = ~new_n42561_ & new_n42564_;
  assign new_n42566_ = ~new_n42173_ & ~new_n42565_;
  assign new_n42567_ = \b[30]  & ~new_n42162_;
  assign new_n42568_ = ~new_n42160_ & new_n42567_;
  assign new_n42569_ = ~new_n42164_ & ~new_n42568_;
  assign new_n42570_ = ~new_n42566_ & new_n42569_;
  assign new_n42571_ = ~new_n42164_ & ~new_n42570_;
  assign new_n42572_ = \b[31]  & ~new_n42153_;
  assign new_n42573_ = ~new_n42151_ & new_n42572_;
  assign new_n42574_ = ~new_n42155_ & ~new_n42573_;
  assign new_n42575_ = ~new_n42571_ & new_n42574_;
  assign new_n42576_ = ~new_n42155_ & ~new_n42575_;
  assign new_n42577_ = \b[32]  & ~new_n42144_;
  assign new_n42578_ = ~new_n42142_ & new_n42577_;
  assign new_n42579_ = ~new_n42146_ & ~new_n42578_;
  assign new_n42580_ = ~new_n42576_ & new_n42579_;
  assign new_n42581_ = ~new_n42146_ & ~new_n42580_;
  assign new_n42582_ = \b[33]  & ~new_n42135_;
  assign new_n42583_ = ~new_n42133_ & new_n42582_;
  assign new_n42584_ = ~new_n42137_ & ~new_n42583_;
  assign new_n42585_ = ~new_n42581_ & new_n42584_;
  assign new_n42586_ = ~new_n42137_ & ~new_n42585_;
  assign new_n42587_ = \b[34]  & ~new_n42126_;
  assign new_n42588_ = ~new_n42124_ & new_n42587_;
  assign new_n42589_ = ~new_n42128_ & ~new_n42588_;
  assign new_n42590_ = ~new_n42586_ & new_n42589_;
  assign new_n42591_ = ~new_n42128_ & ~new_n42590_;
  assign new_n42592_ = \b[35]  & ~new_n42117_;
  assign new_n42593_ = ~new_n42115_ & new_n42592_;
  assign new_n42594_ = ~new_n42119_ & ~new_n42593_;
  assign new_n42595_ = ~new_n42591_ & new_n42594_;
  assign new_n42596_ = ~new_n42119_ & ~new_n42595_;
  assign new_n42597_ = \b[36]  & ~new_n42108_;
  assign new_n42598_ = ~new_n42106_ & new_n42597_;
  assign new_n42599_ = ~new_n42110_ & ~new_n42598_;
  assign new_n42600_ = ~new_n42596_ & new_n42599_;
  assign new_n42601_ = ~new_n42110_ & ~new_n42600_;
  assign new_n42602_ = \b[37]  & ~new_n42099_;
  assign new_n42603_ = ~new_n42097_ & new_n42602_;
  assign new_n42604_ = ~new_n42101_ & ~new_n42603_;
  assign new_n42605_ = ~new_n42601_ & new_n42604_;
  assign new_n42606_ = ~new_n42101_ & ~new_n42605_;
  assign new_n42607_ = \b[38]  & ~new_n42090_;
  assign new_n42608_ = ~new_n42088_ & new_n42607_;
  assign new_n42609_ = ~new_n42092_ & ~new_n42608_;
  assign new_n42610_ = ~new_n42606_ & new_n42609_;
  assign new_n42611_ = ~new_n42092_ & ~new_n42610_;
  assign new_n42612_ = \b[39]  & ~new_n42081_;
  assign new_n42613_ = ~new_n42079_ & new_n42612_;
  assign new_n42614_ = ~new_n42083_ & ~new_n42613_;
  assign new_n42615_ = ~new_n42611_ & new_n42614_;
  assign new_n42616_ = ~new_n42083_ & ~new_n42615_;
  assign new_n42617_ = \b[40]  & ~new_n42072_;
  assign new_n42618_ = ~new_n42070_ & new_n42617_;
  assign new_n42619_ = ~new_n42074_ & ~new_n42618_;
  assign new_n42620_ = ~new_n42616_ & new_n42619_;
  assign new_n42621_ = ~new_n42074_ & ~new_n42620_;
  assign new_n42622_ = \b[41]  & ~new_n42063_;
  assign new_n42623_ = ~new_n42061_ & new_n42622_;
  assign new_n42624_ = ~new_n42065_ & ~new_n42623_;
  assign new_n42625_ = ~new_n42621_ & new_n42624_;
  assign new_n42626_ = ~new_n42065_ & ~new_n42625_;
  assign new_n42627_ = \b[42]  & ~new_n42054_;
  assign new_n42628_ = ~new_n42052_ & new_n42627_;
  assign new_n42629_ = ~new_n42056_ & ~new_n42628_;
  assign new_n42630_ = ~new_n42626_ & new_n42629_;
  assign new_n42631_ = ~new_n42056_ & ~new_n42630_;
  assign new_n42632_ = \b[43]  & ~new_n42045_;
  assign new_n42633_ = ~new_n42043_ & new_n42632_;
  assign new_n42634_ = ~new_n42047_ & ~new_n42633_;
  assign new_n42635_ = ~new_n42631_ & new_n42634_;
  assign new_n42636_ = ~new_n42047_ & ~new_n42635_;
  assign new_n42637_ = ~new_n41448_ & ~new_n42033_;
  assign new_n42638_ = ~new_n42031_ & new_n42637_;
  assign new_n42639_ = ~new_n42022_ & new_n42638_;
  assign new_n42640_ = ~new_n42031_ & ~new_n42033_;
  assign new_n42641_ = ~new_n42023_ & ~new_n42640_;
  assign new_n42642_ = ~new_n42639_ & ~new_n42641_;
  assign new_n42643_ = ~new_n42038_ & ~new_n42642_;
  assign new_n42644_ = ~new_n42030_ & ~new_n42037_;
  assign new_n42645_ = ~new_n42036_ & new_n42644_;
  assign new_n42646_ = ~new_n42643_ & ~new_n42645_;
  assign new_n42647_ = ~\b[44]  & ~new_n42646_;
  assign new_n42648_ = \b[44]  & ~new_n42645_;
  assign new_n42649_ = ~new_n42643_ & new_n42648_;
  assign new_n42650_ = new_n14576_ & ~new_n42649_;
  assign new_n42651_ = ~new_n42647_ & new_n42650_;
  assign new_n42652_ = ~new_n42636_ & new_n42651_;
  assign new_n42653_ = new_n13958_ & ~new_n42646_;
  assign new_n42654_ = ~new_n42652_ & ~new_n42653_;
  assign new_n42655_ = ~new_n42056_ & new_n42634_;
  assign new_n42656_ = ~new_n42630_ & new_n42655_;
  assign new_n42657_ = ~new_n42631_ & ~new_n42634_;
  assign new_n42658_ = ~new_n42656_ & ~new_n42657_;
  assign new_n42659_ = ~new_n42654_ & ~new_n42658_;
  assign new_n42660_ = ~new_n42046_ & ~new_n42653_;
  assign new_n42661_ = ~new_n42652_ & new_n42660_;
  assign new_n42662_ = ~new_n42659_ & ~new_n42661_;
  assign new_n42663_ = ~new_n42047_ & ~new_n42649_;
  assign new_n42664_ = ~new_n42647_ & new_n42663_;
  assign new_n42665_ = ~new_n42635_ & new_n42664_;
  assign new_n42666_ = ~new_n42647_ & ~new_n42649_;
  assign new_n42667_ = ~new_n42636_ & ~new_n42666_;
  assign new_n42668_ = ~new_n42665_ & ~new_n42667_;
  assign new_n42669_ = ~new_n42654_ & ~new_n42668_;
  assign new_n42670_ = ~new_n42646_ & ~new_n42653_;
  assign new_n42671_ = ~new_n42652_ & new_n42670_;
  assign new_n42672_ = ~new_n42669_ & ~new_n42671_;
  assign new_n42673_ = ~\b[45]  & ~new_n42672_;
  assign new_n42674_ = ~\b[44]  & ~new_n42662_;
  assign new_n42675_ = ~new_n42065_ & new_n42629_;
  assign new_n42676_ = ~new_n42625_ & new_n42675_;
  assign new_n42677_ = ~new_n42626_ & ~new_n42629_;
  assign new_n42678_ = ~new_n42676_ & ~new_n42677_;
  assign new_n42679_ = ~new_n42654_ & ~new_n42678_;
  assign new_n42680_ = ~new_n42055_ & ~new_n42653_;
  assign new_n42681_ = ~new_n42652_ & new_n42680_;
  assign new_n42682_ = ~new_n42679_ & ~new_n42681_;
  assign new_n42683_ = ~\b[43]  & ~new_n42682_;
  assign new_n42684_ = ~new_n42074_ & new_n42624_;
  assign new_n42685_ = ~new_n42620_ & new_n42684_;
  assign new_n42686_ = ~new_n42621_ & ~new_n42624_;
  assign new_n42687_ = ~new_n42685_ & ~new_n42686_;
  assign new_n42688_ = ~new_n42654_ & ~new_n42687_;
  assign new_n42689_ = ~new_n42064_ & ~new_n42653_;
  assign new_n42690_ = ~new_n42652_ & new_n42689_;
  assign new_n42691_ = ~new_n42688_ & ~new_n42690_;
  assign new_n42692_ = ~\b[42]  & ~new_n42691_;
  assign new_n42693_ = ~new_n42083_ & new_n42619_;
  assign new_n42694_ = ~new_n42615_ & new_n42693_;
  assign new_n42695_ = ~new_n42616_ & ~new_n42619_;
  assign new_n42696_ = ~new_n42694_ & ~new_n42695_;
  assign new_n42697_ = ~new_n42654_ & ~new_n42696_;
  assign new_n42698_ = ~new_n42073_ & ~new_n42653_;
  assign new_n42699_ = ~new_n42652_ & new_n42698_;
  assign new_n42700_ = ~new_n42697_ & ~new_n42699_;
  assign new_n42701_ = ~\b[41]  & ~new_n42700_;
  assign new_n42702_ = ~new_n42092_ & new_n42614_;
  assign new_n42703_ = ~new_n42610_ & new_n42702_;
  assign new_n42704_ = ~new_n42611_ & ~new_n42614_;
  assign new_n42705_ = ~new_n42703_ & ~new_n42704_;
  assign new_n42706_ = ~new_n42654_ & ~new_n42705_;
  assign new_n42707_ = ~new_n42082_ & ~new_n42653_;
  assign new_n42708_ = ~new_n42652_ & new_n42707_;
  assign new_n42709_ = ~new_n42706_ & ~new_n42708_;
  assign new_n42710_ = ~\b[40]  & ~new_n42709_;
  assign new_n42711_ = ~new_n42101_ & new_n42609_;
  assign new_n42712_ = ~new_n42605_ & new_n42711_;
  assign new_n42713_ = ~new_n42606_ & ~new_n42609_;
  assign new_n42714_ = ~new_n42712_ & ~new_n42713_;
  assign new_n42715_ = ~new_n42654_ & ~new_n42714_;
  assign new_n42716_ = ~new_n42091_ & ~new_n42653_;
  assign new_n42717_ = ~new_n42652_ & new_n42716_;
  assign new_n42718_ = ~new_n42715_ & ~new_n42717_;
  assign new_n42719_ = ~\b[39]  & ~new_n42718_;
  assign new_n42720_ = ~new_n42110_ & new_n42604_;
  assign new_n42721_ = ~new_n42600_ & new_n42720_;
  assign new_n42722_ = ~new_n42601_ & ~new_n42604_;
  assign new_n42723_ = ~new_n42721_ & ~new_n42722_;
  assign new_n42724_ = ~new_n42654_ & ~new_n42723_;
  assign new_n42725_ = ~new_n42100_ & ~new_n42653_;
  assign new_n42726_ = ~new_n42652_ & new_n42725_;
  assign new_n42727_ = ~new_n42724_ & ~new_n42726_;
  assign new_n42728_ = ~\b[38]  & ~new_n42727_;
  assign new_n42729_ = ~new_n42119_ & new_n42599_;
  assign new_n42730_ = ~new_n42595_ & new_n42729_;
  assign new_n42731_ = ~new_n42596_ & ~new_n42599_;
  assign new_n42732_ = ~new_n42730_ & ~new_n42731_;
  assign new_n42733_ = ~new_n42654_ & ~new_n42732_;
  assign new_n42734_ = ~new_n42109_ & ~new_n42653_;
  assign new_n42735_ = ~new_n42652_ & new_n42734_;
  assign new_n42736_ = ~new_n42733_ & ~new_n42735_;
  assign new_n42737_ = ~\b[37]  & ~new_n42736_;
  assign new_n42738_ = ~new_n42128_ & new_n42594_;
  assign new_n42739_ = ~new_n42590_ & new_n42738_;
  assign new_n42740_ = ~new_n42591_ & ~new_n42594_;
  assign new_n42741_ = ~new_n42739_ & ~new_n42740_;
  assign new_n42742_ = ~new_n42654_ & ~new_n42741_;
  assign new_n42743_ = ~new_n42118_ & ~new_n42653_;
  assign new_n42744_ = ~new_n42652_ & new_n42743_;
  assign new_n42745_ = ~new_n42742_ & ~new_n42744_;
  assign new_n42746_ = ~\b[36]  & ~new_n42745_;
  assign new_n42747_ = ~new_n42137_ & new_n42589_;
  assign new_n42748_ = ~new_n42585_ & new_n42747_;
  assign new_n42749_ = ~new_n42586_ & ~new_n42589_;
  assign new_n42750_ = ~new_n42748_ & ~new_n42749_;
  assign new_n42751_ = ~new_n42654_ & ~new_n42750_;
  assign new_n42752_ = ~new_n42127_ & ~new_n42653_;
  assign new_n42753_ = ~new_n42652_ & new_n42752_;
  assign new_n42754_ = ~new_n42751_ & ~new_n42753_;
  assign new_n42755_ = ~\b[35]  & ~new_n42754_;
  assign new_n42756_ = ~new_n42146_ & new_n42584_;
  assign new_n42757_ = ~new_n42580_ & new_n42756_;
  assign new_n42758_ = ~new_n42581_ & ~new_n42584_;
  assign new_n42759_ = ~new_n42757_ & ~new_n42758_;
  assign new_n42760_ = ~new_n42654_ & ~new_n42759_;
  assign new_n42761_ = ~new_n42136_ & ~new_n42653_;
  assign new_n42762_ = ~new_n42652_ & new_n42761_;
  assign new_n42763_ = ~new_n42760_ & ~new_n42762_;
  assign new_n42764_ = ~\b[34]  & ~new_n42763_;
  assign new_n42765_ = ~new_n42155_ & new_n42579_;
  assign new_n42766_ = ~new_n42575_ & new_n42765_;
  assign new_n42767_ = ~new_n42576_ & ~new_n42579_;
  assign new_n42768_ = ~new_n42766_ & ~new_n42767_;
  assign new_n42769_ = ~new_n42654_ & ~new_n42768_;
  assign new_n42770_ = ~new_n42145_ & ~new_n42653_;
  assign new_n42771_ = ~new_n42652_ & new_n42770_;
  assign new_n42772_ = ~new_n42769_ & ~new_n42771_;
  assign new_n42773_ = ~\b[33]  & ~new_n42772_;
  assign new_n42774_ = ~new_n42164_ & new_n42574_;
  assign new_n42775_ = ~new_n42570_ & new_n42774_;
  assign new_n42776_ = ~new_n42571_ & ~new_n42574_;
  assign new_n42777_ = ~new_n42775_ & ~new_n42776_;
  assign new_n42778_ = ~new_n42654_ & ~new_n42777_;
  assign new_n42779_ = ~new_n42154_ & ~new_n42653_;
  assign new_n42780_ = ~new_n42652_ & new_n42779_;
  assign new_n42781_ = ~new_n42778_ & ~new_n42780_;
  assign new_n42782_ = ~\b[32]  & ~new_n42781_;
  assign new_n42783_ = ~new_n42173_ & new_n42569_;
  assign new_n42784_ = ~new_n42565_ & new_n42783_;
  assign new_n42785_ = ~new_n42566_ & ~new_n42569_;
  assign new_n42786_ = ~new_n42784_ & ~new_n42785_;
  assign new_n42787_ = ~new_n42654_ & ~new_n42786_;
  assign new_n42788_ = ~new_n42163_ & ~new_n42653_;
  assign new_n42789_ = ~new_n42652_ & new_n42788_;
  assign new_n42790_ = ~new_n42787_ & ~new_n42789_;
  assign new_n42791_ = ~\b[31]  & ~new_n42790_;
  assign new_n42792_ = ~new_n42182_ & new_n42564_;
  assign new_n42793_ = ~new_n42560_ & new_n42792_;
  assign new_n42794_ = ~new_n42561_ & ~new_n42564_;
  assign new_n42795_ = ~new_n42793_ & ~new_n42794_;
  assign new_n42796_ = ~new_n42654_ & ~new_n42795_;
  assign new_n42797_ = ~new_n42172_ & ~new_n42653_;
  assign new_n42798_ = ~new_n42652_ & new_n42797_;
  assign new_n42799_ = ~new_n42796_ & ~new_n42798_;
  assign new_n42800_ = ~\b[30]  & ~new_n42799_;
  assign new_n42801_ = ~new_n42191_ & new_n42559_;
  assign new_n42802_ = ~new_n42555_ & new_n42801_;
  assign new_n42803_ = ~new_n42556_ & ~new_n42559_;
  assign new_n42804_ = ~new_n42802_ & ~new_n42803_;
  assign new_n42805_ = ~new_n42654_ & ~new_n42804_;
  assign new_n42806_ = ~new_n42181_ & ~new_n42653_;
  assign new_n42807_ = ~new_n42652_ & new_n42806_;
  assign new_n42808_ = ~new_n42805_ & ~new_n42807_;
  assign new_n42809_ = ~\b[29]  & ~new_n42808_;
  assign new_n42810_ = ~new_n42200_ & new_n42554_;
  assign new_n42811_ = ~new_n42550_ & new_n42810_;
  assign new_n42812_ = ~new_n42551_ & ~new_n42554_;
  assign new_n42813_ = ~new_n42811_ & ~new_n42812_;
  assign new_n42814_ = ~new_n42654_ & ~new_n42813_;
  assign new_n42815_ = ~new_n42190_ & ~new_n42653_;
  assign new_n42816_ = ~new_n42652_ & new_n42815_;
  assign new_n42817_ = ~new_n42814_ & ~new_n42816_;
  assign new_n42818_ = ~\b[28]  & ~new_n42817_;
  assign new_n42819_ = ~new_n42209_ & new_n42549_;
  assign new_n42820_ = ~new_n42545_ & new_n42819_;
  assign new_n42821_ = ~new_n42546_ & ~new_n42549_;
  assign new_n42822_ = ~new_n42820_ & ~new_n42821_;
  assign new_n42823_ = ~new_n42654_ & ~new_n42822_;
  assign new_n42824_ = ~new_n42199_ & ~new_n42653_;
  assign new_n42825_ = ~new_n42652_ & new_n42824_;
  assign new_n42826_ = ~new_n42823_ & ~new_n42825_;
  assign new_n42827_ = ~\b[27]  & ~new_n42826_;
  assign new_n42828_ = ~new_n42218_ & new_n42544_;
  assign new_n42829_ = ~new_n42540_ & new_n42828_;
  assign new_n42830_ = ~new_n42541_ & ~new_n42544_;
  assign new_n42831_ = ~new_n42829_ & ~new_n42830_;
  assign new_n42832_ = ~new_n42654_ & ~new_n42831_;
  assign new_n42833_ = ~new_n42208_ & ~new_n42653_;
  assign new_n42834_ = ~new_n42652_ & new_n42833_;
  assign new_n42835_ = ~new_n42832_ & ~new_n42834_;
  assign new_n42836_ = ~\b[26]  & ~new_n42835_;
  assign new_n42837_ = ~new_n42227_ & new_n42539_;
  assign new_n42838_ = ~new_n42535_ & new_n42837_;
  assign new_n42839_ = ~new_n42536_ & ~new_n42539_;
  assign new_n42840_ = ~new_n42838_ & ~new_n42839_;
  assign new_n42841_ = ~new_n42654_ & ~new_n42840_;
  assign new_n42842_ = ~new_n42217_ & ~new_n42653_;
  assign new_n42843_ = ~new_n42652_ & new_n42842_;
  assign new_n42844_ = ~new_n42841_ & ~new_n42843_;
  assign new_n42845_ = ~\b[25]  & ~new_n42844_;
  assign new_n42846_ = ~new_n42236_ & new_n42534_;
  assign new_n42847_ = ~new_n42530_ & new_n42846_;
  assign new_n42848_ = ~new_n42531_ & ~new_n42534_;
  assign new_n42849_ = ~new_n42847_ & ~new_n42848_;
  assign new_n42850_ = ~new_n42654_ & ~new_n42849_;
  assign new_n42851_ = ~new_n42226_ & ~new_n42653_;
  assign new_n42852_ = ~new_n42652_ & new_n42851_;
  assign new_n42853_ = ~new_n42850_ & ~new_n42852_;
  assign new_n42854_ = ~\b[24]  & ~new_n42853_;
  assign new_n42855_ = ~new_n42245_ & new_n42529_;
  assign new_n42856_ = ~new_n42525_ & new_n42855_;
  assign new_n42857_ = ~new_n42526_ & ~new_n42529_;
  assign new_n42858_ = ~new_n42856_ & ~new_n42857_;
  assign new_n42859_ = ~new_n42654_ & ~new_n42858_;
  assign new_n42860_ = ~new_n42235_ & ~new_n42653_;
  assign new_n42861_ = ~new_n42652_ & new_n42860_;
  assign new_n42862_ = ~new_n42859_ & ~new_n42861_;
  assign new_n42863_ = ~\b[23]  & ~new_n42862_;
  assign new_n42864_ = ~new_n42254_ & new_n42524_;
  assign new_n42865_ = ~new_n42520_ & new_n42864_;
  assign new_n42866_ = ~new_n42521_ & ~new_n42524_;
  assign new_n42867_ = ~new_n42865_ & ~new_n42866_;
  assign new_n42868_ = ~new_n42654_ & ~new_n42867_;
  assign new_n42869_ = ~new_n42244_ & ~new_n42653_;
  assign new_n42870_ = ~new_n42652_ & new_n42869_;
  assign new_n42871_ = ~new_n42868_ & ~new_n42870_;
  assign new_n42872_ = ~\b[22]  & ~new_n42871_;
  assign new_n42873_ = ~new_n42263_ & new_n42519_;
  assign new_n42874_ = ~new_n42515_ & new_n42873_;
  assign new_n42875_ = ~new_n42516_ & ~new_n42519_;
  assign new_n42876_ = ~new_n42874_ & ~new_n42875_;
  assign new_n42877_ = ~new_n42654_ & ~new_n42876_;
  assign new_n42878_ = ~new_n42253_ & ~new_n42653_;
  assign new_n42879_ = ~new_n42652_ & new_n42878_;
  assign new_n42880_ = ~new_n42877_ & ~new_n42879_;
  assign new_n42881_ = ~\b[21]  & ~new_n42880_;
  assign new_n42882_ = ~new_n42272_ & new_n42514_;
  assign new_n42883_ = ~new_n42510_ & new_n42882_;
  assign new_n42884_ = ~new_n42511_ & ~new_n42514_;
  assign new_n42885_ = ~new_n42883_ & ~new_n42884_;
  assign new_n42886_ = ~new_n42654_ & ~new_n42885_;
  assign new_n42887_ = ~new_n42262_ & ~new_n42653_;
  assign new_n42888_ = ~new_n42652_ & new_n42887_;
  assign new_n42889_ = ~new_n42886_ & ~new_n42888_;
  assign new_n42890_ = ~\b[20]  & ~new_n42889_;
  assign new_n42891_ = ~new_n42281_ & new_n42509_;
  assign new_n42892_ = ~new_n42505_ & new_n42891_;
  assign new_n42893_ = ~new_n42506_ & ~new_n42509_;
  assign new_n42894_ = ~new_n42892_ & ~new_n42893_;
  assign new_n42895_ = ~new_n42654_ & ~new_n42894_;
  assign new_n42896_ = ~new_n42271_ & ~new_n42653_;
  assign new_n42897_ = ~new_n42652_ & new_n42896_;
  assign new_n42898_ = ~new_n42895_ & ~new_n42897_;
  assign new_n42899_ = ~\b[19]  & ~new_n42898_;
  assign new_n42900_ = ~new_n42290_ & new_n42504_;
  assign new_n42901_ = ~new_n42500_ & new_n42900_;
  assign new_n42902_ = ~new_n42501_ & ~new_n42504_;
  assign new_n42903_ = ~new_n42901_ & ~new_n42902_;
  assign new_n42904_ = ~new_n42654_ & ~new_n42903_;
  assign new_n42905_ = ~new_n42280_ & ~new_n42653_;
  assign new_n42906_ = ~new_n42652_ & new_n42905_;
  assign new_n42907_ = ~new_n42904_ & ~new_n42906_;
  assign new_n42908_ = ~\b[18]  & ~new_n42907_;
  assign new_n42909_ = ~new_n42299_ & new_n42499_;
  assign new_n42910_ = ~new_n42495_ & new_n42909_;
  assign new_n42911_ = ~new_n42496_ & ~new_n42499_;
  assign new_n42912_ = ~new_n42910_ & ~new_n42911_;
  assign new_n42913_ = ~new_n42654_ & ~new_n42912_;
  assign new_n42914_ = ~new_n42289_ & ~new_n42653_;
  assign new_n42915_ = ~new_n42652_ & new_n42914_;
  assign new_n42916_ = ~new_n42913_ & ~new_n42915_;
  assign new_n42917_ = ~\b[17]  & ~new_n42916_;
  assign new_n42918_ = ~new_n42308_ & new_n42494_;
  assign new_n42919_ = ~new_n42490_ & new_n42918_;
  assign new_n42920_ = ~new_n42491_ & ~new_n42494_;
  assign new_n42921_ = ~new_n42919_ & ~new_n42920_;
  assign new_n42922_ = ~new_n42654_ & ~new_n42921_;
  assign new_n42923_ = ~new_n42298_ & ~new_n42653_;
  assign new_n42924_ = ~new_n42652_ & new_n42923_;
  assign new_n42925_ = ~new_n42922_ & ~new_n42924_;
  assign new_n42926_ = ~\b[16]  & ~new_n42925_;
  assign new_n42927_ = ~new_n42317_ & new_n42489_;
  assign new_n42928_ = ~new_n42485_ & new_n42927_;
  assign new_n42929_ = ~new_n42486_ & ~new_n42489_;
  assign new_n42930_ = ~new_n42928_ & ~new_n42929_;
  assign new_n42931_ = ~new_n42654_ & ~new_n42930_;
  assign new_n42932_ = ~new_n42307_ & ~new_n42653_;
  assign new_n42933_ = ~new_n42652_ & new_n42932_;
  assign new_n42934_ = ~new_n42931_ & ~new_n42933_;
  assign new_n42935_ = ~\b[15]  & ~new_n42934_;
  assign new_n42936_ = ~new_n42326_ & new_n42484_;
  assign new_n42937_ = ~new_n42480_ & new_n42936_;
  assign new_n42938_ = ~new_n42481_ & ~new_n42484_;
  assign new_n42939_ = ~new_n42937_ & ~new_n42938_;
  assign new_n42940_ = ~new_n42654_ & ~new_n42939_;
  assign new_n42941_ = ~new_n42316_ & ~new_n42653_;
  assign new_n42942_ = ~new_n42652_ & new_n42941_;
  assign new_n42943_ = ~new_n42940_ & ~new_n42942_;
  assign new_n42944_ = ~\b[14]  & ~new_n42943_;
  assign new_n42945_ = ~new_n42335_ & new_n42479_;
  assign new_n42946_ = ~new_n42475_ & new_n42945_;
  assign new_n42947_ = ~new_n42476_ & ~new_n42479_;
  assign new_n42948_ = ~new_n42946_ & ~new_n42947_;
  assign new_n42949_ = ~new_n42654_ & ~new_n42948_;
  assign new_n42950_ = ~new_n42325_ & ~new_n42653_;
  assign new_n42951_ = ~new_n42652_ & new_n42950_;
  assign new_n42952_ = ~new_n42949_ & ~new_n42951_;
  assign new_n42953_ = ~\b[13]  & ~new_n42952_;
  assign new_n42954_ = ~new_n42344_ & new_n42474_;
  assign new_n42955_ = ~new_n42470_ & new_n42954_;
  assign new_n42956_ = ~new_n42471_ & ~new_n42474_;
  assign new_n42957_ = ~new_n42955_ & ~new_n42956_;
  assign new_n42958_ = ~new_n42654_ & ~new_n42957_;
  assign new_n42959_ = ~new_n42334_ & ~new_n42653_;
  assign new_n42960_ = ~new_n42652_ & new_n42959_;
  assign new_n42961_ = ~new_n42958_ & ~new_n42960_;
  assign new_n42962_ = ~\b[12]  & ~new_n42961_;
  assign new_n42963_ = ~new_n42353_ & new_n42469_;
  assign new_n42964_ = ~new_n42465_ & new_n42963_;
  assign new_n42965_ = ~new_n42466_ & ~new_n42469_;
  assign new_n42966_ = ~new_n42964_ & ~new_n42965_;
  assign new_n42967_ = ~new_n42654_ & ~new_n42966_;
  assign new_n42968_ = ~new_n42343_ & ~new_n42653_;
  assign new_n42969_ = ~new_n42652_ & new_n42968_;
  assign new_n42970_ = ~new_n42967_ & ~new_n42969_;
  assign new_n42971_ = ~\b[11]  & ~new_n42970_;
  assign new_n42972_ = ~new_n42362_ & new_n42464_;
  assign new_n42973_ = ~new_n42460_ & new_n42972_;
  assign new_n42974_ = ~new_n42461_ & ~new_n42464_;
  assign new_n42975_ = ~new_n42973_ & ~new_n42974_;
  assign new_n42976_ = ~new_n42654_ & ~new_n42975_;
  assign new_n42977_ = ~new_n42352_ & ~new_n42653_;
  assign new_n42978_ = ~new_n42652_ & new_n42977_;
  assign new_n42979_ = ~new_n42976_ & ~new_n42978_;
  assign new_n42980_ = ~\b[10]  & ~new_n42979_;
  assign new_n42981_ = ~new_n42371_ & new_n42459_;
  assign new_n42982_ = ~new_n42455_ & new_n42981_;
  assign new_n42983_ = ~new_n42456_ & ~new_n42459_;
  assign new_n42984_ = ~new_n42982_ & ~new_n42983_;
  assign new_n42985_ = ~new_n42654_ & ~new_n42984_;
  assign new_n42986_ = ~new_n42361_ & ~new_n42653_;
  assign new_n42987_ = ~new_n42652_ & new_n42986_;
  assign new_n42988_ = ~new_n42985_ & ~new_n42987_;
  assign new_n42989_ = ~\b[9]  & ~new_n42988_;
  assign new_n42990_ = ~new_n42380_ & new_n42454_;
  assign new_n42991_ = ~new_n42450_ & new_n42990_;
  assign new_n42992_ = ~new_n42451_ & ~new_n42454_;
  assign new_n42993_ = ~new_n42991_ & ~new_n42992_;
  assign new_n42994_ = ~new_n42654_ & ~new_n42993_;
  assign new_n42995_ = ~new_n42370_ & ~new_n42653_;
  assign new_n42996_ = ~new_n42652_ & new_n42995_;
  assign new_n42997_ = ~new_n42994_ & ~new_n42996_;
  assign new_n42998_ = ~\b[8]  & ~new_n42997_;
  assign new_n42999_ = ~new_n42389_ & new_n42449_;
  assign new_n43000_ = ~new_n42445_ & new_n42999_;
  assign new_n43001_ = ~new_n42446_ & ~new_n42449_;
  assign new_n43002_ = ~new_n43000_ & ~new_n43001_;
  assign new_n43003_ = ~new_n42654_ & ~new_n43002_;
  assign new_n43004_ = ~new_n42379_ & ~new_n42653_;
  assign new_n43005_ = ~new_n42652_ & new_n43004_;
  assign new_n43006_ = ~new_n43003_ & ~new_n43005_;
  assign new_n43007_ = ~\b[7]  & ~new_n43006_;
  assign new_n43008_ = ~new_n42398_ & new_n42444_;
  assign new_n43009_ = ~new_n42440_ & new_n43008_;
  assign new_n43010_ = ~new_n42441_ & ~new_n42444_;
  assign new_n43011_ = ~new_n43009_ & ~new_n43010_;
  assign new_n43012_ = ~new_n42654_ & ~new_n43011_;
  assign new_n43013_ = ~new_n42388_ & ~new_n42653_;
  assign new_n43014_ = ~new_n42652_ & new_n43013_;
  assign new_n43015_ = ~new_n43012_ & ~new_n43014_;
  assign new_n43016_ = ~\b[6]  & ~new_n43015_;
  assign new_n43017_ = ~new_n42407_ & new_n42439_;
  assign new_n43018_ = ~new_n42435_ & new_n43017_;
  assign new_n43019_ = ~new_n42436_ & ~new_n42439_;
  assign new_n43020_ = ~new_n43018_ & ~new_n43019_;
  assign new_n43021_ = ~new_n42654_ & ~new_n43020_;
  assign new_n43022_ = ~new_n42397_ & ~new_n42653_;
  assign new_n43023_ = ~new_n42652_ & new_n43022_;
  assign new_n43024_ = ~new_n43021_ & ~new_n43023_;
  assign new_n43025_ = ~\b[5]  & ~new_n43024_;
  assign new_n43026_ = ~new_n42415_ & new_n42434_;
  assign new_n43027_ = ~new_n42430_ & new_n43026_;
  assign new_n43028_ = ~new_n42431_ & ~new_n42434_;
  assign new_n43029_ = ~new_n43027_ & ~new_n43028_;
  assign new_n43030_ = ~new_n42654_ & ~new_n43029_;
  assign new_n43031_ = ~new_n42406_ & ~new_n42653_;
  assign new_n43032_ = ~new_n42652_ & new_n43031_;
  assign new_n43033_ = ~new_n43030_ & ~new_n43032_;
  assign new_n43034_ = ~\b[4]  & ~new_n43033_;
  assign new_n43035_ = ~new_n42425_ & new_n42429_;
  assign new_n43036_ = ~new_n42424_ & new_n43035_;
  assign new_n43037_ = ~new_n42426_ & ~new_n42429_;
  assign new_n43038_ = ~new_n43036_ & ~new_n43037_;
  assign new_n43039_ = ~new_n42654_ & ~new_n43038_;
  assign new_n43040_ = ~new_n42414_ & ~new_n42653_;
  assign new_n43041_ = ~new_n42652_ & new_n43040_;
  assign new_n43042_ = ~new_n43039_ & ~new_n43041_;
  assign new_n43043_ = ~\b[3]  & ~new_n43042_;
  assign new_n43044_ = new_n14349_ & ~new_n42422_;
  assign new_n43045_ = ~new_n42420_ & new_n43044_;
  assign new_n43046_ = ~new_n42424_ & ~new_n43045_;
  assign new_n43047_ = ~new_n42654_ & new_n43046_;
  assign new_n43048_ = ~new_n42419_ & ~new_n42653_;
  assign new_n43049_ = ~new_n42652_ & new_n43048_;
  assign new_n43050_ = ~new_n43047_ & ~new_n43049_;
  assign new_n43051_ = ~\b[2]  & ~new_n43050_;
  assign new_n43052_ = \b[0]  & ~new_n42654_;
  assign new_n43053_ = \a[19]  & ~new_n43052_;
  assign new_n43054_ = new_n14349_ & ~new_n42654_;
  assign new_n43055_ = ~new_n43053_ & ~new_n43054_;
  assign new_n43056_ = \b[1]  & ~new_n43055_;
  assign new_n43057_ = ~\b[1]  & ~new_n43054_;
  assign new_n43058_ = ~new_n43053_ & new_n43057_;
  assign new_n43059_ = ~new_n43056_ & ~new_n43058_;
  assign new_n43060_ = ~new_n14987_ & ~new_n43059_;
  assign new_n43061_ = ~\b[1]  & ~new_n43055_;
  assign new_n43062_ = ~new_n43060_ & ~new_n43061_;
  assign new_n43063_ = \b[2]  & ~new_n43049_;
  assign new_n43064_ = ~new_n43047_ & new_n43063_;
  assign new_n43065_ = ~new_n43051_ & ~new_n43064_;
  assign new_n43066_ = ~new_n43062_ & new_n43065_;
  assign new_n43067_ = ~new_n43051_ & ~new_n43066_;
  assign new_n43068_ = \b[3]  & ~new_n43041_;
  assign new_n43069_ = ~new_n43039_ & new_n43068_;
  assign new_n43070_ = ~new_n43043_ & ~new_n43069_;
  assign new_n43071_ = ~new_n43067_ & new_n43070_;
  assign new_n43072_ = ~new_n43043_ & ~new_n43071_;
  assign new_n43073_ = \b[4]  & ~new_n43032_;
  assign new_n43074_ = ~new_n43030_ & new_n43073_;
  assign new_n43075_ = ~new_n43034_ & ~new_n43074_;
  assign new_n43076_ = ~new_n43072_ & new_n43075_;
  assign new_n43077_ = ~new_n43034_ & ~new_n43076_;
  assign new_n43078_ = \b[5]  & ~new_n43023_;
  assign new_n43079_ = ~new_n43021_ & new_n43078_;
  assign new_n43080_ = ~new_n43025_ & ~new_n43079_;
  assign new_n43081_ = ~new_n43077_ & new_n43080_;
  assign new_n43082_ = ~new_n43025_ & ~new_n43081_;
  assign new_n43083_ = \b[6]  & ~new_n43014_;
  assign new_n43084_ = ~new_n43012_ & new_n43083_;
  assign new_n43085_ = ~new_n43016_ & ~new_n43084_;
  assign new_n43086_ = ~new_n43082_ & new_n43085_;
  assign new_n43087_ = ~new_n43016_ & ~new_n43086_;
  assign new_n43088_ = \b[7]  & ~new_n43005_;
  assign new_n43089_ = ~new_n43003_ & new_n43088_;
  assign new_n43090_ = ~new_n43007_ & ~new_n43089_;
  assign new_n43091_ = ~new_n43087_ & new_n43090_;
  assign new_n43092_ = ~new_n43007_ & ~new_n43091_;
  assign new_n43093_ = \b[8]  & ~new_n42996_;
  assign new_n43094_ = ~new_n42994_ & new_n43093_;
  assign new_n43095_ = ~new_n42998_ & ~new_n43094_;
  assign new_n43096_ = ~new_n43092_ & new_n43095_;
  assign new_n43097_ = ~new_n42998_ & ~new_n43096_;
  assign new_n43098_ = \b[9]  & ~new_n42987_;
  assign new_n43099_ = ~new_n42985_ & new_n43098_;
  assign new_n43100_ = ~new_n42989_ & ~new_n43099_;
  assign new_n43101_ = ~new_n43097_ & new_n43100_;
  assign new_n43102_ = ~new_n42989_ & ~new_n43101_;
  assign new_n43103_ = \b[10]  & ~new_n42978_;
  assign new_n43104_ = ~new_n42976_ & new_n43103_;
  assign new_n43105_ = ~new_n42980_ & ~new_n43104_;
  assign new_n43106_ = ~new_n43102_ & new_n43105_;
  assign new_n43107_ = ~new_n42980_ & ~new_n43106_;
  assign new_n43108_ = \b[11]  & ~new_n42969_;
  assign new_n43109_ = ~new_n42967_ & new_n43108_;
  assign new_n43110_ = ~new_n42971_ & ~new_n43109_;
  assign new_n43111_ = ~new_n43107_ & new_n43110_;
  assign new_n43112_ = ~new_n42971_ & ~new_n43111_;
  assign new_n43113_ = \b[12]  & ~new_n42960_;
  assign new_n43114_ = ~new_n42958_ & new_n43113_;
  assign new_n43115_ = ~new_n42962_ & ~new_n43114_;
  assign new_n43116_ = ~new_n43112_ & new_n43115_;
  assign new_n43117_ = ~new_n42962_ & ~new_n43116_;
  assign new_n43118_ = \b[13]  & ~new_n42951_;
  assign new_n43119_ = ~new_n42949_ & new_n43118_;
  assign new_n43120_ = ~new_n42953_ & ~new_n43119_;
  assign new_n43121_ = ~new_n43117_ & new_n43120_;
  assign new_n43122_ = ~new_n42953_ & ~new_n43121_;
  assign new_n43123_ = \b[14]  & ~new_n42942_;
  assign new_n43124_ = ~new_n42940_ & new_n43123_;
  assign new_n43125_ = ~new_n42944_ & ~new_n43124_;
  assign new_n43126_ = ~new_n43122_ & new_n43125_;
  assign new_n43127_ = ~new_n42944_ & ~new_n43126_;
  assign new_n43128_ = \b[15]  & ~new_n42933_;
  assign new_n43129_ = ~new_n42931_ & new_n43128_;
  assign new_n43130_ = ~new_n42935_ & ~new_n43129_;
  assign new_n43131_ = ~new_n43127_ & new_n43130_;
  assign new_n43132_ = ~new_n42935_ & ~new_n43131_;
  assign new_n43133_ = \b[16]  & ~new_n42924_;
  assign new_n43134_ = ~new_n42922_ & new_n43133_;
  assign new_n43135_ = ~new_n42926_ & ~new_n43134_;
  assign new_n43136_ = ~new_n43132_ & new_n43135_;
  assign new_n43137_ = ~new_n42926_ & ~new_n43136_;
  assign new_n43138_ = \b[17]  & ~new_n42915_;
  assign new_n43139_ = ~new_n42913_ & new_n43138_;
  assign new_n43140_ = ~new_n42917_ & ~new_n43139_;
  assign new_n43141_ = ~new_n43137_ & new_n43140_;
  assign new_n43142_ = ~new_n42917_ & ~new_n43141_;
  assign new_n43143_ = \b[18]  & ~new_n42906_;
  assign new_n43144_ = ~new_n42904_ & new_n43143_;
  assign new_n43145_ = ~new_n42908_ & ~new_n43144_;
  assign new_n43146_ = ~new_n43142_ & new_n43145_;
  assign new_n43147_ = ~new_n42908_ & ~new_n43146_;
  assign new_n43148_ = \b[19]  & ~new_n42897_;
  assign new_n43149_ = ~new_n42895_ & new_n43148_;
  assign new_n43150_ = ~new_n42899_ & ~new_n43149_;
  assign new_n43151_ = ~new_n43147_ & new_n43150_;
  assign new_n43152_ = ~new_n42899_ & ~new_n43151_;
  assign new_n43153_ = \b[20]  & ~new_n42888_;
  assign new_n43154_ = ~new_n42886_ & new_n43153_;
  assign new_n43155_ = ~new_n42890_ & ~new_n43154_;
  assign new_n43156_ = ~new_n43152_ & new_n43155_;
  assign new_n43157_ = ~new_n42890_ & ~new_n43156_;
  assign new_n43158_ = \b[21]  & ~new_n42879_;
  assign new_n43159_ = ~new_n42877_ & new_n43158_;
  assign new_n43160_ = ~new_n42881_ & ~new_n43159_;
  assign new_n43161_ = ~new_n43157_ & new_n43160_;
  assign new_n43162_ = ~new_n42881_ & ~new_n43161_;
  assign new_n43163_ = \b[22]  & ~new_n42870_;
  assign new_n43164_ = ~new_n42868_ & new_n43163_;
  assign new_n43165_ = ~new_n42872_ & ~new_n43164_;
  assign new_n43166_ = ~new_n43162_ & new_n43165_;
  assign new_n43167_ = ~new_n42872_ & ~new_n43166_;
  assign new_n43168_ = \b[23]  & ~new_n42861_;
  assign new_n43169_ = ~new_n42859_ & new_n43168_;
  assign new_n43170_ = ~new_n42863_ & ~new_n43169_;
  assign new_n43171_ = ~new_n43167_ & new_n43170_;
  assign new_n43172_ = ~new_n42863_ & ~new_n43171_;
  assign new_n43173_ = \b[24]  & ~new_n42852_;
  assign new_n43174_ = ~new_n42850_ & new_n43173_;
  assign new_n43175_ = ~new_n42854_ & ~new_n43174_;
  assign new_n43176_ = ~new_n43172_ & new_n43175_;
  assign new_n43177_ = ~new_n42854_ & ~new_n43176_;
  assign new_n43178_ = \b[25]  & ~new_n42843_;
  assign new_n43179_ = ~new_n42841_ & new_n43178_;
  assign new_n43180_ = ~new_n42845_ & ~new_n43179_;
  assign new_n43181_ = ~new_n43177_ & new_n43180_;
  assign new_n43182_ = ~new_n42845_ & ~new_n43181_;
  assign new_n43183_ = \b[26]  & ~new_n42834_;
  assign new_n43184_ = ~new_n42832_ & new_n43183_;
  assign new_n43185_ = ~new_n42836_ & ~new_n43184_;
  assign new_n43186_ = ~new_n43182_ & new_n43185_;
  assign new_n43187_ = ~new_n42836_ & ~new_n43186_;
  assign new_n43188_ = \b[27]  & ~new_n42825_;
  assign new_n43189_ = ~new_n42823_ & new_n43188_;
  assign new_n43190_ = ~new_n42827_ & ~new_n43189_;
  assign new_n43191_ = ~new_n43187_ & new_n43190_;
  assign new_n43192_ = ~new_n42827_ & ~new_n43191_;
  assign new_n43193_ = \b[28]  & ~new_n42816_;
  assign new_n43194_ = ~new_n42814_ & new_n43193_;
  assign new_n43195_ = ~new_n42818_ & ~new_n43194_;
  assign new_n43196_ = ~new_n43192_ & new_n43195_;
  assign new_n43197_ = ~new_n42818_ & ~new_n43196_;
  assign new_n43198_ = \b[29]  & ~new_n42807_;
  assign new_n43199_ = ~new_n42805_ & new_n43198_;
  assign new_n43200_ = ~new_n42809_ & ~new_n43199_;
  assign new_n43201_ = ~new_n43197_ & new_n43200_;
  assign new_n43202_ = ~new_n42809_ & ~new_n43201_;
  assign new_n43203_ = \b[30]  & ~new_n42798_;
  assign new_n43204_ = ~new_n42796_ & new_n43203_;
  assign new_n43205_ = ~new_n42800_ & ~new_n43204_;
  assign new_n43206_ = ~new_n43202_ & new_n43205_;
  assign new_n43207_ = ~new_n42800_ & ~new_n43206_;
  assign new_n43208_ = \b[31]  & ~new_n42789_;
  assign new_n43209_ = ~new_n42787_ & new_n43208_;
  assign new_n43210_ = ~new_n42791_ & ~new_n43209_;
  assign new_n43211_ = ~new_n43207_ & new_n43210_;
  assign new_n43212_ = ~new_n42791_ & ~new_n43211_;
  assign new_n43213_ = \b[32]  & ~new_n42780_;
  assign new_n43214_ = ~new_n42778_ & new_n43213_;
  assign new_n43215_ = ~new_n42782_ & ~new_n43214_;
  assign new_n43216_ = ~new_n43212_ & new_n43215_;
  assign new_n43217_ = ~new_n42782_ & ~new_n43216_;
  assign new_n43218_ = \b[33]  & ~new_n42771_;
  assign new_n43219_ = ~new_n42769_ & new_n43218_;
  assign new_n43220_ = ~new_n42773_ & ~new_n43219_;
  assign new_n43221_ = ~new_n43217_ & new_n43220_;
  assign new_n43222_ = ~new_n42773_ & ~new_n43221_;
  assign new_n43223_ = \b[34]  & ~new_n42762_;
  assign new_n43224_ = ~new_n42760_ & new_n43223_;
  assign new_n43225_ = ~new_n42764_ & ~new_n43224_;
  assign new_n43226_ = ~new_n43222_ & new_n43225_;
  assign new_n43227_ = ~new_n42764_ & ~new_n43226_;
  assign new_n43228_ = \b[35]  & ~new_n42753_;
  assign new_n43229_ = ~new_n42751_ & new_n43228_;
  assign new_n43230_ = ~new_n42755_ & ~new_n43229_;
  assign new_n43231_ = ~new_n43227_ & new_n43230_;
  assign new_n43232_ = ~new_n42755_ & ~new_n43231_;
  assign new_n43233_ = \b[36]  & ~new_n42744_;
  assign new_n43234_ = ~new_n42742_ & new_n43233_;
  assign new_n43235_ = ~new_n42746_ & ~new_n43234_;
  assign new_n43236_ = ~new_n43232_ & new_n43235_;
  assign new_n43237_ = ~new_n42746_ & ~new_n43236_;
  assign new_n43238_ = \b[37]  & ~new_n42735_;
  assign new_n43239_ = ~new_n42733_ & new_n43238_;
  assign new_n43240_ = ~new_n42737_ & ~new_n43239_;
  assign new_n43241_ = ~new_n43237_ & new_n43240_;
  assign new_n43242_ = ~new_n42737_ & ~new_n43241_;
  assign new_n43243_ = \b[38]  & ~new_n42726_;
  assign new_n43244_ = ~new_n42724_ & new_n43243_;
  assign new_n43245_ = ~new_n42728_ & ~new_n43244_;
  assign new_n43246_ = ~new_n43242_ & new_n43245_;
  assign new_n43247_ = ~new_n42728_ & ~new_n43246_;
  assign new_n43248_ = \b[39]  & ~new_n42717_;
  assign new_n43249_ = ~new_n42715_ & new_n43248_;
  assign new_n43250_ = ~new_n42719_ & ~new_n43249_;
  assign new_n43251_ = ~new_n43247_ & new_n43250_;
  assign new_n43252_ = ~new_n42719_ & ~new_n43251_;
  assign new_n43253_ = \b[40]  & ~new_n42708_;
  assign new_n43254_ = ~new_n42706_ & new_n43253_;
  assign new_n43255_ = ~new_n42710_ & ~new_n43254_;
  assign new_n43256_ = ~new_n43252_ & new_n43255_;
  assign new_n43257_ = ~new_n42710_ & ~new_n43256_;
  assign new_n43258_ = \b[41]  & ~new_n42699_;
  assign new_n43259_ = ~new_n42697_ & new_n43258_;
  assign new_n43260_ = ~new_n42701_ & ~new_n43259_;
  assign new_n43261_ = ~new_n43257_ & new_n43260_;
  assign new_n43262_ = ~new_n42701_ & ~new_n43261_;
  assign new_n43263_ = \b[42]  & ~new_n42690_;
  assign new_n43264_ = ~new_n42688_ & new_n43263_;
  assign new_n43265_ = ~new_n42692_ & ~new_n43264_;
  assign new_n43266_ = ~new_n43262_ & new_n43265_;
  assign new_n43267_ = ~new_n42692_ & ~new_n43266_;
  assign new_n43268_ = \b[43]  & ~new_n42681_;
  assign new_n43269_ = ~new_n42679_ & new_n43268_;
  assign new_n43270_ = ~new_n42683_ & ~new_n43269_;
  assign new_n43271_ = ~new_n43267_ & new_n43270_;
  assign new_n43272_ = ~new_n42683_ & ~new_n43271_;
  assign new_n43273_ = \b[44]  & ~new_n42661_;
  assign new_n43274_ = ~new_n42659_ & new_n43273_;
  assign new_n43275_ = ~new_n42674_ & ~new_n43274_;
  assign new_n43276_ = ~new_n43272_ & new_n43275_;
  assign new_n43277_ = ~new_n42674_ & ~new_n43276_;
  assign new_n43278_ = \b[45]  & ~new_n42671_;
  assign new_n43279_ = ~new_n42669_ & new_n43278_;
  assign new_n43280_ = ~new_n42673_ & ~new_n43279_;
  assign new_n43281_ = ~new_n43277_ & new_n43280_;
  assign new_n43282_ = ~new_n42673_ & ~new_n43281_;
  assign new_n43283_ = new_n15212_ & ~new_n43282_;
  assign new_n43284_ = ~new_n42662_ & ~new_n43283_;
  assign new_n43285_ = ~new_n42683_ & new_n43275_;
  assign new_n43286_ = ~new_n43271_ & new_n43285_;
  assign new_n43287_ = ~new_n43272_ & ~new_n43275_;
  assign new_n43288_ = ~new_n43286_ & ~new_n43287_;
  assign new_n43289_ = new_n15212_ & ~new_n43288_;
  assign new_n43290_ = ~new_n43282_ & new_n43289_;
  assign new_n43291_ = ~new_n43284_ & ~new_n43290_;
  assign new_n43292_ = ~\b[45]  & ~new_n43291_;
  assign new_n43293_ = ~new_n42682_ & ~new_n43283_;
  assign new_n43294_ = ~new_n42692_ & new_n43270_;
  assign new_n43295_ = ~new_n43266_ & new_n43294_;
  assign new_n43296_ = ~new_n43267_ & ~new_n43270_;
  assign new_n43297_ = ~new_n43295_ & ~new_n43296_;
  assign new_n43298_ = new_n15212_ & ~new_n43297_;
  assign new_n43299_ = ~new_n43282_ & new_n43298_;
  assign new_n43300_ = ~new_n43293_ & ~new_n43299_;
  assign new_n43301_ = ~\b[44]  & ~new_n43300_;
  assign new_n43302_ = ~new_n42691_ & ~new_n43283_;
  assign new_n43303_ = ~new_n42701_ & new_n43265_;
  assign new_n43304_ = ~new_n43261_ & new_n43303_;
  assign new_n43305_ = ~new_n43262_ & ~new_n43265_;
  assign new_n43306_ = ~new_n43304_ & ~new_n43305_;
  assign new_n43307_ = new_n15212_ & ~new_n43306_;
  assign new_n43308_ = ~new_n43282_ & new_n43307_;
  assign new_n43309_ = ~new_n43302_ & ~new_n43308_;
  assign new_n43310_ = ~\b[43]  & ~new_n43309_;
  assign new_n43311_ = ~new_n42700_ & ~new_n43283_;
  assign new_n43312_ = ~new_n42710_ & new_n43260_;
  assign new_n43313_ = ~new_n43256_ & new_n43312_;
  assign new_n43314_ = ~new_n43257_ & ~new_n43260_;
  assign new_n43315_ = ~new_n43313_ & ~new_n43314_;
  assign new_n43316_ = new_n15212_ & ~new_n43315_;
  assign new_n43317_ = ~new_n43282_ & new_n43316_;
  assign new_n43318_ = ~new_n43311_ & ~new_n43317_;
  assign new_n43319_ = ~\b[42]  & ~new_n43318_;
  assign new_n43320_ = ~new_n42709_ & ~new_n43283_;
  assign new_n43321_ = ~new_n42719_ & new_n43255_;
  assign new_n43322_ = ~new_n43251_ & new_n43321_;
  assign new_n43323_ = ~new_n43252_ & ~new_n43255_;
  assign new_n43324_ = ~new_n43322_ & ~new_n43323_;
  assign new_n43325_ = new_n15212_ & ~new_n43324_;
  assign new_n43326_ = ~new_n43282_ & new_n43325_;
  assign new_n43327_ = ~new_n43320_ & ~new_n43326_;
  assign new_n43328_ = ~\b[41]  & ~new_n43327_;
  assign new_n43329_ = ~new_n42718_ & ~new_n43283_;
  assign new_n43330_ = ~new_n42728_ & new_n43250_;
  assign new_n43331_ = ~new_n43246_ & new_n43330_;
  assign new_n43332_ = ~new_n43247_ & ~new_n43250_;
  assign new_n43333_ = ~new_n43331_ & ~new_n43332_;
  assign new_n43334_ = new_n15212_ & ~new_n43333_;
  assign new_n43335_ = ~new_n43282_ & new_n43334_;
  assign new_n43336_ = ~new_n43329_ & ~new_n43335_;
  assign new_n43337_ = ~\b[40]  & ~new_n43336_;
  assign new_n43338_ = ~new_n42727_ & ~new_n43283_;
  assign new_n43339_ = ~new_n42737_ & new_n43245_;
  assign new_n43340_ = ~new_n43241_ & new_n43339_;
  assign new_n43341_ = ~new_n43242_ & ~new_n43245_;
  assign new_n43342_ = ~new_n43340_ & ~new_n43341_;
  assign new_n43343_ = new_n15212_ & ~new_n43342_;
  assign new_n43344_ = ~new_n43282_ & new_n43343_;
  assign new_n43345_ = ~new_n43338_ & ~new_n43344_;
  assign new_n43346_ = ~\b[39]  & ~new_n43345_;
  assign new_n43347_ = ~new_n42736_ & ~new_n43283_;
  assign new_n43348_ = ~new_n42746_ & new_n43240_;
  assign new_n43349_ = ~new_n43236_ & new_n43348_;
  assign new_n43350_ = ~new_n43237_ & ~new_n43240_;
  assign new_n43351_ = ~new_n43349_ & ~new_n43350_;
  assign new_n43352_ = new_n15212_ & ~new_n43351_;
  assign new_n43353_ = ~new_n43282_ & new_n43352_;
  assign new_n43354_ = ~new_n43347_ & ~new_n43353_;
  assign new_n43355_ = ~\b[38]  & ~new_n43354_;
  assign new_n43356_ = ~new_n42745_ & ~new_n43283_;
  assign new_n43357_ = ~new_n42755_ & new_n43235_;
  assign new_n43358_ = ~new_n43231_ & new_n43357_;
  assign new_n43359_ = ~new_n43232_ & ~new_n43235_;
  assign new_n43360_ = ~new_n43358_ & ~new_n43359_;
  assign new_n43361_ = new_n15212_ & ~new_n43360_;
  assign new_n43362_ = ~new_n43282_ & new_n43361_;
  assign new_n43363_ = ~new_n43356_ & ~new_n43362_;
  assign new_n43364_ = ~\b[37]  & ~new_n43363_;
  assign new_n43365_ = ~new_n42754_ & ~new_n43283_;
  assign new_n43366_ = ~new_n42764_ & new_n43230_;
  assign new_n43367_ = ~new_n43226_ & new_n43366_;
  assign new_n43368_ = ~new_n43227_ & ~new_n43230_;
  assign new_n43369_ = ~new_n43367_ & ~new_n43368_;
  assign new_n43370_ = new_n15212_ & ~new_n43369_;
  assign new_n43371_ = ~new_n43282_ & new_n43370_;
  assign new_n43372_ = ~new_n43365_ & ~new_n43371_;
  assign new_n43373_ = ~\b[36]  & ~new_n43372_;
  assign new_n43374_ = ~new_n42763_ & ~new_n43283_;
  assign new_n43375_ = ~new_n42773_ & new_n43225_;
  assign new_n43376_ = ~new_n43221_ & new_n43375_;
  assign new_n43377_ = ~new_n43222_ & ~new_n43225_;
  assign new_n43378_ = ~new_n43376_ & ~new_n43377_;
  assign new_n43379_ = new_n15212_ & ~new_n43378_;
  assign new_n43380_ = ~new_n43282_ & new_n43379_;
  assign new_n43381_ = ~new_n43374_ & ~new_n43380_;
  assign new_n43382_ = ~\b[35]  & ~new_n43381_;
  assign new_n43383_ = ~new_n42772_ & ~new_n43283_;
  assign new_n43384_ = ~new_n42782_ & new_n43220_;
  assign new_n43385_ = ~new_n43216_ & new_n43384_;
  assign new_n43386_ = ~new_n43217_ & ~new_n43220_;
  assign new_n43387_ = ~new_n43385_ & ~new_n43386_;
  assign new_n43388_ = new_n15212_ & ~new_n43387_;
  assign new_n43389_ = ~new_n43282_ & new_n43388_;
  assign new_n43390_ = ~new_n43383_ & ~new_n43389_;
  assign new_n43391_ = ~\b[34]  & ~new_n43390_;
  assign new_n43392_ = ~new_n42781_ & ~new_n43283_;
  assign new_n43393_ = ~new_n42791_ & new_n43215_;
  assign new_n43394_ = ~new_n43211_ & new_n43393_;
  assign new_n43395_ = ~new_n43212_ & ~new_n43215_;
  assign new_n43396_ = ~new_n43394_ & ~new_n43395_;
  assign new_n43397_ = new_n15212_ & ~new_n43396_;
  assign new_n43398_ = ~new_n43282_ & new_n43397_;
  assign new_n43399_ = ~new_n43392_ & ~new_n43398_;
  assign new_n43400_ = ~\b[33]  & ~new_n43399_;
  assign new_n43401_ = ~new_n42790_ & ~new_n43283_;
  assign new_n43402_ = ~new_n42800_ & new_n43210_;
  assign new_n43403_ = ~new_n43206_ & new_n43402_;
  assign new_n43404_ = ~new_n43207_ & ~new_n43210_;
  assign new_n43405_ = ~new_n43403_ & ~new_n43404_;
  assign new_n43406_ = new_n15212_ & ~new_n43405_;
  assign new_n43407_ = ~new_n43282_ & new_n43406_;
  assign new_n43408_ = ~new_n43401_ & ~new_n43407_;
  assign new_n43409_ = ~\b[32]  & ~new_n43408_;
  assign new_n43410_ = ~new_n42799_ & ~new_n43283_;
  assign new_n43411_ = ~new_n42809_ & new_n43205_;
  assign new_n43412_ = ~new_n43201_ & new_n43411_;
  assign new_n43413_ = ~new_n43202_ & ~new_n43205_;
  assign new_n43414_ = ~new_n43412_ & ~new_n43413_;
  assign new_n43415_ = new_n15212_ & ~new_n43414_;
  assign new_n43416_ = ~new_n43282_ & new_n43415_;
  assign new_n43417_ = ~new_n43410_ & ~new_n43416_;
  assign new_n43418_ = ~\b[31]  & ~new_n43417_;
  assign new_n43419_ = ~new_n42808_ & ~new_n43283_;
  assign new_n43420_ = ~new_n42818_ & new_n43200_;
  assign new_n43421_ = ~new_n43196_ & new_n43420_;
  assign new_n43422_ = ~new_n43197_ & ~new_n43200_;
  assign new_n43423_ = ~new_n43421_ & ~new_n43422_;
  assign new_n43424_ = new_n15212_ & ~new_n43423_;
  assign new_n43425_ = ~new_n43282_ & new_n43424_;
  assign new_n43426_ = ~new_n43419_ & ~new_n43425_;
  assign new_n43427_ = ~\b[30]  & ~new_n43426_;
  assign new_n43428_ = ~new_n42817_ & ~new_n43283_;
  assign new_n43429_ = ~new_n42827_ & new_n43195_;
  assign new_n43430_ = ~new_n43191_ & new_n43429_;
  assign new_n43431_ = ~new_n43192_ & ~new_n43195_;
  assign new_n43432_ = ~new_n43430_ & ~new_n43431_;
  assign new_n43433_ = new_n15212_ & ~new_n43432_;
  assign new_n43434_ = ~new_n43282_ & new_n43433_;
  assign new_n43435_ = ~new_n43428_ & ~new_n43434_;
  assign new_n43436_ = ~\b[29]  & ~new_n43435_;
  assign new_n43437_ = ~new_n42826_ & ~new_n43283_;
  assign new_n43438_ = ~new_n42836_ & new_n43190_;
  assign new_n43439_ = ~new_n43186_ & new_n43438_;
  assign new_n43440_ = ~new_n43187_ & ~new_n43190_;
  assign new_n43441_ = ~new_n43439_ & ~new_n43440_;
  assign new_n43442_ = new_n15212_ & ~new_n43441_;
  assign new_n43443_ = ~new_n43282_ & new_n43442_;
  assign new_n43444_ = ~new_n43437_ & ~new_n43443_;
  assign new_n43445_ = ~\b[28]  & ~new_n43444_;
  assign new_n43446_ = ~new_n42835_ & ~new_n43283_;
  assign new_n43447_ = ~new_n42845_ & new_n43185_;
  assign new_n43448_ = ~new_n43181_ & new_n43447_;
  assign new_n43449_ = ~new_n43182_ & ~new_n43185_;
  assign new_n43450_ = ~new_n43448_ & ~new_n43449_;
  assign new_n43451_ = new_n15212_ & ~new_n43450_;
  assign new_n43452_ = ~new_n43282_ & new_n43451_;
  assign new_n43453_ = ~new_n43446_ & ~new_n43452_;
  assign new_n43454_ = ~\b[27]  & ~new_n43453_;
  assign new_n43455_ = ~new_n42844_ & ~new_n43283_;
  assign new_n43456_ = ~new_n42854_ & new_n43180_;
  assign new_n43457_ = ~new_n43176_ & new_n43456_;
  assign new_n43458_ = ~new_n43177_ & ~new_n43180_;
  assign new_n43459_ = ~new_n43457_ & ~new_n43458_;
  assign new_n43460_ = new_n15212_ & ~new_n43459_;
  assign new_n43461_ = ~new_n43282_ & new_n43460_;
  assign new_n43462_ = ~new_n43455_ & ~new_n43461_;
  assign new_n43463_ = ~\b[26]  & ~new_n43462_;
  assign new_n43464_ = ~new_n42853_ & ~new_n43283_;
  assign new_n43465_ = ~new_n42863_ & new_n43175_;
  assign new_n43466_ = ~new_n43171_ & new_n43465_;
  assign new_n43467_ = ~new_n43172_ & ~new_n43175_;
  assign new_n43468_ = ~new_n43466_ & ~new_n43467_;
  assign new_n43469_ = new_n15212_ & ~new_n43468_;
  assign new_n43470_ = ~new_n43282_ & new_n43469_;
  assign new_n43471_ = ~new_n43464_ & ~new_n43470_;
  assign new_n43472_ = ~\b[25]  & ~new_n43471_;
  assign new_n43473_ = ~new_n42862_ & ~new_n43283_;
  assign new_n43474_ = ~new_n42872_ & new_n43170_;
  assign new_n43475_ = ~new_n43166_ & new_n43474_;
  assign new_n43476_ = ~new_n43167_ & ~new_n43170_;
  assign new_n43477_ = ~new_n43475_ & ~new_n43476_;
  assign new_n43478_ = new_n15212_ & ~new_n43477_;
  assign new_n43479_ = ~new_n43282_ & new_n43478_;
  assign new_n43480_ = ~new_n43473_ & ~new_n43479_;
  assign new_n43481_ = ~\b[24]  & ~new_n43480_;
  assign new_n43482_ = ~new_n42871_ & ~new_n43283_;
  assign new_n43483_ = ~new_n42881_ & new_n43165_;
  assign new_n43484_ = ~new_n43161_ & new_n43483_;
  assign new_n43485_ = ~new_n43162_ & ~new_n43165_;
  assign new_n43486_ = ~new_n43484_ & ~new_n43485_;
  assign new_n43487_ = new_n15212_ & ~new_n43486_;
  assign new_n43488_ = ~new_n43282_ & new_n43487_;
  assign new_n43489_ = ~new_n43482_ & ~new_n43488_;
  assign new_n43490_ = ~\b[23]  & ~new_n43489_;
  assign new_n43491_ = ~new_n42880_ & ~new_n43283_;
  assign new_n43492_ = ~new_n42890_ & new_n43160_;
  assign new_n43493_ = ~new_n43156_ & new_n43492_;
  assign new_n43494_ = ~new_n43157_ & ~new_n43160_;
  assign new_n43495_ = ~new_n43493_ & ~new_n43494_;
  assign new_n43496_ = new_n15212_ & ~new_n43495_;
  assign new_n43497_ = ~new_n43282_ & new_n43496_;
  assign new_n43498_ = ~new_n43491_ & ~new_n43497_;
  assign new_n43499_ = ~\b[22]  & ~new_n43498_;
  assign new_n43500_ = ~new_n42889_ & ~new_n43283_;
  assign new_n43501_ = ~new_n42899_ & new_n43155_;
  assign new_n43502_ = ~new_n43151_ & new_n43501_;
  assign new_n43503_ = ~new_n43152_ & ~new_n43155_;
  assign new_n43504_ = ~new_n43502_ & ~new_n43503_;
  assign new_n43505_ = new_n15212_ & ~new_n43504_;
  assign new_n43506_ = ~new_n43282_ & new_n43505_;
  assign new_n43507_ = ~new_n43500_ & ~new_n43506_;
  assign new_n43508_ = ~\b[21]  & ~new_n43507_;
  assign new_n43509_ = ~new_n42898_ & ~new_n43283_;
  assign new_n43510_ = ~new_n42908_ & new_n43150_;
  assign new_n43511_ = ~new_n43146_ & new_n43510_;
  assign new_n43512_ = ~new_n43147_ & ~new_n43150_;
  assign new_n43513_ = ~new_n43511_ & ~new_n43512_;
  assign new_n43514_ = new_n15212_ & ~new_n43513_;
  assign new_n43515_ = ~new_n43282_ & new_n43514_;
  assign new_n43516_ = ~new_n43509_ & ~new_n43515_;
  assign new_n43517_ = ~\b[20]  & ~new_n43516_;
  assign new_n43518_ = ~new_n42907_ & ~new_n43283_;
  assign new_n43519_ = ~new_n42917_ & new_n43145_;
  assign new_n43520_ = ~new_n43141_ & new_n43519_;
  assign new_n43521_ = ~new_n43142_ & ~new_n43145_;
  assign new_n43522_ = ~new_n43520_ & ~new_n43521_;
  assign new_n43523_ = new_n15212_ & ~new_n43522_;
  assign new_n43524_ = ~new_n43282_ & new_n43523_;
  assign new_n43525_ = ~new_n43518_ & ~new_n43524_;
  assign new_n43526_ = ~\b[19]  & ~new_n43525_;
  assign new_n43527_ = ~new_n42916_ & ~new_n43283_;
  assign new_n43528_ = ~new_n42926_ & new_n43140_;
  assign new_n43529_ = ~new_n43136_ & new_n43528_;
  assign new_n43530_ = ~new_n43137_ & ~new_n43140_;
  assign new_n43531_ = ~new_n43529_ & ~new_n43530_;
  assign new_n43532_ = new_n15212_ & ~new_n43531_;
  assign new_n43533_ = ~new_n43282_ & new_n43532_;
  assign new_n43534_ = ~new_n43527_ & ~new_n43533_;
  assign new_n43535_ = ~\b[18]  & ~new_n43534_;
  assign new_n43536_ = ~new_n42925_ & ~new_n43283_;
  assign new_n43537_ = ~new_n42935_ & new_n43135_;
  assign new_n43538_ = ~new_n43131_ & new_n43537_;
  assign new_n43539_ = ~new_n43132_ & ~new_n43135_;
  assign new_n43540_ = ~new_n43538_ & ~new_n43539_;
  assign new_n43541_ = new_n15212_ & ~new_n43540_;
  assign new_n43542_ = ~new_n43282_ & new_n43541_;
  assign new_n43543_ = ~new_n43536_ & ~new_n43542_;
  assign new_n43544_ = ~\b[17]  & ~new_n43543_;
  assign new_n43545_ = ~new_n42934_ & ~new_n43283_;
  assign new_n43546_ = ~new_n42944_ & new_n43130_;
  assign new_n43547_ = ~new_n43126_ & new_n43546_;
  assign new_n43548_ = ~new_n43127_ & ~new_n43130_;
  assign new_n43549_ = ~new_n43547_ & ~new_n43548_;
  assign new_n43550_ = new_n15212_ & ~new_n43549_;
  assign new_n43551_ = ~new_n43282_ & new_n43550_;
  assign new_n43552_ = ~new_n43545_ & ~new_n43551_;
  assign new_n43553_ = ~\b[16]  & ~new_n43552_;
  assign new_n43554_ = ~new_n42943_ & ~new_n43283_;
  assign new_n43555_ = ~new_n42953_ & new_n43125_;
  assign new_n43556_ = ~new_n43121_ & new_n43555_;
  assign new_n43557_ = ~new_n43122_ & ~new_n43125_;
  assign new_n43558_ = ~new_n43556_ & ~new_n43557_;
  assign new_n43559_ = new_n15212_ & ~new_n43558_;
  assign new_n43560_ = ~new_n43282_ & new_n43559_;
  assign new_n43561_ = ~new_n43554_ & ~new_n43560_;
  assign new_n43562_ = ~\b[15]  & ~new_n43561_;
  assign new_n43563_ = ~new_n42952_ & ~new_n43283_;
  assign new_n43564_ = ~new_n42962_ & new_n43120_;
  assign new_n43565_ = ~new_n43116_ & new_n43564_;
  assign new_n43566_ = ~new_n43117_ & ~new_n43120_;
  assign new_n43567_ = ~new_n43565_ & ~new_n43566_;
  assign new_n43568_ = new_n15212_ & ~new_n43567_;
  assign new_n43569_ = ~new_n43282_ & new_n43568_;
  assign new_n43570_ = ~new_n43563_ & ~new_n43569_;
  assign new_n43571_ = ~\b[14]  & ~new_n43570_;
  assign new_n43572_ = ~new_n42961_ & ~new_n43283_;
  assign new_n43573_ = ~new_n42971_ & new_n43115_;
  assign new_n43574_ = ~new_n43111_ & new_n43573_;
  assign new_n43575_ = ~new_n43112_ & ~new_n43115_;
  assign new_n43576_ = ~new_n43574_ & ~new_n43575_;
  assign new_n43577_ = new_n15212_ & ~new_n43576_;
  assign new_n43578_ = ~new_n43282_ & new_n43577_;
  assign new_n43579_ = ~new_n43572_ & ~new_n43578_;
  assign new_n43580_ = ~\b[13]  & ~new_n43579_;
  assign new_n43581_ = ~new_n42970_ & ~new_n43283_;
  assign new_n43582_ = ~new_n42980_ & new_n43110_;
  assign new_n43583_ = ~new_n43106_ & new_n43582_;
  assign new_n43584_ = ~new_n43107_ & ~new_n43110_;
  assign new_n43585_ = ~new_n43583_ & ~new_n43584_;
  assign new_n43586_ = new_n15212_ & ~new_n43585_;
  assign new_n43587_ = ~new_n43282_ & new_n43586_;
  assign new_n43588_ = ~new_n43581_ & ~new_n43587_;
  assign new_n43589_ = ~\b[12]  & ~new_n43588_;
  assign new_n43590_ = ~new_n42979_ & ~new_n43283_;
  assign new_n43591_ = ~new_n42989_ & new_n43105_;
  assign new_n43592_ = ~new_n43101_ & new_n43591_;
  assign new_n43593_ = ~new_n43102_ & ~new_n43105_;
  assign new_n43594_ = ~new_n43592_ & ~new_n43593_;
  assign new_n43595_ = new_n15212_ & ~new_n43594_;
  assign new_n43596_ = ~new_n43282_ & new_n43595_;
  assign new_n43597_ = ~new_n43590_ & ~new_n43596_;
  assign new_n43598_ = ~\b[11]  & ~new_n43597_;
  assign new_n43599_ = ~new_n42988_ & ~new_n43283_;
  assign new_n43600_ = ~new_n42998_ & new_n43100_;
  assign new_n43601_ = ~new_n43096_ & new_n43600_;
  assign new_n43602_ = ~new_n43097_ & ~new_n43100_;
  assign new_n43603_ = ~new_n43601_ & ~new_n43602_;
  assign new_n43604_ = new_n15212_ & ~new_n43603_;
  assign new_n43605_ = ~new_n43282_ & new_n43604_;
  assign new_n43606_ = ~new_n43599_ & ~new_n43605_;
  assign new_n43607_ = ~\b[10]  & ~new_n43606_;
  assign new_n43608_ = ~new_n42997_ & ~new_n43283_;
  assign new_n43609_ = ~new_n43007_ & new_n43095_;
  assign new_n43610_ = ~new_n43091_ & new_n43609_;
  assign new_n43611_ = ~new_n43092_ & ~new_n43095_;
  assign new_n43612_ = ~new_n43610_ & ~new_n43611_;
  assign new_n43613_ = new_n15212_ & ~new_n43612_;
  assign new_n43614_ = ~new_n43282_ & new_n43613_;
  assign new_n43615_ = ~new_n43608_ & ~new_n43614_;
  assign new_n43616_ = ~\b[9]  & ~new_n43615_;
  assign new_n43617_ = ~new_n43006_ & ~new_n43283_;
  assign new_n43618_ = ~new_n43016_ & new_n43090_;
  assign new_n43619_ = ~new_n43086_ & new_n43618_;
  assign new_n43620_ = ~new_n43087_ & ~new_n43090_;
  assign new_n43621_ = ~new_n43619_ & ~new_n43620_;
  assign new_n43622_ = new_n15212_ & ~new_n43621_;
  assign new_n43623_ = ~new_n43282_ & new_n43622_;
  assign new_n43624_ = ~new_n43617_ & ~new_n43623_;
  assign new_n43625_ = ~\b[8]  & ~new_n43624_;
  assign new_n43626_ = ~new_n43015_ & ~new_n43283_;
  assign new_n43627_ = ~new_n43025_ & new_n43085_;
  assign new_n43628_ = ~new_n43081_ & new_n43627_;
  assign new_n43629_ = ~new_n43082_ & ~new_n43085_;
  assign new_n43630_ = ~new_n43628_ & ~new_n43629_;
  assign new_n43631_ = new_n15212_ & ~new_n43630_;
  assign new_n43632_ = ~new_n43282_ & new_n43631_;
  assign new_n43633_ = ~new_n43626_ & ~new_n43632_;
  assign new_n43634_ = ~\b[7]  & ~new_n43633_;
  assign new_n43635_ = ~new_n43024_ & ~new_n43283_;
  assign new_n43636_ = ~new_n43034_ & new_n43080_;
  assign new_n43637_ = ~new_n43076_ & new_n43636_;
  assign new_n43638_ = ~new_n43077_ & ~new_n43080_;
  assign new_n43639_ = ~new_n43637_ & ~new_n43638_;
  assign new_n43640_ = new_n15212_ & ~new_n43639_;
  assign new_n43641_ = ~new_n43282_ & new_n43640_;
  assign new_n43642_ = ~new_n43635_ & ~new_n43641_;
  assign new_n43643_ = ~\b[6]  & ~new_n43642_;
  assign new_n43644_ = ~new_n43033_ & ~new_n43283_;
  assign new_n43645_ = ~new_n43043_ & new_n43075_;
  assign new_n43646_ = ~new_n43071_ & new_n43645_;
  assign new_n43647_ = ~new_n43072_ & ~new_n43075_;
  assign new_n43648_ = ~new_n43646_ & ~new_n43647_;
  assign new_n43649_ = new_n15212_ & ~new_n43648_;
  assign new_n43650_ = ~new_n43282_ & new_n43649_;
  assign new_n43651_ = ~new_n43644_ & ~new_n43650_;
  assign new_n43652_ = ~\b[5]  & ~new_n43651_;
  assign new_n43653_ = ~new_n43042_ & ~new_n43283_;
  assign new_n43654_ = ~new_n43051_ & new_n43070_;
  assign new_n43655_ = ~new_n43066_ & new_n43654_;
  assign new_n43656_ = ~new_n43067_ & ~new_n43070_;
  assign new_n43657_ = ~new_n43655_ & ~new_n43656_;
  assign new_n43658_ = new_n15212_ & ~new_n43657_;
  assign new_n43659_ = ~new_n43282_ & new_n43658_;
  assign new_n43660_ = ~new_n43653_ & ~new_n43659_;
  assign new_n43661_ = ~\b[4]  & ~new_n43660_;
  assign new_n43662_ = ~new_n43050_ & ~new_n43283_;
  assign new_n43663_ = ~new_n43061_ & new_n43065_;
  assign new_n43664_ = ~new_n43060_ & new_n43663_;
  assign new_n43665_ = ~new_n43062_ & ~new_n43065_;
  assign new_n43666_ = ~new_n43664_ & ~new_n43665_;
  assign new_n43667_ = new_n15212_ & ~new_n43666_;
  assign new_n43668_ = ~new_n43282_ & new_n43667_;
  assign new_n43669_ = ~new_n43662_ & ~new_n43668_;
  assign new_n43670_ = ~\b[3]  & ~new_n43669_;
  assign new_n43671_ = ~new_n43055_ & ~new_n43283_;
  assign new_n43672_ = new_n14987_ & ~new_n43058_;
  assign new_n43673_ = ~new_n43056_ & new_n43672_;
  assign new_n43674_ = new_n15212_ & ~new_n43673_;
  assign new_n43675_ = ~new_n43060_ & new_n43674_;
  assign new_n43676_ = ~new_n43282_ & new_n43675_;
  assign new_n43677_ = ~new_n43671_ & ~new_n43676_;
  assign new_n43678_ = ~\b[2]  & ~new_n43677_;
  assign new_n43679_ = new_n15612_ & ~new_n43282_;
  assign new_n43680_ = \a[18]  & ~new_n43679_;
  assign new_n43681_ = new_n15617_ & ~new_n43282_;
  assign new_n43682_ = ~new_n43680_ & ~new_n43681_;
  assign new_n43683_ = \b[1]  & ~new_n43682_;
  assign new_n43684_ = ~\b[1]  & ~new_n43681_;
  assign new_n43685_ = ~new_n43680_ & new_n43684_;
  assign new_n43686_ = ~new_n43683_ & ~new_n43685_;
  assign new_n43687_ = ~new_n15624_ & ~new_n43686_;
  assign new_n43688_ = ~\b[1]  & ~new_n43682_;
  assign new_n43689_ = ~new_n43687_ & ~new_n43688_;
  assign new_n43690_ = \b[2]  & ~new_n43676_;
  assign new_n43691_ = ~new_n43671_ & new_n43690_;
  assign new_n43692_ = ~new_n43678_ & ~new_n43691_;
  assign new_n43693_ = ~new_n43689_ & new_n43692_;
  assign new_n43694_ = ~new_n43678_ & ~new_n43693_;
  assign new_n43695_ = \b[3]  & ~new_n43668_;
  assign new_n43696_ = ~new_n43662_ & new_n43695_;
  assign new_n43697_ = ~new_n43670_ & ~new_n43696_;
  assign new_n43698_ = ~new_n43694_ & new_n43697_;
  assign new_n43699_ = ~new_n43670_ & ~new_n43698_;
  assign new_n43700_ = \b[4]  & ~new_n43659_;
  assign new_n43701_ = ~new_n43653_ & new_n43700_;
  assign new_n43702_ = ~new_n43661_ & ~new_n43701_;
  assign new_n43703_ = ~new_n43699_ & new_n43702_;
  assign new_n43704_ = ~new_n43661_ & ~new_n43703_;
  assign new_n43705_ = \b[5]  & ~new_n43650_;
  assign new_n43706_ = ~new_n43644_ & new_n43705_;
  assign new_n43707_ = ~new_n43652_ & ~new_n43706_;
  assign new_n43708_ = ~new_n43704_ & new_n43707_;
  assign new_n43709_ = ~new_n43652_ & ~new_n43708_;
  assign new_n43710_ = \b[6]  & ~new_n43641_;
  assign new_n43711_ = ~new_n43635_ & new_n43710_;
  assign new_n43712_ = ~new_n43643_ & ~new_n43711_;
  assign new_n43713_ = ~new_n43709_ & new_n43712_;
  assign new_n43714_ = ~new_n43643_ & ~new_n43713_;
  assign new_n43715_ = \b[7]  & ~new_n43632_;
  assign new_n43716_ = ~new_n43626_ & new_n43715_;
  assign new_n43717_ = ~new_n43634_ & ~new_n43716_;
  assign new_n43718_ = ~new_n43714_ & new_n43717_;
  assign new_n43719_ = ~new_n43634_ & ~new_n43718_;
  assign new_n43720_ = \b[8]  & ~new_n43623_;
  assign new_n43721_ = ~new_n43617_ & new_n43720_;
  assign new_n43722_ = ~new_n43625_ & ~new_n43721_;
  assign new_n43723_ = ~new_n43719_ & new_n43722_;
  assign new_n43724_ = ~new_n43625_ & ~new_n43723_;
  assign new_n43725_ = \b[9]  & ~new_n43614_;
  assign new_n43726_ = ~new_n43608_ & new_n43725_;
  assign new_n43727_ = ~new_n43616_ & ~new_n43726_;
  assign new_n43728_ = ~new_n43724_ & new_n43727_;
  assign new_n43729_ = ~new_n43616_ & ~new_n43728_;
  assign new_n43730_ = \b[10]  & ~new_n43605_;
  assign new_n43731_ = ~new_n43599_ & new_n43730_;
  assign new_n43732_ = ~new_n43607_ & ~new_n43731_;
  assign new_n43733_ = ~new_n43729_ & new_n43732_;
  assign new_n43734_ = ~new_n43607_ & ~new_n43733_;
  assign new_n43735_ = \b[11]  & ~new_n43596_;
  assign new_n43736_ = ~new_n43590_ & new_n43735_;
  assign new_n43737_ = ~new_n43598_ & ~new_n43736_;
  assign new_n43738_ = ~new_n43734_ & new_n43737_;
  assign new_n43739_ = ~new_n43598_ & ~new_n43738_;
  assign new_n43740_ = \b[12]  & ~new_n43587_;
  assign new_n43741_ = ~new_n43581_ & new_n43740_;
  assign new_n43742_ = ~new_n43589_ & ~new_n43741_;
  assign new_n43743_ = ~new_n43739_ & new_n43742_;
  assign new_n43744_ = ~new_n43589_ & ~new_n43743_;
  assign new_n43745_ = \b[13]  & ~new_n43578_;
  assign new_n43746_ = ~new_n43572_ & new_n43745_;
  assign new_n43747_ = ~new_n43580_ & ~new_n43746_;
  assign new_n43748_ = ~new_n43744_ & new_n43747_;
  assign new_n43749_ = ~new_n43580_ & ~new_n43748_;
  assign new_n43750_ = \b[14]  & ~new_n43569_;
  assign new_n43751_ = ~new_n43563_ & new_n43750_;
  assign new_n43752_ = ~new_n43571_ & ~new_n43751_;
  assign new_n43753_ = ~new_n43749_ & new_n43752_;
  assign new_n43754_ = ~new_n43571_ & ~new_n43753_;
  assign new_n43755_ = \b[15]  & ~new_n43560_;
  assign new_n43756_ = ~new_n43554_ & new_n43755_;
  assign new_n43757_ = ~new_n43562_ & ~new_n43756_;
  assign new_n43758_ = ~new_n43754_ & new_n43757_;
  assign new_n43759_ = ~new_n43562_ & ~new_n43758_;
  assign new_n43760_ = \b[16]  & ~new_n43551_;
  assign new_n43761_ = ~new_n43545_ & new_n43760_;
  assign new_n43762_ = ~new_n43553_ & ~new_n43761_;
  assign new_n43763_ = ~new_n43759_ & new_n43762_;
  assign new_n43764_ = ~new_n43553_ & ~new_n43763_;
  assign new_n43765_ = \b[17]  & ~new_n43542_;
  assign new_n43766_ = ~new_n43536_ & new_n43765_;
  assign new_n43767_ = ~new_n43544_ & ~new_n43766_;
  assign new_n43768_ = ~new_n43764_ & new_n43767_;
  assign new_n43769_ = ~new_n43544_ & ~new_n43768_;
  assign new_n43770_ = \b[18]  & ~new_n43533_;
  assign new_n43771_ = ~new_n43527_ & new_n43770_;
  assign new_n43772_ = ~new_n43535_ & ~new_n43771_;
  assign new_n43773_ = ~new_n43769_ & new_n43772_;
  assign new_n43774_ = ~new_n43535_ & ~new_n43773_;
  assign new_n43775_ = \b[19]  & ~new_n43524_;
  assign new_n43776_ = ~new_n43518_ & new_n43775_;
  assign new_n43777_ = ~new_n43526_ & ~new_n43776_;
  assign new_n43778_ = ~new_n43774_ & new_n43777_;
  assign new_n43779_ = ~new_n43526_ & ~new_n43778_;
  assign new_n43780_ = \b[20]  & ~new_n43515_;
  assign new_n43781_ = ~new_n43509_ & new_n43780_;
  assign new_n43782_ = ~new_n43517_ & ~new_n43781_;
  assign new_n43783_ = ~new_n43779_ & new_n43782_;
  assign new_n43784_ = ~new_n43517_ & ~new_n43783_;
  assign new_n43785_ = \b[21]  & ~new_n43506_;
  assign new_n43786_ = ~new_n43500_ & new_n43785_;
  assign new_n43787_ = ~new_n43508_ & ~new_n43786_;
  assign new_n43788_ = ~new_n43784_ & new_n43787_;
  assign new_n43789_ = ~new_n43508_ & ~new_n43788_;
  assign new_n43790_ = \b[22]  & ~new_n43497_;
  assign new_n43791_ = ~new_n43491_ & new_n43790_;
  assign new_n43792_ = ~new_n43499_ & ~new_n43791_;
  assign new_n43793_ = ~new_n43789_ & new_n43792_;
  assign new_n43794_ = ~new_n43499_ & ~new_n43793_;
  assign new_n43795_ = \b[23]  & ~new_n43488_;
  assign new_n43796_ = ~new_n43482_ & new_n43795_;
  assign new_n43797_ = ~new_n43490_ & ~new_n43796_;
  assign new_n43798_ = ~new_n43794_ & new_n43797_;
  assign new_n43799_ = ~new_n43490_ & ~new_n43798_;
  assign new_n43800_ = \b[24]  & ~new_n43479_;
  assign new_n43801_ = ~new_n43473_ & new_n43800_;
  assign new_n43802_ = ~new_n43481_ & ~new_n43801_;
  assign new_n43803_ = ~new_n43799_ & new_n43802_;
  assign new_n43804_ = ~new_n43481_ & ~new_n43803_;
  assign new_n43805_ = \b[25]  & ~new_n43470_;
  assign new_n43806_ = ~new_n43464_ & new_n43805_;
  assign new_n43807_ = ~new_n43472_ & ~new_n43806_;
  assign new_n43808_ = ~new_n43804_ & new_n43807_;
  assign new_n43809_ = ~new_n43472_ & ~new_n43808_;
  assign new_n43810_ = \b[26]  & ~new_n43461_;
  assign new_n43811_ = ~new_n43455_ & new_n43810_;
  assign new_n43812_ = ~new_n43463_ & ~new_n43811_;
  assign new_n43813_ = ~new_n43809_ & new_n43812_;
  assign new_n43814_ = ~new_n43463_ & ~new_n43813_;
  assign new_n43815_ = \b[27]  & ~new_n43452_;
  assign new_n43816_ = ~new_n43446_ & new_n43815_;
  assign new_n43817_ = ~new_n43454_ & ~new_n43816_;
  assign new_n43818_ = ~new_n43814_ & new_n43817_;
  assign new_n43819_ = ~new_n43454_ & ~new_n43818_;
  assign new_n43820_ = \b[28]  & ~new_n43443_;
  assign new_n43821_ = ~new_n43437_ & new_n43820_;
  assign new_n43822_ = ~new_n43445_ & ~new_n43821_;
  assign new_n43823_ = ~new_n43819_ & new_n43822_;
  assign new_n43824_ = ~new_n43445_ & ~new_n43823_;
  assign new_n43825_ = \b[29]  & ~new_n43434_;
  assign new_n43826_ = ~new_n43428_ & new_n43825_;
  assign new_n43827_ = ~new_n43436_ & ~new_n43826_;
  assign new_n43828_ = ~new_n43824_ & new_n43827_;
  assign new_n43829_ = ~new_n43436_ & ~new_n43828_;
  assign new_n43830_ = \b[30]  & ~new_n43425_;
  assign new_n43831_ = ~new_n43419_ & new_n43830_;
  assign new_n43832_ = ~new_n43427_ & ~new_n43831_;
  assign new_n43833_ = ~new_n43829_ & new_n43832_;
  assign new_n43834_ = ~new_n43427_ & ~new_n43833_;
  assign new_n43835_ = \b[31]  & ~new_n43416_;
  assign new_n43836_ = ~new_n43410_ & new_n43835_;
  assign new_n43837_ = ~new_n43418_ & ~new_n43836_;
  assign new_n43838_ = ~new_n43834_ & new_n43837_;
  assign new_n43839_ = ~new_n43418_ & ~new_n43838_;
  assign new_n43840_ = \b[32]  & ~new_n43407_;
  assign new_n43841_ = ~new_n43401_ & new_n43840_;
  assign new_n43842_ = ~new_n43409_ & ~new_n43841_;
  assign new_n43843_ = ~new_n43839_ & new_n43842_;
  assign new_n43844_ = ~new_n43409_ & ~new_n43843_;
  assign new_n43845_ = \b[33]  & ~new_n43398_;
  assign new_n43846_ = ~new_n43392_ & new_n43845_;
  assign new_n43847_ = ~new_n43400_ & ~new_n43846_;
  assign new_n43848_ = ~new_n43844_ & new_n43847_;
  assign new_n43849_ = ~new_n43400_ & ~new_n43848_;
  assign new_n43850_ = \b[34]  & ~new_n43389_;
  assign new_n43851_ = ~new_n43383_ & new_n43850_;
  assign new_n43852_ = ~new_n43391_ & ~new_n43851_;
  assign new_n43853_ = ~new_n43849_ & new_n43852_;
  assign new_n43854_ = ~new_n43391_ & ~new_n43853_;
  assign new_n43855_ = \b[35]  & ~new_n43380_;
  assign new_n43856_ = ~new_n43374_ & new_n43855_;
  assign new_n43857_ = ~new_n43382_ & ~new_n43856_;
  assign new_n43858_ = ~new_n43854_ & new_n43857_;
  assign new_n43859_ = ~new_n43382_ & ~new_n43858_;
  assign new_n43860_ = \b[36]  & ~new_n43371_;
  assign new_n43861_ = ~new_n43365_ & new_n43860_;
  assign new_n43862_ = ~new_n43373_ & ~new_n43861_;
  assign new_n43863_ = ~new_n43859_ & new_n43862_;
  assign new_n43864_ = ~new_n43373_ & ~new_n43863_;
  assign new_n43865_ = \b[37]  & ~new_n43362_;
  assign new_n43866_ = ~new_n43356_ & new_n43865_;
  assign new_n43867_ = ~new_n43364_ & ~new_n43866_;
  assign new_n43868_ = ~new_n43864_ & new_n43867_;
  assign new_n43869_ = ~new_n43364_ & ~new_n43868_;
  assign new_n43870_ = \b[38]  & ~new_n43353_;
  assign new_n43871_ = ~new_n43347_ & new_n43870_;
  assign new_n43872_ = ~new_n43355_ & ~new_n43871_;
  assign new_n43873_ = ~new_n43869_ & new_n43872_;
  assign new_n43874_ = ~new_n43355_ & ~new_n43873_;
  assign new_n43875_ = \b[39]  & ~new_n43344_;
  assign new_n43876_ = ~new_n43338_ & new_n43875_;
  assign new_n43877_ = ~new_n43346_ & ~new_n43876_;
  assign new_n43878_ = ~new_n43874_ & new_n43877_;
  assign new_n43879_ = ~new_n43346_ & ~new_n43878_;
  assign new_n43880_ = \b[40]  & ~new_n43335_;
  assign new_n43881_ = ~new_n43329_ & new_n43880_;
  assign new_n43882_ = ~new_n43337_ & ~new_n43881_;
  assign new_n43883_ = ~new_n43879_ & new_n43882_;
  assign new_n43884_ = ~new_n43337_ & ~new_n43883_;
  assign new_n43885_ = \b[41]  & ~new_n43326_;
  assign new_n43886_ = ~new_n43320_ & new_n43885_;
  assign new_n43887_ = ~new_n43328_ & ~new_n43886_;
  assign new_n43888_ = ~new_n43884_ & new_n43887_;
  assign new_n43889_ = ~new_n43328_ & ~new_n43888_;
  assign new_n43890_ = \b[42]  & ~new_n43317_;
  assign new_n43891_ = ~new_n43311_ & new_n43890_;
  assign new_n43892_ = ~new_n43319_ & ~new_n43891_;
  assign new_n43893_ = ~new_n43889_ & new_n43892_;
  assign new_n43894_ = ~new_n43319_ & ~new_n43893_;
  assign new_n43895_ = \b[43]  & ~new_n43308_;
  assign new_n43896_ = ~new_n43302_ & new_n43895_;
  assign new_n43897_ = ~new_n43310_ & ~new_n43896_;
  assign new_n43898_ = ~new_n43894_ & new_n43897_;
  assign new_n43899_ = ~new_n43310_ & ~new_n43898_;
  assign new_n43900_ = \b[44]  & ~new_n43299_;
  assign new_n43901_ = ~new_n43293_ & new_n43900_;
  assign new_n43902_ = ~new_n43301_ & ~new_n43901_;
  assign new_n43903_ = ~new_n43899_ & new_n43902_;
  assign new_n43904_ = ~new_n43301_ & ~new_n43903_;
  assign new_n43905_ = \b[45]  & ~new_n43290_;
  assign new_n43906_ = ~new_n43284_ & new_n43905_;
  assign new_n43907_ = ~new_n43292_ & ~new_n43906_;
  assign new_n43908_ = ~new_n43904_ & new_n43907_;
  assign new_n43909_ = ~new_n43292_ & ~new_n43908_;
  assign new_n43910_ = ~new_n42672_ & ~new_n43283_;
  assign new_n43911_ = ~new_n42674_ & new_n43280_;
  assign new_n43912_ = ~new_n43276_ & new_n43911_;
  assign new_n43913_ = ~new_n43277_ & ~new_n43280_;
  assign new_n43914_ = ~new_n43912_ & ~new_n43913_;
  assign new_n43915_ = new_n43283_ & ~new_n43914_;
  assign new_n43916_ = ~new_n43910_ & ~new_n43915_;
  assign new_n43917_ = ~\b[46]  & ~new_n43916_;
  assign new_n43918_ = \b[46]  & ~new_n43910_;
  assign new_n43919_ = ~new_n43915_ & new_n43918_;
  assign new_n43920_ = new_n15859_ & ~new_n43919_;
  assign new_n43921_ = ~new_n43917_ & new_n43920_;
  assign new_n43922_ = ~new_n43909_ & new_n43921_;
  assign new_n43923_ = new_n15212_ & ~new_n43916_;
  assign new_n43924_ = ~new_n43922_ & ~new_n43923_;
  assign new_n43925_ = ~new_n43301_ & new_n43907_;
  assign new_n43926_ = ~new_n43903_ & new_n43925_;
  assign new_n43927_ = ~new_n43904_ & ~new_n43907_;
  assign new_n43928_ = ~new_n43926_ & ~new_n43927_;
  assign new_n43929_ = ~new_n43924_ & ~new_n43928_;
  assign new_n43930_ = ~new_n43291_ & ~new_n43923_;
  assign new_n43931_ = ~new_n43922_ & new_n43930_;
  assign new_n43932_ = ~new_n43929_ & ~new_n43931_;
  assign new_n43933_ = ~\b[46]  & ~new_n43932_;
  assign new_n43934_ = ~new_n43310_ & new_n43902_;
  assign new_n43935_ = ~new_n43898_ & new_n43934_;
  assign new_n43936_ = ~new_n43899_ & ~new_n43902_;
  assign new_n43937_ = ~new_n43935_ & ~new_n43936_;
  assign new_n43938_ = ~new_n43924_ & ~new_n43937_;
  assign new_n43939_ = ~new_n43300_ & ~new_n43923_;
  assign new_n43940_ = ~new_n43922_ & new_n43939_;
  assign new_n43941_ = ~new_n43938_ & ~new_n43940_;
  assign new_n43942_ = ~\b[45]  & ~new_n43941_;
  assign new_n43943_ = ~new_n43319_ & new_n43897_;
  assign new_n43944_ = ~new_n43893_ & new_n43943_;
  assign new_n43945_ = ~new_n43894_ & ~new_n43897_;
  assign new_n43946_ = ~new_n43944_ & ~new_n43945_;
  assign new_n43947_ = ~new_n43924_ & ~new_n43946_;
  assign new_n43948_ = ~new_n43309_ & ~new_n43923_;
  assign new_n43949_ = ~new_n43922_ & new_n43948_;
  assign new_n43950_ = ~new_n43947_ & ~new_n43949_;
  assign new_n43951_ = ~\b[44]  & ~new_n43950_;
  assign new_n43952_ = ~new_n43328_ & new_n43892_;
  assign new_n43953_ = ~new_n43888_ & new_n43952_;
  assign new_n43954_ = ~new_n43889_ & ~new_n43892_;
  assign new_n43955_ = ~new_n43953_ & ~new_n43954_;
  assign new_n43956_ = ~new_n43924_ & ~new_n43955_;
  assign new_n43957_ = ~new_n43318_ & ~new_n43923_;
  assign new_n43958_ = ~new_n43922_ & new_n43957_;
  assign new_n43959_ = ~new_n43956_ & ~new_n43958_;
  assign new_n43960_ = ~\b[43]  & ~new_n43959_;
  assign new_n43961_ = ~new_n43337_ & new_n43887_;
  assign new_n43962_ = ~new_n43883_ & new_n43961_;
  assign new_n43963_ = ~new_n43884_ & ~new_n43887_;
  assign new_n43964_ = ~new_n43962_ & ~new_n43963_;
  assign new_n43965_ = ~new_n43924_ & ~new_n43964_;
  assign new_n43966_ = ~new_n43327_ & ~new_n43923_;
  assign new_n43967_ = ~new_n43922_ & new_n43966_;
  assign new_n43968_ = ~new_n43965_ & ~new_n43967_;
  assign new_n43969_ = ~\b[42]  & ~new_n43968_;
  assign new_n43970_ = ~new_n43346_ & new_n43882_;
  assign new_n43971_ = ~new_n43878_ & new_n43970_;
  assign new_n43972_ = ~new_n43879_ & ~new_n43882_;
  assign new_n43973_ = ~new_n43971_ & ~new_n43972_;
  assign new_n43974_ = ~new_n43924_ & ~new_n43973_;
  assign new_n43975_ = ~new_n43336_ & ~new_n43923_;
  assign new_n43976_ = ~new_n43922_ & new_n43975_;
  assign new_n43977_ = ~new_n43974_ & ~new_n43976_;
  assign new_n43978_ = ~\b[41]  & ~new_n43977_;
  assign new_n43979_ = ~new_n43355_ & new_n43877_;
  assign new_n43980_ = ~new_n43873_ & new_n43979_;
  assign new_n43981_ = ~new_n43874_ & ~new_n43877_;
  assign new_n43982_ = ~new_n43980_ & ~new_n43981_;
  assign new_n43983_ = ~new_n43924_ & ~new_n43982_;
  assign new_n43984_ = ~new_n43345_ & ~new_n43923_;
  assign new_n43985_ = ~new_n43922_ & new_n43984_;
  assign new_n43986_ = ~new_n43983_ & ~new_n43985_;
  assign new_n43987_ = ~\b[40]  & ~new_n43986_;
  assign new_n43988_ = ~new_n43364_ & new_n43872_;
  assign new_n43989_ = ~new_n43868_ & new_n43988_;
  assign new_n43990_ = ~new_n43869_ & ~new_n43872_;
  assign new_n43991_ = ~new_n43989_ & ~new_n43990_;
  assign new_n43992_ = ~new_n43924_ & ~new_n43991_;
  assign new_n43993_ = ~new_n43354_ & ~new_n43923_;
  assign new_n43994_ = ~new_n43922_ & new_n43993_;
  assign new_n43995_ = ~new_n43992_ & ~new_n43994_;
  assign new_n43996_ = ~\b[39]  & ~new_n43995_;
  assign new_n43997_ = ~new_n43373_ & new_n43867_;
  assign new_n43998_ = ~new_n43863_ & new_n43997_;
  assign new_n43999_ = ~new_n43864_ & ~new_n43867_;
  assign new_n44000_ = ~new_n43998_ & ~new_n43999_;
  assign new_n44001_ = ~new_n43924_ & ~new_n44000_;
  assign new_n44002_ = ~new_n43363_ & ~new_n43923_;
  assign new_n44003_ = ~new_n43922_ & new_n44002_;
  assign new_n44004_ = ~new_n44001_ & ~new_n44003_;
  assign new_n44005_ = ~\b[38]  & ~new_n44004_;
  assign new_n44006_ = ~new_n43382_ & new_n43862_;
  assign new_n44007_ = ~new_n43858_ & new_n44006_;
  assign new_n44008_ = ~new_n43859_ & ~new_n43862_;
  assign new_n44009_ = ~new_n44007_ & ~new_n44008_;
  assign new_n44010_ = ~new_n43924_ & ~new_n44009_;
  assign new_n44011_ = ~new_n43372_ & ~new_n43923_;
  assign new_n44012_ = ~new_n43922_ & new_n44011_;
  assign new_n44013_ = ~new_n44010_ & ~new_n44012_;
  assign new_n44014_ = ~\b[37]  & ~new_n44013_;
  assign new_n44015_ = ~new_n43391_ & new_n43857_;
  assign new_n44016_ = ~new_n43853_ & new_n44015_;
  assign new_n44017_ = ~new_n43854_ & ~new_n43857_;
  assign new_n44018_ = ~new_n44016_ & ~new_n44017_;
  assign new_n44019_ = ~new_n43924_ & ~new_n44018_;
  assign new_n44020_ = ~new_n43381_ & ~new_n43923_;
  assign new_n44021_ = ~new_n43922_ & new_n44020_;
  assign new_n44022_ = ~new_n44019_ & ~new_n44021_;
  assign new_n44023_ = ~\b[36]  & ~new_n44022_;
  assign new_n44024_ = ~new_n43400_ & new_n43852_;
  assign new_n44025_ = ~new_n43848_ & new_n44024_;
  assign new_n44026_ = ~new_n43849_ & ~new_n43852_;
  assign new_n44027_ = ~new_n44025_ & ~new_n44026_;
  assign new_n44028_ = ~new_n43924_ & ~new_n44027_;
  assign new_n44029_ = ~new_n43390_ & ~new_n43923_;
  assign new_n44030_ = ~new_n43922_ & new_n44029_;
  assign new_n44031_ = ~new_n44028_ & ~new_n44030_;
  assign new_n44032_ = ~\b[35]  & ~new_n44031_;
  assign new_n44033_ = ~new_n43409_ & new_n43847_;
  assign new_n44034_ = ~new_n43843_ & new_n44033_;
  assign new_n44035_ = ~new_n43844_ & ~new_n43847_;
  assign new_n44036_ = ~new_n44034_ & ~new_n44035_;
  assign new_n44037_ = ~new_n43924_ & ~new_n44036_;
  assign new_n44038_ = ~new_n43399_ & ~new_n43923_;
  assign new_n44039_ = ~new_n43922_ & new_n44038_;
  assign new_n44040_ = ~new_n44037_ & ~new_n44039_;
  assign new_n44041_ = ~\b[34]  & ~new_n44040_;
  assign new_n44042_ = ~new_n43418_ & new_n43842_;
  assign new_n44043_ = ~new_n43838_ & new_n44042_;
  assign new_n44044_ = ~new_n43839_ & ~new_n43842_;
  assign new_n44045_ = ~new_n44043_ & ~new_n44044_;
  assign new_n44046_ = ~new_n43924_ & ~new_n44045_;
  assign new_n44047_ = ~new_n43408_ & ~new_n43923_;
  assign new_n44048_ = ~new_n43922_ & new_n44047_;
  assign new_n44049_ = ~new_n44046_ & ~new_n44048_;
  assign new_n44050_ = ~\b[33]  & ~new_n44049_;
  assign new_n44051_ = ~new_n43427_ & new_n43837_;
  assign new_n44052_ = ~new_n43833_ & new_n44051_;
  assign new_n44053_ = ~new_n43834_ & ~new_n43837_;
  assign new_n44054_ = ~new_n44052_ & ~new_n44053_;
  assign new_n44055_ = ~new_n43924_ & ~new_n44054_;
  assign new_n44056_ = ~new_n43417_ & ~new_n43923_;
  assign new_n44057_ = ~new_n43922_ & new_n44056_;
  assign new_n44058_ = ~new_n44055_ & ~new_n44057_;
  assign new_n44059_ = ~\b[32]  & ~new_n44058_;
  assign new_n44060_ = ~new_n43436_ & new_n43832_;
  assign new_n44061_ = ~new_n43828_ & new_n44060_;
  assign new_n44062_ = ~new_n43829_ & ~new_n43832_;
  assign new_n44063_ = ~new_n44061_ & ~new_n44062_;
  assign new_n44064_ = ~new_n43924_ & ~new_n44063_;
  assign new_n44065_ = ~new_n43426_ & ~new_n43923_;
  assign new_n44066_ = ~new_n43922_ & new_n44065_;
  assign new_n44067_ = ~new_n44064_ & ~new_n44066_;
  assign new_n44068_ = ~\b[31]  & ~new_n44067_;
  assign new_n44069_ = ~new_n43445_ & new_n43827_;
  assign new_n44070_ = ~new_n43823_ & new_n44069_;
  assign new_n44071_ = ~new_n43824_ & ~new_n43827_;
  assign new_n44072_ = ~new_n44070_ & ~new_n44071_;
  assign new_n44073_ = ~new_n43924_ & ~new_n44072_;
  assign new_n44074_ = ~new_n43435_ & ~new_n43923_;
  assign new_n44075_ = ~new_n43922_ & new_n44074_;
  assign new_n44076_ = ~new_n44073_ & ~new_n44075_;
  assign new_n44077_ = ~\b[30]  & ~new_n44076_;
  assign new_n44078_ = ~new_n43454_ & new_n43822_;
  assign new_n44079_ = ~new_n43818_ & new_n44078_;
  assign new_n44080_ = ~new_n43819_ & ~new_n43822_;
  assign new_n44081_ = ~new_n44079_ & ~new_n44080_;
  assign new_n44082_ = ~new_n43924_ & ~new_n44081_;
  assign new_n44083_ = ~new_n43444_ & ~new_n43923_;
  assign new_n44084_ = ~new_n43922_ & new_n44083_;
  assign new_n44085_ = ~new_n44082_ & ~new_n44084_;
  assign new_n44086_ = ~\b[29]  & ~new_n44085_;
  assign new_n44087_ = ~new_n43463_ & new_n43817_;
  assign new_n44088_ = ~new_n43813_ & new_n44087_;
  assign new_n44089_ = ~new_n43814_ & ~new_n43817_;
  assign new_n44090_ = ~new_n44088_ & ~new_n44089_;
  assign new_n44091_ = ~new_n43924_ & ~new_n44090_;
  assign new_n44092_ = ~new_n43453_ & ~new_n43923_;
  assign new_n44093_ = ~new_n43922_ & new_n44092_;
  assign new_n44094_ = ~new_n44091_ & ~new_n44093_;
  assign new_n44095_ = ~\b[28]  & ~new_n44094_;
  assign new_n44096_ = ~new_n43472_ & new_n43812_;
  assign new_n44097_ = ~new_n43808_ & new_n44096_;
  assign new_n44098_ = ~new_n43809_ & ~new_n43812_;
  assign new_n44099_ = ~new_n44097_ & ~new_n44098_;
  assign new_n44100_ = ~new_n43924_ & ~new_n44099_;
  assign new_n44101_ = ~new_n43462_ & ~new_n43923_;
  assign new_n44102_ = ~new_n43922_ & new_n44101_;
  assign new_n44103_ = ~new_n44100_ & ~new_n44102_;
  assign new_n44104_ = ~\b[27]  & ~new_n44103_;
  assign new_n44105_ = ~new_n43481_ & new_n43807_;
  assign new_n44106_ = ~new_n43803_ & new_n44105_;
  assign new_n44107_ = ~new_n43804_ & ~new_n43807_;
  assign new_n44108_ = ~new_n44106_ & ~new_n44107_;
  assign new_n44109_ = ~new_n43924_ & ~new_n44108_;
  assign new_n44110_ = ~new_n43471_ & ~new_n43923_;
  assign new_n44111_ = ~new_n43922_ & new_n44110_;
  assign new_n44112_ = ~new_n44109_ & ~new_n44111_;
  assign new_n44113_ = ~\b[26]  & ~new_n44112_;
  assign new_n44114_ = ~new_n43490_ & new_n43802_;
  assign new_n44115_ = ~new_n43798_ & new_n44114_;
  assign new_n44116_ = ~new_n43799_ & ~new_n43802_;
  assign new_n44117_ = ~new_n44115_ & ~new_n44116_;
  assign new_n44118_ = ~new_n43924_ & ~new_n44117_;
  assign new_n44119_ = ~new_n43480_ & ~new_n43923_;
  assign new_n44120_ = ~new_n43922_ & new_n44119_;
  assign new_n44121_ = ~new_n44118_ & ~new_n44120_;
  assign new_n44122_ = ~\b[25]  & ~new_n44121_;
  assign new_n44123_ = ~new_n43499_ & new_n43797_;
  assign new_n44124_ = ~new_n43793_ & new_n44123_;
  assign new_n44125_ = ~new_n43794_ & ~new_n43797_;
  assign new_n44126_ = ~new_n44124_ & ~new_n44125_;
  assign new_n44127_ = ~new_n43924_ & ~new_n44126_;
  assign new_n44128_ = ~new_n43489_ & ~new_n43923_;
  assign new_n44129_ = ~new_n43922_ & new_n44128_;
  assign new_n44130_ = ~new_n44127_ & ~new_n44129_;
  assign new_n44131_ = ~\b[24]  & ~new_n44130_;
  assign new_n44132_ = ~new_n43508_ & new_n43792_;
  assign new_n44133_ = ~new_n43788_ & new_n44132_;
  assign new_n44134_ = ~new_n43789_ & ~new_n43792_;
  assign new_n44135_ = ~new_n44133_ & ~new_n44134_;
  assign new_n44136_ = ~new_n43924_ & ~new_n44135_;
  assign new_n44137_ = ~new_n43498_ & ~new_n43923_;
  assign new_n44138_ = ~new_n43922_ & new_n44137_;
  assign new_n44139_ = ~new_n44136_ & ~new_n44138_;
  assign new_n44140_ = ~\b[23]  & ~new_n44139_;
  assign new_n44141_ = ~new_n43517_ & new_n43787_;
  assign new_n44142_ = ~new_n43783_ & new_n44141_;
  assign new_n44143_ = ~new_n43784_ & ~new_n43787_;
  assign new_n44144_ = ~new_n44142_ & ~new_n44143_;
  assign new_n44145_ = ~new_n43924_ & ~new_n44144_;
  assign new_n44146_ = ~new_n43507_ & ~new_n43923_;
  assign new_n44147_ = ~new_n43922_ & new_n44146_;
  assign new_n44148_ = ~new_n44145_ & ~new_n44147_;
  assign new_n44149_ = ~\b[22]  & ~new_n44148_;
  assign new_n44150_ = ~new_n43526_ & new_n43782_;
  assign new_n44151_ = ~new_n43778_ & new_n44150_;
  assign new_n44152_ = ~new_n43779_ & ~new_n43782_;
  assign new_n44153_ = ~new_n44151_ & ~new_n44152_;
  assign new_n44154_ = ~new_n43924_ & ~new_n44153_;
  assign new_n44155_ = ~new_n43516_ & ~new_n43923_;
  assign new_n44156_ = ~new_n43922_ & new_n44155_;
  assign new_n44157_ = ~new_n44154_ & ~new_n44156_;
  assign new_n44158_ = ~\b[21]  & ~new_n44157_;
  assign new_n44159_ = ~new_n43535_ & new_n43777_;
  assign new_n44160_ = ~new_n43773_ & new_n44159_;
  assign new_n44161_ = ~new_n43774_ & ~new_n43777_;
  assign new_n44162_ = ~new_n44160_ & ~new_n44161_;
  assign new_n44163_ = ~new_n43924_ & ~new_n44162_;
  assign new_n44164_ = ~new_n43525_ & ~new_n43923_;
  assign new_n44165_ = ~new_n43922_ & new_n44164_;
  assign new_n44166_ = ~new_n44163_ & ~new_n44165_;
  assign new_n44167_ = ~\b[20]  & ~new_n44166_;
  assign new_n44168_ = ~new_n43544_ & new_n43772_;
  assign new_n44169_ = ~new_n43768_ & new_n44168_;
  assign new_n44170_ = ~new_n43769_ & ~new_n43772_;
  assign new_n44171_ = ~new_n44169_ & ~new_n44170_;
  assign new_n44172_ = ~new_n43924_ & ~new_n44171_;
  assign new_n44173_ = ~new_n43534_ & ~new_n43923_;
  assign new_n44174_ = ~new_n43922_ & new_n44173_;
  assign new_n44175_ = ~new_n44172_ & ~new_n44174_;
  assign new_n44176_ = ~\b[19]  & ~new_n44175_;
  assign new_n44177_ = ~new_n43553_ & new_n43767_;
  assign new_n44178_ = ~new_n43763_ & new_n44177_;
  assign new_n44179_ = ~new_n43764_ & ~new_n43767_;
  assign new_n44180_ = ~new_n44178_ & ~new_n44179_;
  assign new_n44181_ = ~new_n43924_ & ~new_n44180_;
  assign new_n44182_ = ~new_n43543_ & ~new_n43923_;
  assign new_n44183_ = ~new_n43922_ & new_n44182_;
  assign new_n44184_ = ~new_n44181_ & ~new_n44183_;
  assign new_n44185_ = ~\b[18]  & ~new_n44184_;
  assign new_n44186_ = ~new_n43562_ & new_n43762_;
  assign new_n44187_ = ~new_n43758_ & new_n44186_;
  assign new_n44188_ = ~new_n43759_ & ~new_n43762_;
  assign new_n44189_ = ~new_n44187_ & ~new_n44188_;
  assign new_n44190_ = ~new_n43924_ & ~new_n44189_;
  assign new_n44191_ = ~new_n43552_ & ~new_n43923_;
  assign new_n44192_ = ~new_n43922_ & new_n44191_;
  assign new_n44193_ = ~new_n44190_ & ~new_n44192_;
  assign new_n44194_ = ~\b[17]  & ~new_n44193_;
  assign new_n44195_ = ~new_n43571_ & new_n43757_;
  assign new_n44196_ = ~new_n43753_ & new_n44195_;
  assign new_n44197_ = ~new_n43754_ & ~new_n43757_;
  assign new_n44198_ = ~new_n44196_ & ~new_n44197_;
  assign new_n44199_ = ~new_n43924_ & ~new_n44198_;
  assign new_n44200_ = ~new_n43561_ & ~new_n43923_;
  assign new_n44201_ = ~new_n43922_ & new_n44200_;
  assign new_n44202_ = ~new_n44199_ & ~new_n44201_;
  assign new_n44203_ = ~\b[16]  & ~new_n44202_;
  assign new_n44204_ = ~new_n43580_ & new_n43752_;
  assign new_n44205_ = ~new_n43748_ & new_n44204_;
  assign new_n44206_ = ~new_n43749_ & ~new_n43752_;
  assign new_n44207_ = ~new_n44205_ & ~new_n44206_;
  assign new_n44208_ = ~new_n43924_ & ~new_n44207_;
  assign new_n44209_ = ~new_n43570_ & ~new_n43923_;
  assign new_n44210_ = ~new_n43922_ & new_n44209_;
  assign new_n44211_ = ~new_n44208_ & ~new_n44210_;
  assign new_n44212_ = ~\b[15]  & ~new_n44211_;
  assign new_n44213_ = ~new_n43589_ & new_n43747_;
  assign new_n44214_ = ~new_n43743_ & new_n44213_;
  assign new_n44215_ = ~new_n43744_ & ~new_n43747_;
  assign new_n44216_ = ~new_n44214_ & ~new_n44215_;
  assign new_n44217_ = ~new_n43924_ & ~new_n44216_;
  assign new_n44218_ = ~new_n43579_ & ~new_n43923_;
  assign new_n44219_ = ~new_n43922_ & new_n44218_;
  assign new_n44220_ = ~new_n44217_ & ~new_n44219_;
  assign new_n44221_ = ~\b[14]  & ~new_n44220_;
  assign new_n44222_ = ~new_n43598_ & new_n43742_;
  assign new_n44223_ = ~new_n43738_ & new_n44222_;
  assign new_n44224_ = ~new_n43739_ & ~new_n43742_;
  assign new_n44225_ = ~new_n44223_ & ~new_n44224_;
  assign new_n44226_ = ~new_n43924_ & ~new_n44225_;
  assign new_n44227_ = ~new_n43588_ & ~new_n43923_;
  assign new_n44228_ = ~new_n43922_ & new_n44227_;
  assign new_n44229_ = ~new_n44226_ & ~new_n44228_;
  assign new_n44230_ = ~\b[13]  & ~new_n44229_;
  assign new_n44231_ = ~new_n43607_ & new_n43737_;
  assign new_n44232_ = ~new_n43733_ & new_n44231_;
  assign new_n44233_ = ~new_n43734_ & ~new_n43737_;
  assign new_n44234_ = ~new_n44232_ & ~new_n44233_;
  assign new_n44235_ = ~new_n43924_ & ~new_n44234_;
  assign new_n44236_ = ~new_n43597_ & ~new_n43923_;
  assign new_n44237_ = ~new_n43922_ & new_n44236_;
  assign new_n44238_ = ~new_n44235_ & ~new_n44237_;
  assign new_n44239_ = ~\b[12]  & ~new_n44238_;
  assign new_n44240_ = ~new_n43616_ & new_n43732_;
  assign new_n44241_ = ~new_n43728_ & new_n44240_;
  assign new_n44242_ = ~new_n43729_ & ~new_n43732_;
  assign new_n44243_ = ~new_n44241_ & ~new_n44242_;
  assign new_n44244_ = ~new_n43924_ & ~new_n44243_;
  assign new_n44245_ = ~new_n43606_ & ~new_n43923_;
  assign new_n44246_ = ~new_n43922_ & new_n44245_;
  assign new_n44247_ = ~new_n44244_ & ~new_n44246_;
  assign new_n44248_ = ~\b[11]  & ~new_n44247_;
  assign new_n44249_ = ~new_n43625_ & new_n43727_;
  assign new_n44250_ = ~new_n43723_ & new_n44249_;
  assign new_n44251_ = ~new_n43724_ & ~new_n43727_;
  assign new_n44252_ = ~new_n44250_ & ~new_n44251_;
  assign new_n44253_ = ~new_n43924_ & ~new_n44252_;
  assign new_n44254_ = ~new_n43615_ & ~new_n43923_;
  assign new_n44255_ = ~new_n43922_ & new_n44254_;
  assign new_n44256_ = ~new_n44253_ & ~new_n44255_;
  assign new_n44257_ = ~\b[10]  & ~new_n44256_;
  assign new_n44258_ = ~new_n43634_ & new_n43722_;
  assign new_n44259_ = ~new_n43718_ & new_n44258_;
  assign new_n44260_ = ~new_n43719_ & ~new_n43722_;
  assign new_n44261_ = ~new_n44259_ & ~new_n44260_;
  assign new_n44262_ = ~new_n43924_ & ~new_n44261_;
  assign new_n44263_ = ~new_n43624_ & ~new_n43923_;
  assign new_n44264_ = ~new_n43922_ & new_n44263_;
  assign new_n44265_ = ~new_n44262_ & ~new_n44264_;
  assign new_n44266_ = ~\b[9]  & ~new_n44265_;
  assign new_n44267_ = ~new_n43643_ & new_n43717_;
  assign new_n44268_ = ~new_n43713_ & new_n44267_;
  assign new_n44269_ = ~new_n43714_ & ~new_n43717_;
  assign new_n44270_ = ~new_n44268_ & ~new_n44269_;
  assign new_n44271_ = ~new_n43924_ & ~new_n44270_;
  assign new_n44272_ = ~new_n43633_ & ~new_n43923_;
  assign new_n44273_ = ~new_n43922_ & new_n44272_;
  assign new_n44274_ = ~new_n44271_ & ~new_n44273_;
  assign new_n44275_ = ~\b[8]  & ~new_n44274_;
  assign new_n44276_ = ~new_n43652_ & new_n43712_;
  assign new_n44277_ = ~new_n43708_ & new_n44276_;
  assign new_n44278_ = ~new_n43709_ & ~new_n43712_;
  assign new_n44279_ = ~new_n44277_ & ~new_n44278_;
  assign new_n44280_ = ~new_n43924_ & ~new_n44279_;
  assign new_n44281_ = ~new_n43642_ & ~new_n43923_;
  assign new_n44282_ = ~new_n43922_ & new_n44281_;
  assign new_n44283_ = ~new_n44280_ & ~new_n44282_;
  assign new_n44284_ = ~\b[7]  & ~new_n44283_;
  assign new_n44285_ = ~new_n43661_ & new_n43707_;
  assign new_n44286_ = ~new_n43703_ & new_n44285_;
  assign new_n44287_ = ~new_n43704_ & ~new_n43707_;
  assign new_n44288_ = ~new_n44286_ & ~new_n44287_;
  assign new_n44289_ = ~new_n43924_ & ~new_n44288_;
  assign new_n44290_ = ~new_n43651_ & ~new_n43923_;
  assign new_n44291_ = ~new_n43922_ & new_n44290_;
  assign new_n44292_ = ~new_n44289_ & ~new_n44291_;
  assign new_n44293_ = ~\b[6]  & ~new_n44292_;
  assign new_n44294_ = ~new_n43670_ & new_n43702_;
  assign new_n44295_ = ~new_n43698_ & new_n44294_;
  assign new_n44296_ = ~new_n43699_ & ~new_n43702_;
  assign new_n44297_ = ~new_n44295_ & ~new_n44296_;
  assign new_n44298_ = ~new_n43924_ & ~new_n44297_;
  assign new_n44299_ = ~new_n43660_ & ~new_n43923_;
  assign new_n44300_ = ~new_n43922_ & new_n44299_;
  assign new_n44301_ = ~new_n44298_ & ~new_n44300_;
  assign new_n44302_ = ~\b[5]  & ~new_n44301_;
  assign new_n44303_ = ~new_n43678_ & new_n43697_;
  assign new_n44304_ = ~new_n43693_ & new_n44303_;
  assign new_n44305_ = ~new_n43694_ & ~new_n43697_;
  assign new_n44306_ = ~new_n44304_ & ~new_n44305_;
  assign new_n44307_ = ~new_n43924_ & ~new_n44306_;
  assign new_n44308_ = ~new_n43669_ & ~new_n43923_;
  assign new_n44309_ = ~new_n43922_ & new_n44308_;
  assign new_n44310_ = ~new_n44307_ & ~new_n44309_;
  assign new_n44311_ = ~\b[4]  & ~new_n44310_;
  assign new_n44312_ = ~new_n43688_ & new_n43692_;
  assign new_n44313_ = ~new_n43687_ & new_n44312_;
  assign new_n44314_ = ~new_n43689_ & ~new_n43692_;
  assign new_n44315_ = ~new_n44313_ & ~new_n44314_;
  assign new_n44316_ = ~new_n43924_ & ~new_n44315_;
  assign new_n44317_ = ~new_n43677_ & ~new_n43923_;
  assign new_n44318_ = ~new_n43922_ & new_n44317_;
  assign new_n44319_ = ~new_n44316_ & ~new_n44318_;
  assign new_n44320_ = ~\b[3]  & ~new_n44319_;
  assign new_n44321_ = new_n15624_ & ~new_n43685_;
  assign new_n44322_ = ~new_n43683_ & new_n44321_;
  assign new_n44323_ = ~new_n43687_ & ~new_n44322_;
  assign new_n44324_ = ~new_n43924_ & new_n44323_;
  assign new_n44325_ = ~new_n43682_ & ~new_n43923_;
  assign new_n44326_ = ~new_n43922_ & new_n44325_;
  assign new_n44327_ = ~new_n44324_ & ~new_n44326_;
  assign new_n44328_ = ~\b[2]  & ~new_n44327_;
  assign new_n44329_ = \b[0]  & ~new_n43924_;
  assign new_n44330_ = \a[17]  & ~new_n44329_;
  assign new_n44331_ = new_n15624_ & ~new_n43924_;
  assign new_n44332_ = ~new_n44330_ & ~new_n44331_;
  assign new_n44333_ = \b[1]  & ~new_n44332_;
  assign new_n44334_ = ~\b[1]  & ~new_n44331_;
  assign new_n44335_ = ~new_n44330_ & new_n44334_;
  assign new_n44336_ = ~new_n44333_ & ~new_n44335_;
  assign new_n44337_ = ~new_n16277_ & ~new_n44336_;
  assign new_n44338_ = ~\b[1]  & ~new_n44332_;
  assign new_n44339_ = ~new_n44337_ & ~new_n44338_;
  assign new_n44340_ = \b[2]  & ~new_n44326_;
  assign new_n44341_ = ~new_n44324_ & new_n44340_;
  assign new_n44342_ = ~new_n44328_ & ~new_n44341_;
  assign new_n44343_ = ~new_n44339_ & new_n44342_;
  assign new_n44344_ = ~new_n44328_ & ~new_n44343_;
  assign new_n44345_ = \b[3]  & ~new_n44318_;
  assign new_n44346_ = ~new_n44316_ & new_n44345_;
  assign new_n44347_ = ~new_n44320_ & ~new_n44346_;
  assign new_n44348_ = ~new_n44344_ & new_n44347_;
  assign new_n44349_ = ~new_n44320_ & ~new_n44348_;
  assign new_n44350_ = \b[4]  & ~new_n44309_;
  assign new_n44351_ = ~new_n44307_ & new_n44350_;
  assign new_n44352_ = ~new_n44311_ & ~new_n44351_;
  assign new_n44353_ = ~new_n44349_ & new_n44352_;
  assign new_n44354_ = ~new_n44311_ & ~new_n44353_;
  assign new_n44355_ = \b[5]  & ~new_n44300_;
  assign new_n44356_ = ~new_n44298_ & new_n44355_;
  assign new_n44357_ = ~new_n44302_ & ~new_n44356_;
  assign new_n44358_ = ~new_n44354_ & new_n44357_;
  assign new_n44359_ = ~new_n44302_ & ~new_n44358_;
  assign new_n44360_ = \b[6]  & ~new_n44291_;
  assign new_n44361_ = ~new_n44289_ & new_n44360_;
  assign new_n44362_ = ~new_n44293_ & ~new_n44361_;
  assign new_n44363_ = ~new_n44359_ & new_n44362_;
  assign new_n44364_ = ~new_n44293_ & ~new_n44363_;
  assign new_n44365_ = \b[7]  & ~new_n44282_;
  assign new_n44366_ = ~new_n44280_ & new_n44365_;
  assign new_n44367_ = ~new_n44284_ & ~new_n44366_;
  assign new_n44368_ = ~new_n44364_ & new_n44367_;
  assign new_n44369_ = ~new_n44284_ & ~new_n44368_;
  assign new_n44370_ = \b[8]  & ~new_n44273_;
  assign new_n44371_ = ~new_n44271_ & new_n44370_;
  assign new_n44372_ = ~new_n44275_ & ~new_n44371_;
  assign new_n44373_ = ~new_n44369_ & new_n44372_;
  assign new_n44374_ = ~new_n44275_ & ~new_n44373_;
  assign new_n44375_ = \b[9]  & ~new_n44264_;
  assign new_n44376_ = ~new_n44262_ & new_n44375_;
  assign new_n44377_ = ~new_n44266_ & ~new_n44376_;
  assign new_n44378_ = ~new_n44374_ & new_n44377_;
  assign new_n44379_ = ~new_n44266_ & ~new_n44378_;
  assign new_n44380_ = \b[10]  & ~new_n44255_;
  assign new_n44381_ = ~new_n44253_ & new_n44380_;
  assign new_n44382_ = ~new_n44257_ & ~new_n44381_;
  assign new_n44383_ = ~new_n44379_ & new_n44382_;
  assign new_n44384_ = ~new_n44257_ & ~new_n44383_;
  assign new_n44385_ = \b[11]  & ~new_n44246_;
  assign new_n44386_ = ~new_n44244_ & new_n44385_;
  assign new_n44387_ = ~new_n44248_ & ~new_n44386_;
  assign new_n44388_ = ~new_n44384_ & new_n44387_;
  assign new_n44389_ = ~new_n44248_ & ~new_n44388_;
  assign new_n44390_ = \b[12]  & ~new_n44237_;
  assign new_n44391_ = ~new_n44235_ & new_n44390_;
  assign new_n44392_ = ~new_n44239_ & ~new_n44391_;
  assign new_n44393_ = ~new_n44389_ & new_n44392_;
  assign new_n44394_ = ~new_n44239_ & ~new_n44393_;
  assign new_n44395_ = \b[13]  & ~new_n44228_;
  assign new_n44396_ = ~new_n44226_ & new_n44395_;
  assign new_n44397_ = ~new_n44230_ & ~new_n44396_;
  assign new_n44398_ = ~new_n44394_ & new_n44397_;
  assign new_n44399_ = ~new_n44230_ & ~new_n44398_;
  assign new_n44400_ = \b[14]  & ~new_n44219_;
  assign new_n44401_ = ~new_n44217_ & new_n44400_;
  assign new_n44402_ = ~new_n44221_ & ~new_n44401_;
  assign new_n44403_ = ~new_n44399_ & new_n44402_;
  assign new_n44404_ = ~new_n44221_ & ~new_n44403_;
  assign new_n44405_ = \b[15]  & ~new_n44210_;
  assign new_n44406_ = ~new_n44208_ & new_n44405_;
  assign new_n44407_ = ~new_n44212_ & ~new_n44406_;
  assign new_n44408_ = ~new_n44404_ & new_n44407_;
  assign new_n44409_ = ~new_n44212_ & ~new_n44408_;
  assign new_n44410_ = \b[16]  & ~new_n44201_;
  assign new_n44411_ = ~new_n44199_ & new_n44410_;
  assign new_n44412_ = ~new_n44203_ & ~new_n44411_;
  assign new_n44413_ = ~new_n44409_ & new_n44412_;
  assign new_n44414_ = ~new_n44203_ & ~new_n44413_;
  assign new_n44415_ = \b[17]  & ~new_n44192_;
  assign new_n44416_ = ~new_n44190_ & new_n44415_;
  assign new_n44417_ = ~new_n44194_ & ~new_n44416_;
  assign new_n44418_ = ~new_n44414_ & new_n44417_;
  assign new_n44419_ = ~new_n44194_ & ~new_n44418_;
  assign new_n44420_ = \b[18]  & ~new_n44183_;
  assign new_n44421_ = ~new_n44181_ & new_n44420_;
  assign new_n44422_ = ~new_n44185_ & ~new_n44421_;
  assign new_n44423_ = ~new_n44419_ & new_n44422_;
  assign new_n44424_ = ~new_n44185_ & ~new_n44423_;
  assign new_n44425_ = \b[19]  & ~new_n44174_;
  assign new_n44426_ = ~new_n44172_ & new_n44425_;
  assign new_n44427_ = ~new_n44176_ & ~new_n44426_;
  assign new_n44428_ = ~new_n44424_ & new_n44427_;
  assign new_n44429_ = ~new_n44176_ & ~new_n44428_;
  assign new_n44430_ = \b[20]  & ~new_n44165_;
  assign new_n44431_ = ~new_n44163_ & new_n44430_;
  assign new_n44432_ = ~new_n44167_ & ~new_n44431_;
  assign new_n44433_ = ~new_n44429_ & new_n44432_;
  assign new_n44434_ = ~new_n44167_ & ~new_n44433_;
  assign new_n44435_ = \b[21]  & ~new_n44156_;
  assign new_n44436_ = ~new_n44154_ & new_n44435_;
  assign new_n44437_ = ~new_n44158_ & ~new_n44436_;
  assign new_n44438_ = ~new_n44434_ & new_n44437_;
  assign new_n44439_ = ~new_n44158_ & ~new_n44438_;
  assign new_n44440_ = \b[22]  & ~new_n44147_;
  assign new_n44441_ = ~new_n44145_ & new_n44440_;
  assign new_n44442_ = ~new_n44149_ & ~new_n44441_;
  assign new_n44443_ = ~new_n44439_ & new_n44442_;
  assign new_n44444_ = ~new_n44149_ & ~new_n44443_;
  assign new_n44445_ = \b[23]  & ~new_n44138_;
  assign new_n44446_ = ~new_n44136_ & new_n44445_;
  assign new_n44447_ = ~new_n44140_ & ~new_n44446_;
  assign new_n44448_ = ~new_n44444_ & new_n44447_;
  assign new_n44449_ = ~new_n44140_ & ~new_n44448_;
  assign new_n44450_ = \b[24]  & ~new_n44129_;
  assign new_n44451_ = ~new_n44127_ & new_n44450_;
  assign new_n44452_ = ~new_n44131_ & ~new_n44451_;
  assign new_n44453_ = ~new_n44449_ & new_n44452_;
  assign new_n44454_ = ~new_n44131_ & ~new_n44453_;
  assign new_n44455_ = \b[25]  & ~new_n44120_;
  assign new_n44456_ = ~new_n44118_ & new_n44455_;
  assign new_n44457_ = ~new_n44122_ & ~new_n44456_;
  assign new_n44458_ = ~new_n44454_ & new_n44457_;
  assign new_n44459_ = ~new_n44122_ & ~new_n44458_;
  assign new_n44460_ = \b[26]  & ~new_n44111_;
  assign new_n44461_ = ~new_n44109_ & new_n44460_;
  assign new_n44462_ = ~new_n44113_ & ~new_n44461_;
  assign new_n44463_ = ~new_n44459_ & new_n44462_;
  assign new_n44464_ = ~new_n44113_ & ~new_n44463_;
  assign new_n44465_ = \b[27]  & ~new_n44102_;
  assign new_n44466_ = ~new_n44100_ & new_n44465_;
  assign new_n44467_ = ~new_n44104_ & ~new_n44466_;
  assign new_n44468_ = ~new_n44464_ & new_n44467_;
  assign new_n44469_ = ~new_n44104_ & ~new_n44468_;
  assign new_n44470_ = \b[28]  & ~new_n44093_;
  assign new_n44471_ = ~new_n44091_ & new_n44470_;
  assign new_n44472_ = ~new_n44095_ & ~new_n44471_;
  assign new_n44473_ = ~new_n44469_ & new_n44472_;
  assign new_n44474_ = ~new_n44095_ & ~new_n44473_;
  assign new_n44475_ = \b[29]  & ~new_n44084_;
  assign new_n44476_ = ~new_n44082_ & new_n44475_;
  assign new_n44477_ = ~new_n44086_ & ~new_n44476_;
  assign new_n44478_ = ~new_n44474_ & new_n44477_;
  assign new_n44479_ = ~new_n44086_ & ~new_n44478_;
  assign new_n44480_ = \b[30]  & ~new_n44075_;
  assign new_n44481_ = ~new_n44073_ & new_n44480_;
  assign new_n44482_ = ~new_n44077_ & ~new_n44481_;
  assign new_n44483_ = ~new_n44479_ & new_n44482_;
  assign new_n44484_ = ~new_n44077_ & ~new_n44483_;
  assign new_n44485_ = \b[31]  & ~new_n44066_;
  assign new_n44486_ = ~new_n44064_ & new_n44485_;
  assign new_n44487_ = ~new_n44068_ & ~new_n44486_;
  assign new_n44488_ = ~new_n44484_ & new_n44487_;
  assign new_n44489_ = ~new_n44068_ & ~new_n44488_;
  assign new_n44490_ = \b[32]  & ~new_n44057_;
  assign new_n44491_ = ~new_n44055_ & new_n44490_;
  assign new_n44492_ = ~new_n44059_ & ~new_n44491_;
  assign new_n44493_ = ~new_n44489_ & new_n44492_;
  assign new_n44494_ = ~new_n44059_ & ~new_n44493_;
  assign new_n44495_ = \b[33]  & ~new_n44048_;
  assign new_n44496_ = ~new_n44046_ & new_n44495_;
  assign new_n44497_ = ~new_n44050_ & ~new_n44496_;
  assign new_n44498_ = ~new_n44494_ & new_n44497_;
  assign new_n44499_ = ~new_n44050_ & ~new_n44498_;
  assign new_n44500_ = \b[34]  & ~new_n44039_;
  assign new_n44501_ = ~new_n44037_ & new_n44500_;
  assign new_n44502_ = ~new_n44041_ & ~new_n44501_;
  assign new_n44503_ = ~new_n44499_ & new_n44502_;
  assign new_n44504_ = ~new_n44041_ & ~new_n44503_;
  assign new_n44505_ = \b[35]  & ~new_n44030_;
  assign new_n44506_ = ~new_n44028_ & new_n44505_;
  assign new_n44507_ = ~new_n44032_ & ~new_n44506_;
  assign new_n44508_ = ~new_n44504_ & new_n44507_;
  assign new_n44509_ = ~new_n44032_ & ~new_n44508_;
  assign new_n44510_ = \b[36]  & ~new_n44021_;
  assign new_n44511_ = ~new_n44019_ & new_n44510_;
  assign new_n44512_ = ~new_n44023_ & ~new_n44511_;
  assign new_n44513_ = ~new_n44509_ & new_n44512_;
  assign new_n44514_ = ~new_n44023_ & ~new_n44513_;
  assign new_n44515_ = \b[37]  & ~new_n44012_;
  assign new_n44516_ = ~new_n44010_ & new_n44515_;
  assign new_n44517_ = ~new_n44014_ & ~new_n44516_;
  assign new_n44518_ = ~new_n44514_ & new_n44517_;
  assign new_n44519_ = ~new_n44014_ & ~new_n44518_;
  assign new_n44520_ = \b[38]  & ~new_n44003_;
  assign new_n44521_ = ~new_n44001_ & new_n44520_;
  assign new_n44522_ = ~new_n44005_ & ~new_n44521_;
  assign new_n44523_ = ~new_n44519_ & new_n44522_;
  assign new_n44524_ = ~new_n44005_ & ~new_n44523_;
  assign new_n44525_ = \b[39]  & ~new_n43994_;
  assign new_n44526_ = ~new_n43992_ & new_n44525_;
  assign new_n44527_ = ~new_n43996_ & ~new_n44526_;
  assign new_n44528_ = ~new_n44524_ & new_n44527_;
  assign new_n44529_ = ~new_n43996_ & ~new_n44528_;
  assign new_n44530_ = \b[40]  & ~new_n43985_;
  assign new_n44531_ = ~new_n43983_ & new_n44530_;
  assign new_n44532_ = ~new_n43987_ & ~new_n44531_;
  assign new_n44533_ = ~new_n44529_ & new_n44532_;
  assign new_n44534_ = ~new_n43987_ & ~new_n44533_;
  assign new_n44535_ = \b[41]  & ~new_n43976_;
  assign new_n44536_ = ~new_n43974_ & new_n44535_;
  assign new_n44537_ = ~new_n43978_ & ~new_n44536_;
  assign new_n44538_ = ~new_n44534_ & new_n44537_;
  assign new_n44539_ = ~new_n43978_ & ~new_n44538_;
  assign new_n44540_ = \b[42]  & ~new_n43967_;
  assign new_n44541_ = ~new_n43965_ & new_n44540_;
  assign new_n44542_ = ~new_n43969_ & ~new_n44541_;
  assign new_n44543_ = ~new_n44539_ & new_n44542_;
  assign new_n44544_ = ~new_n43969_ & ~new_n44543_;
  assign new_n44545_ = \b[43]  & ~new_n43958_;
  assign new_n44546_ = ~new_n43956_ & new_n44545_;
  assign new_n44547_ = ~new_n43960_ & ~new_n44546_;
  assign new_n44548_ = ~new_n44544_ & new_n44547_;
  assign new_n44549_ = ~new_n43960_ & ~new_n44548_;
  assign new_n44550_ = \b[44]  & ~new_n43949_;
  assign new_n44551_ = ~new_n43947_ & new_n44550_;
  assign new_n44552_ = ~new_n43951_ & ~new_n44551_;
  assign new_n44553_ = ~new_n44549_ & new_n44552_;
  assign new_n44554_ = ~new_n43951_ & ~new_n44553_;
  assign new_n44555_ = \b[45]  & ~new_n43940_;
  assign new_n44556_ = ~new_n43938_ & new_n44555_;
  assign new_n44557_ = ~new_n43942_ & ~new_n44556_;
  assign new_n44558_ = ~new_n44554_ & new_n44557_;
  assign new_n44559_ = ~new_n43942_ & ~new_n44558_;
  assign new_n44560_ = \b[46]  & ~new_n43931_;
  assign new_n44561_ = ~new_n43929_ & new_n44560_;
  assign new_n44562_ = ~new_n43933_ & ~new_n44561_;
  assign new_n44563_ = ~new_n44559_ & new_n44562_;
  assign new_n44564_ = ~new_n43933_ & ~new_n44563_;
  assign new_n44565_ = ~new_n43292_ & ~new_n43919_;
  assign new_n44566_ = ~new_n43917_ & new_n44565_;
  assign new_n44567_ = ~new_n43908_ & new_n44566_;
  assign new_n44568_ = ~new_n43917_ & ~new_n43919_;
  assign new_n44569_ = ~new_n43909_ & ~new_n44568_;
  assign new_n44570_ = ~new_n44567_ & ~new_n44569_;
  assign new_n44571_ = ~new_n43924_ & ~new_n44570_;
  assign new_n44572_ = ~new_n43916_ & ~new_n43923_;
  assign new_n44573_ = ~new_n43922_ & new_n44572_;
  assign new_n44574_ = ~new_n44571_ & ~new_n44573_;
  assign new_n44575_ = ~\b[47]  & ~new_n44574_;
  assign new_n44576_ = \b[47]  & ~new_n44573_;
  assign new_n44577_ = ~new_n44571_ & new_n44576_;
  assign new_n44578_ = new_n338_ & ~new_n44577_;
  assign new_n44579_ = ~new_n44575_ & new_n44578_;
  assign new_n44580_ = ~new_n44564_ & new_n44579_;
  assign new_n44581_ = new_n15859_ & ~new_n44574_;
  assign new_n44582_ = ~new_n44580_ & ~new_n44581_;
  assign new_n44583_ = ~new_n43942_ & new_n44562_;
  assign new_n44584_ = ~new_n44558_ & new_n44583_;
  assign new_n44585_ = ~new_n44559_ & ~new_n44562_;
  assign new_n44586_ = ~new_n44584_ & ~new_n44585_;
  assign new_n44587_ = ~new_n44582_ & ~new_n44586_;
  assign new_n44588_ = ~new_n43932_ & ~new_n44581_;
  assign new_n44589_ = ~new_n44580_ & new_n44588_;
  assign new_n44590_ = ~new_n44587_ & ~new_n44589_;
  assign new_n44591_ = ~new_n43933_ & ~new_n44577_;
  assign new_n44592_ = ~new_n44575_ & new_n44591_;
  assign new_n44593_ = ~new_n44563_ & new_n44592_;
  assign new_n44594_ = ~new_n44575_ & ~new_n44577_;
  assign new_n44595_ = ~new_n44564_ & ~new_n44594_;
  assign new_n44596_ = ~new_n44593_ & ~new_n44595_;
  assign new_n44597_ = ~new_n44582_ & ~new_n44596_;
  assign new_n44598_ = ~new_n44574_ & ~new_n44581_;
  assign new_n44599_ = ~new_n44580_ & new_n44598_;
  assign new_n44600_ = ~new_n44597_ & ~new_n44599_;
  assign new_n44601_ = ~\b[48]  & ~new_n44600_;
  assign new_n44602_ = ~\b[47]  & ~new_n44590_;
  assign new_n44603_ = ~new_n43951_ & new_n44557_;
  assign new_n44604_ = ~new_n44553_ & new_n44603_;
  assign new_n44605_ = ~new_n44554_ & ~new_n44557_;
  assign new_n44606_ = ~new_n44604_ & ~new_n44605_;
  assign new_n44607_ = ~new_n44582_ & ~new_n44606_;
  assign new_n44608_ = ~new_n43941_ & ~new_n44581_;
  assign new_n44609_ = ~new_n44580_ & new_n44608_;
  assign new_n44610_ = ~new_n44607_ & ~new_n44609_;
  assign new_n44611_ = ~\b[46]  & ~new_n44610_;
  assign new_n44612_ = ~new_n43960_ & new_n44552_;
  assign new_n44613_ = ~new_n44548_ & new_n44612_;
  assign new_n44614_ = ~new_n44549_ & ~new_n44552_;
  assign new_n44615_ = ~new_n44613_ & ~new_n44614_;
  assign new_n44616_ = ~new_n44582_ & ~new_n44615_;
  assign new_n44617_ = ~new_n43950_ & ~new_n44581_;
  assign new_n44618_ = ~new_n44580_ & new_n44617_;
  assign new_n44619_ = ~new_n44616_ & ~new_n44618_;
  assign new_n44620_ = ~\b[45]  & ~new_n44619_;
  assign new_n44621_ = ~new_n43969_ & new_n44547_;
  assign new_n44622_ = ~new_n44543_ & new_n44621_;
  assign new_n44623_ = ~new_n44544_ & ~new_n44547_;
  assign new_n44624_ = ~new_n44622_ & ~new_n44623_;
  assign new_n44625_ = ~new_n44582_ & ~new_n44624_;
  assign new_n44626_ = ~new_n43959_ & ~new_n44581_;
  assign new_n44627_ = ~new_n44580_ & new_n44626_;
  assign new_n44628_ = ~new_n44625_ & ~new_n44627_;
  assign new_n44629_ = ~\b[44]  & ~new_n44628_;
  assign new_n44630_ = ~new_n43978_ & new_n44542_;
  assign new_n44631_ = ~new_n44538_ & new_n44630_;
  assign new_n44632_ = ~new_n44539_ & ~new_n44542_;
  assign new_n44633_ = ~new_n44631_ & ~new_n44632_;
  assign new_n44634_ = ~new_n44582_ & ~new_n44633_;
  assign new_n44635_ = ~new_n43968_ & ~new_n44581_;
  assign new_n44636_ = ~new_n44580_ & new_n44635_;
  assign new_n44637_ = ~new_n44634_ & ~new_n44636_;
  assign new_n44638_ = ~\b[43]  & ~new_n44637_;
  assign new_n44639_ = ~new_n43987_ & new_n44537_;
  assign new_n44640_ = ~new_n44533_ & new_n44639_;
  assign new_n44641_ = ~new_n44534_ & ~new_n44537_;
  assign new_n44642_ = ~new_n44640_ & ~new_n44641_;
  assign new_n44643_ = ~new_n44582_ & ~new_n44642_;
  assign new_n44644_ = ~new_n43977_ & ~new_n44581_;
  assign new_n44645_ = ~new_n44580_ & new_n44644_;
  assign new_n44646_ = ~new_n44643_ & ~new_n44645_;
  assign new_n44647_ = ~\b[42]  & ~new_n44646_;
  assign new_n44648_ = ~new_n43996_ & new_n44532_;
  assign new_n44649_ = ~new_n44528_ & new_n44648_;
  assign new_n44650_ = ~new_n44529_ & ~new_n44532_;
  assign new_n44651_ = ~new_n44649_ & ~new_n44650_;
  assign new_n44652_ = ~new_n44582_ & ~new_n44651_;
  assign new_n44653_ = ~new_n43986_ & ~new_n44581_;
  assign new_n44654_ = ~new_n44580_ & new_n44653_;
  assign new_n44655_ = ~new_n44652_ & ~new_n44654_;
  assign new_n44656_ = ~\b[41]  & ~new_n44655_;
  assign new_n44657_ = ~new_n44005_ & new_n44527_;
  assign new_n44658_ = ~new_n44523_ & new_n44657_;
  assign new_n44659_ = ~new_n44524_ & ~new_n44527_;
  assign new_n44660_ = ~new_n44658_ & ~new_n44659_;
  assign new_n44661_ = ~new_n44582_ & ~new_n44660_;
  assign new_n44662_ = ~new_n43995_ & ~new_n44581_;
  assign new_n44663_ = ~new_n44580_ & new_n44662_;
  assign new_n44664_ = ~new_n44661_ & ~new_n44663_;
  assign new_n44665_ = ~\b[40]  & ~new_n44664_;
  assign new_n44666_ = ~new_n44014_ & new_n44522_;
  assign new_n44667_ = ~new_n44518_ & new_n44666_;
  assign new_n44668_ = ~new_n44519_ & ~new_n44522_;
  assign new_n44669_ = ~new_n44667_ & ~new_n44668_;
  assign new_n44670_ = ~new_n44582_ & ~new_n44669_;
  assign new_n44671_ = ~new_n44004_ & ~new_n44581_;
  assign new_n44672_ = ~new_n44580_ & new_n44671_;
  assign new_n44673_ = ~new_n44670_ & ~new_n44672_;
  assign new_n44674_ = ~\b[39]  & ~new_n44673_;
  assign new_n44675_ = ~new_n44023_ & new_n44517_;
  assign new_n44676_ = ~new_n44513_ & new_n44675_;
  assign new_n44677_ = ~new_n44514_ & ~new_n44517_;
  assign new_n44678_ = ~new_n44676_ & ~new_n44677_;
  assign new_n44679_ = ~new_n44582_ & ~new_n44678_;
  assign new_n44680_ = ~new_n44013_ & ~new_n44581_;
  assign new_n44681_ = ~new_n44580_ & new_n44680_;
  assign new_n44682_ = ~new_n44679_ & ~new_n44681_;
  assign new_n44683_ = ~\b[38]  & ~new_n44682_;
  assign new_n44684_ = ~new_n44032_ & new_n44512_;
  assign new_n44685_ = ~new_n44508_ & new_n44684_;
  assign new_n44686_ = ~new_n44509_ & ~new_n44512_;
  assign new_n44687_ = ~new_n44685_ & ~new_n44686_;
  assign new_n44688_ = ~new_n44582_ & ~new_n44687_;
  assign new_n44689_ = ~new_n44022_ & ~new_n44581_;
  assign new_n44690_ = ~new_n44580_ & new_n44689_;
  assign new_n44691_ = ~new_n44688_ & ~new_n44690_;
  assign new_n44692_ = ~\b[37]  & ~new_n44691_;
  assign new_n44693_ = ~new_n44041_ & new_n44507_;
  assign new_n44694_ = ~new_n44503_ & new_n44693_;
  assign new_n44695_ = ~new_n44504_ & ~new_n44507_;
  assign new_n44696_ = ~new_n44694_ & ~new_n44695_;
  assign new_n44697_ = ~new_n44582_ & ~new_n44696_;
  assign new_n44698_ = ~new_n44031_ & ~new_n44581_;
  assign new_n44699_ = ~new_n44580_ & new_n44698_;
  assign new_n44700_ = ~new_n44697_ & ~new_n44699_;
  assign new_n44701_ = ~\b[36]  & ~new_n44700_;
  assign new_n44702_ = ~new_n44050_ & new_n44502_;
  assign new_n44703_ = ~new_n44498_ & new_n44702_;
  assign new_n44704_ = ~new_n44499_ & ~new_n44502_;
  assign new_n44705_ = ~new_n44703_ & ~new_n44704_;
  assign new_n44706_ = ~new_n44582_ & ~new_n44705_;
  assign new_n44707_ = ~new_n44040_ & ~new_n44581_;
  assign new_n44708_ = ~new_n44580_ & new_n44707_;
  assign new_n44709_ = ~new_n44706_ & ~new_n44708_;
  assign new_n44710_ = ~\b[35]  & ~new_n44709_;
  assign new_n44711_ = ~new_n44059_ & new_n44497_;
  assign new_n44712_ = ~new_n44493_ & new_n44711_;
  assign new_n44713_ = ~new_n44494_ & ~new_n44497_;
  assign new_n44714_ = ~new_n44712_ & ~new_n44713_;
  assign new_n44715_ = ~new_n44582_ & ~new_n44714_;
  assign new_n44716_ = ~new_n44049_ & ~new_n44581_;
  assign new_n44717_ = ~new_n44580_ & new_n44716_;
  assign new_n44718_ = ~new_n44715_ & ~new_n44717_;
  assign new_n44719_ = ~\b[34]  & ~new_n44718_;
  assign new_n44720_ = ~new_n44068_ & new_n44492_;
  assign new_n44721_ = ~new_n44488_ & new_n44720_;
  assign new_n44722_ = ~new_n44489_ & ~new_n44492_;
  assign new_n44723_ = ~new_n44721_ & ~new_n44722_;
  assign new_n44724_ = ~new_n44582_ & ~new_n44723_;
  assign new_n44725_ = ~new_n44058_ & ~new_n44581_;
  assign new_n44726_ = ~new_n44580_ & new_n44725_;
  assign new_n44727_ = ~new_n44724_ & ~new_n44726_;
  assign new_n44728_ = ~\b[33]  & ~new_n44727_;
  assign new_n44729_ = ~new_n44077_ & new_n44487_;
  assign new_n44730_ = ~new_n44483_ & new_n44729_;
  assign new_n44731_ = ~new_n44484_ & ~new_n44487_;
  assign new_n44732_ = ~new_n44730_ & ~new_n44731_;
  assign new_n44733_ = ~new_n44582_ & ~new_n44732_;
  assign new_n44734_ = ~new_n44067_ & ~new_n44581_;
  assign new_n44735_ = ~new_n44580_ & new_n44734_;
  assign new_n44736_ = ~new_n44733_ & ~new_n44735_;
  assign new_n44737_ = ~\b[32]  & ~new_n44736_;
  assign new_n44738_ = ~new_n44086_ & new_n44482_;
  assign new_n44739_ = ~new_n44478_ & new_n44738_;
  assign new_n44740_ = ~new_n44479_ & ~new_n44482_;
  assign new_n44741_ = ~new_n44739_ & ~new_n44740_;
  assign new_n44742_ = ~new_n44582_ & ~new_n44741_;
  assign new_n44743_ = ~new_n44076_ & ~new_n44581_;
  assign new_n44744_ = ~new_n44580_ & new_n44743_;
  assign new_n44745_ = ~new_n44742_ & ~new_n44744_;
  assign new_n44746_ = ~\b[31]  & ~new_n44745_;
  assign new_n44747_ = ~new_n44095_ & new_n44477_;
  assign new_n44748_ = ~new_n44473_ & new_n44747_;
  assign new_n44749_ = ~new_n44474_ & ~new_n44477_;
  assign new_n44750_ = ~new_n44748_ & ~new_n44749_;
  assign new_n44751_ = ~new_n44582_ & ~new_n44750_;
  assign new_n44752_ = ~new_n44085_ & ~new_n44581_;
  assign new_n44753_ = ~new_n44580_ & new_n44752_;
  assign new_n44754_ = ~new_n44751_ & ~new_n44753_;
  assign new_n44755_ = ~\b[30]  & ~new_n44754_;
  assign new_n44756_ = ~new_n44104_ & new_n44472_;
  assign new_n44757_ = ~new_n44468_ & new_n44756_;
  assign new_n44758_ = ~new_n44469_ & ~new_n44472_;
  assign new_n44759_ = ~new_n44757_ & ~new_n44758_;
  assign new_n44760_ = ~new_n44582_ & ~new_n44759_;
  assign new_n44761_ = ~new_n44094_ & ~new_n44581_;
  assign new_n44762_ = ~new_n44580_ & new_n44761_;
  assign new_n44763_ = ~new_n44760_ & ~new_n44762_;
  assign new_n44764_ = ~\b[29]  & ~new_n44763_;
  assign new_n44765_ = ~new_n44113_ & new_n44467_;
  assign new_n44766_ = ~new_n44463_ & new_n44765_;
  assign new_n44767_ = ~new_n44464_ & ~new_n44467_;
  assign new_n44768_ = ~new_n44766_ & ~new_n44767_;
  assign new_n44769_ = ~new_n44582_ & ~new_n44768_;
  assign new_n44770_ = ~new_n44103_ & ~new_n44581_;
  assign new_n44771_ = ~new_n44580_ & new_n44770_;
  assign new_n44772_ = ~new_n44769_ & ~new_n44771_;
  assign new_n44773_ = ~\b[28]  & ~new_n44772_;
  assign new_n44774_ = ~new_n44122_ & new_n44462_;
  assign new_n44775_ = ~new_n44458_ & new_n44774_;
  assign new_n44776_ = ~new_n44459_ & ~new_n44462_;
  assign new_n44777_ = ~new_n44775_ & ~new_n44776_;
  assign new_n44778_ = ~new_n44582_ & ~new_n44777_;
  assign new_n44779_ = ~new_n44112_ & ~new_n44581_;
  assign new_n44780_ = ~new_n44580_ & new_n44779_;
  assign new_n44781_ = ~new_n44778_ & ~new_n44780_;
  assign new_n44782_ = ~\b[27]  & ~new_n44781_;
  assign new_n44783_ = ~new_n44131_ & new_n44457_;
  assign new_n44784_ = ~new_n44453_ & new_n44783_;
  assign new_n44785_ = ~new_n44454_ & ~new_n44457_;
  assign new_n44786_ = ~new_n44784_ & ~new_n44785_;
  assign new_n44787_ = ~new_n44582_ & ~new_n44786_;
  assign new_n44788_ = ~new_n44121_ & ~new_n44581_;
  assign new_n44789_ = ~new_n44580_ & new_n44788_;
  assign new_n44790_ = ~new_n44787_ & ~new_n44789_;
  assign new_n44791_ = ~\b[26]  & ~new_n44790_;
  assign new_n44792_ = ~new_n44140_ & new_n44452_;
  assign new_n44793_ = ~new_n44448_ & new_n44792_;
  assign new_n44794_ = ~new_n44449_ & ~new_n44452_;
  assign new_n44795_ = ~new_n44793_ & ~new_n44794_;
  assign new_n44796_ = ~new_n44582_ & ~new_n44795_;
  assign new_n44797_ = ~new_n44130_ & ~new_n44581_;
  assign new_n44798_ = ~new_n44580_ & new_n44797_;
  assign new_n44799_ = ~new_n44796_ & ~new_n44798_;
  assign new_n44800_ = ~\b[25]  & ~new_n44799_;
  assign new_n44801_ = ~new_n44149_ & new_n44447_;
  assign new_n44802_ = ~new_n44443_ & new_n44801_;
  assign new_n44803_ = ~new_n44444_ & ~new_n44447_;
  assign new_n44804_ = ~new_n44802_ & ~new_n44803_;
  assign new_n44805_ = ~new_n44582_ & ~new_n44804_;
  assign new_n44806_ = ~new_n44139_ & ~new_n44581_;
  assign new_n44807_ = ~new_n44580_ & new_n44806_;
  assign new_n44808_ = ~new_n44805_ & ~new_n44807_;
  assign new_n44809_ = ~\b[24]  & ~new_n44808_;
  assign new_n44810_ = ~new_n44158_ & new_n44442_;
  assign new_n44811_ = ~new_n44438_ & new_n44810_;
  assign new_n44812_ = ~new_n44439_ & ~new_n44442_;
  assign new_n44813_ = ~new_n44811_ & ~new_n44812_;
  assign new_n44814_ = ~new_n44582_ & ~new_n44813_;
  assign new_n44815_ = ~new_n44148_ & ~new_n44581_;
  assign new_n44816_ = ~new_n44580_ & new_n44815_;
  assign new_n44817_ = ~new_n44814_ & ~new_n44816_;
  assign new_n44818_ = ~\b[23]  & ~new_n44817_;
  assign new_n44819_ = ~new_n44167_ & new_n44437_;
  assign new_n44820_ = ~new_n44433_ & new_n44819_;
  assign new_n44821_ = ~new_n44434_ & ~new_n44437_;
  assign new_n44822_ = ~new_n44820_ & ~new_n44821_;
  assign new_n44823_ = ~new_n44582_ & ~new_n44822_;
  assign new_n44824_ = ~new_n44157_ & ~new_n44581_;
  assign new_n44825_ = ~new_n44580_ & new_n44824_;
  assign new_n44826_ = ~new_n44823_ & ~new_n44825_;
  assign new_n44827_ = ~\b[22]  & ~new_n44826_;
  assign new_n44828_ = ~new_n44176_ & new_n44432_;
  assign new_n44829_ = ~new_n44428_ & new_n44828_;
  assign new_n44830_ = ~new_n44429_ & ~new_n44432_;
  assign new_n44831_ = ~new_n44829_ & ~new_n44830_;
  assign new_n44832_ = ~new_n44582_ & ~new_n44831_;
  assign new_n44833_ = ~new_n44166_ & ~new_n44581_;
  assign new_n44834_ = ~new_n44580_ & new_n44833_;
  assign new_n44835_ = ~new_n44832_ & ~new_n44834_;
  assign new_n44836_ = ~\b[21]  & ~new_n44835_;
  assign new_n44837_ = ~new_n44185_ & new_n44427_;
  assign new_n44838_ = ~new_n44423_ & new_n44837_;
  assign new_n44839_ = ~new_n44424_ & ~new_n44427_;
  assign new_n44840_ = ~new_n44838_ & ~new_n44839_;
  assign new_n44841_ = ~new_n44582_ & ~new_n44840_;
  assign new_n44842_ = ~new_n44175_ & ~new_n44581_;
  assign new_n44843_ = ~new_n44580_ & new_n44842_;
  assign new_n44844_ = ~new_n44841_ & ~new_n44843_;
  assign new_n44845_ = ~\b[20]  & ~new_n44844_;
  assign new_n44846_ = ~new_n44194_ & new_n44422_;
  assign new_n44847_ = ~new_n44418_ & new_n44846_;
  assign new_n44848_ = ~new_n44419_ & ~new_n44422_;
  assign new_n44849_ = ~new_n44847_ & ~new_n44848_;
  assign new_n44850_ = ~new_n44582_ & ~new_n44849_;
  assign new_n44851_ = ~new_n44184_ & ~new_n44581_;
  assign new_n44852_ = ~new_n44580_ & new_n44851_;
  assign new_n44853_ = ~new_n44850_ & ~new_n44852_;
  assign new_n44854_ = ~\b[19]  & ~new_n44853_;
  assign new_n44855_ = ~new_n44203_ & new_n44417_;
  assign new_n44856_ = ~new_n44413_ & new_n44855_;
  assign new_n44857_ = ~new_n44414_ & ~new_n44417_;
  assign new_n44858_ = ~new_n44856_ & ~new_n44857_;
  assign new_n44859_ = ~new_n44582_ & ~new_n44858_;
  assign new_n44860_ = ~new_n44193_ & ~new_n44581_;
  assign new_n44861_ = ~new_n44580_ & new_n44860_;
  assign new_n44862_ = ~new_n44859_ & ~new_n44861_;
  assign new_n44863_ = ~\b[18]  & ~new_n44862_;
  assign new_n44864_ = ~new_n44212_ & new_n44412_;
  assign new_n44865_ = ~new_n44408_ & new_n44864_;
  assign new_n44866_ = ~new_n44409_ & ~new_n44412_;
  assign new_n44867_ = ~new_n44865_ & ~new_n44866_;
  assign new_n44868_ = ~new_n44582_ & ~new_n44867_;
  assign new_n44869_ = ~new_n44202_ & ~new_n44581_;
  assign new_n44870_ = ~new_n44580_ & new_n44869_;
  assign new_n44871_ = ~new_n44868_ & ~new_n44870_;
  assign new_n44872_ = ~\b[17]  & ~new_n44871_;
  assign new_n44873_ = ~new_n44221_ & new_n44407_;
  assign new_n44874_ = ~new_n44403_ & new_n44873_;
  assign new_n44875_ = ~new_n44404_ & ~new_n44407_;
  assign new_n44876_ = ~new_n44874_ & ~new_n44875_;
  assign new_n44877_ = ~new_n44582_ & ~new_n44876_;
  assign new_n44878_ = ~new_n44211_ & ~new_n44581_;
  assign new_n44879_ = ~new_n44580_ & new_n44878_;
  assign new_n44880_ = ~new_n44877_ & ~new_n44879_;
  assign new_n44881_ = ~\b[16]  & ~new_n44880_;
  assign new_n44882_ = ~new_n44230_ & new_n44402_;
  assign new_n44883_ = ~new_n44398_ & new_n44882_;
  assign new_n44884_ = ~new_n44399_ & ~new_n44402_;
  assign new_n44885_ = ~new_n44883_ & ~new_n44884_;
  assign new_n44886_ = ~new_n44582_ & ~new_n44885_;
  assign new_n44887_ = ~new_n44220_ & ~new_n44581_;
  assign new_n44888_ = ~new_n44580_ & new_n44887_;
  assign new_n44889_ = ~new_n44886_ & ~new_n44888_;
  assign new_n44890_ = ~\b[15]  & ~new_n44889_;
  assign new_n44891_ = ~new_n44239_ & new_n44397_;
  assign new_n44892_ = ~new_n44393_ & new_n44891_;
  assign new_n44893_ = ~new_n44394_ & ~new_n44397_;
  assign new_n44894_ = ~new_n44892_ & ~new_n44893_;
  assign new_n44895_ = ~new_n44582_ & ~new_n44894_;
  assign new_n44896_ = ~new_n44229_ & ~new_n44581_;
  assign new_n44897_ = ~new_n44580_ & new_n44896_;
  assign new_n44898_ = ~new_n44895_ & ~new_n44897_;
  assign new_n44899_ = ~\b[14]  & ~new_n44898_;
  assign new_n44900_ = ~new_n44248_ & new_n44392_;
  assign new_n44901_ = ~new_n44388_ & new_n44900_;
  assign new_n44902_ = ~new_n44389_ & ~new_n44392_;
  assign new_n44903_ = ~new_n44901_ & ~new_n44902_;
  assign new_n44904_ = ~new_n44582_ & ~new_n44903_;
  assign new_n44905_ = ~new_n44238_ & ~new_n44581_;
  assign new_n44906_ = ~new_n44580_ & new_n44905_;
  assign new_n44907_ = ~new_n44904_ & ~new_n44906_;
  assign new_n44908_ = ~\b[13]  & ~new_n44907_;
  assign new_n44909_ = ~new_n44257_ & new_n44387_;
  assign new_n44910_ = ~new_n44383_ & new_n44909_;
  assign new_n44911_ = ~new_n44384_ & ~new_n44387_;
  assign new_n44912_ = ~new_n44910_ & ~new_n44911_;
  assign new_n44913_ = ~new_n44582_ & ~new_n44912_;
  assign new_n44914_ = ~new_n44247_ & ~new_n44581_;
  assign new_n44915_ = ~new_n44580_ & new_n44914_;
  assign new_n44916_ = ~new_n44913_ & ~new_n44915_;
  assign new_n44917_ = ~\b[12]  & ~new_n44916_;
  assign new_n44918_ = ~new_n44266_ & new_n44382_;
  assign new_n44919_ = ~new_n44378_ & new_n44918_;
  assign new_n44920_ = ~new_n44379_ & ~new_n44382_;
  assign new_n44921_ = ~new_n44919_ & ~new_n44920_;
  assign new_n44922_ = ~new_n44582_ & ~new_n44921_;
  assign new_n44923_ = ~new_n44256_ & ~new_n44581_;
  assign new_n44924_ = ~new_n44580_ & new_n44923_;
  assign new_n44925_ = ~new_n44922_ & ~new_n44924_;
  assign new_n44926_ = ~\b[11]  & ~new_n44925_;
  assign new_n44927_ = ~new_n44275_ & new_n44377_;
  assign new_n44928_ = ~new_n44373_ & new_n44927_;
  assign new_n44929_ = ~new_n44374_ & ~new_n44377_;
  assign new_n44930_ = ~new_n44928_ & ~new_n44929_;
  assign new_n44931_ = ~new_n44582_ & ~new_n44930_;
  assign new_n44932_ = ~new_n44265_ & ~new_n44581_;
  assign new_n44933_ = ~new_n44580_ & new_n44932_;
  assign new_n44934_ = ~new_n44931_ & ~new_n44933_;
  assign new_n44935_ = ~\b[10]  & ~new_n44934_;
  assign new_n44936_ = ~new_n44284_ & new_n44372_;
  assign new_n44937_ = ~new_n44368_ & new_n44936_;
  assign new_n44938_ = ~new_n44369_ & ~new_n44372_;
  assign new_n44939_ = ~new_n44937_ & ~new_n44938_;
  assign new_n44940_ = ~new_n44582_ & ~new_n44939_;
  assign new_n44941_ = ~new_n44274_ & ~new_n44581_;
  assign new_n44942_ = ~new_n44580_ & new_n44941_;
  assign new_n44943_ = ~new_n44940_ & ~new_n44942_;
  assign new_n44944_ = ~\b[9]  & ~new_n44943_;
  assign new_n44945_ = ~new_n44293_ & new_n44367_;
  assign new_n44946_ = ~new_n44363_ & new_n44945_;
  assign new_n44947_ = ~new_n44364_ & ~new_n44367_;
  assign new_n44948_ = ~new_n44946_ & ~new_n44947_;
  assign new_n44949_ = ~new_n44582_ & ~new_n44948_;
  assign new_n44950_ = ~new_n44283_ & ~new_n44581_;
  assign new_n44951_ = ~new_n44580_ & new_n44950_;
  assign new_n44952_ = ~new_n44949_ & ~new_n44951_;
  assign new_n44953_ = ~\b[8]  & ~new_n44952_;
  assign new_n44954_ = ~new_n44302_ & new_n44362_;
  assign new_n44955_ = ~new_n44358_ & new_n44954_;
  assign new_n44956_ = ~new_n44359_ & ~new_n44362_;
  assign new_n44957_ = ~new_n44955_ & ~new_n44956_;
  assign new_n44958_ = ~new_n44582_ & ~new_n44957_;
  assign new_n44959_ = ~new_n44292_ & ~new_n44581_;
  assign new_n44960_ = ~new_n44580_ & new_n44959_;
  assign new_n44961_ = ~new_n44958_ & ~new_n44960_;
  assign new_n44962_ = ~\b[7]  & ~new_n44961_;
  assign new_n44963_ = ~new_n44311_ & new_n44357_;
  assign new_n44964_ = ~new_n44353_ & new_n44963_;
  assign new_n44965_ = ~new_n44354_ & ~new_n44357_;
  assign new_n44966_ = ~new_n44964_ & ~new_n44965_;
  assign new_n44967_ = ~new_n44582_ & ~new_n44966_;
  assign new_n44968_ = ~new_n44301_ & ~new_n44581_;
  assign new_n44969_ = ~new_n44580_ & new_n44968_;
  assign new_n44970_ = ~new_n44967_ & ~new_n44969_;
  assign new_n44971_ = ~\b[6]  & ~new_n44970_;
  assign new_n44972_ = ~new_n44320_ & new_n44352_;
  assign new_n44973_ = ~new_n44348_ & new_n44972_;
  assign new_n44974_ = ~new_n44349_ & ~new_n44352_;
  assign new_n44975_ = ~new_n44973_ & ~new_n44974_;
  assign new_n44976_ = ~new_n44582_ & ~new_n44975_;
  assign new_n44977_ = ~new_n44310_ & ~new_n44581_;
  assign new_n44978_ = ~new_n44580_ & new_n44977_;
  assign new_n44979_ = ~new_n44976_ & ~new_n44978_;
  assign new_n44980_ = ~\b[5]  & ~new_n44979_;
  assign new_n44981_ = ~new_n44328_ & new_n44347_;
  assign new_n44982_ = ~new_n44343_ & new_n44981_;
  assign new_n44983_ = ~new_n44344_ & ~new_n44347_;
  assign new_n44984_ = ~new_n44982_ & ~new_n44983_;
  assign new_n44985_ = ~new_n44582_ & ~new_n44984_;
  assign new_n44986_ = ~new_n44319_ & ~new_n44581_;
  assign new_n44987_ = ~new_n44580_ & new_n44986_;
  assign new_n44988_ = ~new_n44985_ & ~new_n44987_;
  assign new_n44989_ = ~\b[4]  & ~new_n44988_;
  assign new_n44990_ = ~new_n44338_ & new_n44342_;
  assign new_n44991_ = ~new_n44337_ & new_n44990_;
  assign new_n44992_ = ~new_n44339_ & ~new_n44342_;
  assign new_n44993_ = ~new_n44991_ & ~new_n44992_;
  assign new_n44994_ = ~new_n44582_ & ~new_n44993_;
  assign new_n44995_ = ~new_n44327_ & ~new_n44581_;
  assign new_n44996_ = ~new_n44580_ & new_n44995_;
  assign new_n44997_ = ~new_n44994_ & ~new_n44996_;
  assign new_n44998_ = ~\b[3]  & ~new_n44997_;
  assign new_n44999_ = new_n16277_ & ~new_n44335_;
  assign new_n45000_ = ~new_n44333_ & new_n44999_;
  assign new_n45001_ = ~new_n44337_ & ~new_n45000_;
  assign new_n45002_ = ~new_n44582_ & new_n45001_;
  assign new_n45003_ = ~new_n44332_ & ~new_n44581_;
  assign new_n45004_ = ~new_n44580_ & new_n45003_;
  assign new_n45005_ = ~new_n45002_ & ~new_n45004_;
  assign new_n45006_ = ~\b[2]  & ~new_n45005_;
  assign new_n45007_ = \b[0]  & ~new_n44582_;
  assign new_n45008_ = \a[16]  & ~new_n45007_;
  assign new_n45009_ = new_n16277_ & ~new_n44582_;
  assign new_n45010_ = ~new_n45008_ & ~new_n45009_;
  assign new_n45011_ = \b[1]  & ~new_n45010_;
  assign new_n45012_ = ~\b[1]  & ~new_n45009_;
  assign new_n45013_ = ~new_n45008_ & new_n45012_;
  assign new_n45014_ = ~new_n45011_ & ~new_n45013_;
  assign new_n45015_ = ~new_n16956_ & ~new_n45014_;
  assign new_n45016_ = ~\b[1]  & ~new_n45010_;
  assign new_n45017_ = ~new_n45015_ & ~new_n45016_;
  assign new_n45018_ = \b[2]  & ~new_n45004_;
  assign new_n45019_ = ~new_n45002_ & new_n45018_;
  assign new_n45020_ = ~new_n45006_ & ~new_n45019_;
  assign new_n45021_ = ~new_n45017_ & new_n45020_;
  assign new_n45022_ = ~new_n45006_ & ~new_n45021_;
  assign new_n45023_ = \b[3]  & ~new_n44996_;
  assign new_n45024_ = ~new_n44994_ & new_n45023_;
  assign new_n45025_ = ~new_n44998_ & ~new_n45024_;
  assign new_n45026_ = ~new_n45022_ & new_n45025_;
  assign new_n45027_ = ~new_n44998_ & ~new_n45026_;
  assign new_n45028_ = \b[4]  & ~new_n44987_;
  assign new_n45029_ = ~new_n44985_ & new_n45028_;
  assign new_n45030_ = ~new_n44989_ & ~new_n45029_;
  assign new_n45031_ = ~new_n45027_ & new_n45030_;
  assign new_n45032_ = ~new_n44989_ & ~new_n45031_;
  assign new_n45033_ = \b[5]  & ~new_n44978_;
  assign new_n45034_ = ~new_n44976_ & new_n45033_;
  assign new_n45035_ = ~new_n44980_ & ~new_n45034_;
  assign new_n45036_ = ~new_n45032_ & new_n45035_;
  assign new_n45037_ = ~new_n44980_ & ~new_n45036_;
  assign new_n45038_ = \b[6]  & ~new_n44969_;
  assign new_n45039_ = ~new_n44967_ & new_n45038_;
  assign new_n45040_ = ~new_n44971_ & ~new_n45039_;
  assign new_n45041_ = ~new_n45037_ & new_n45040_;
  assign new_n45042_ = ~new_n44971_ & ~new_n45041_;
  assign new_n45043_ = \b[7]  & ~new_n44960_;
  assign new_n45044_ = ~new_n44958_ & new_n45043_;
  assign new_n45045_ = ~new_n44962_ & ~new_n45044_;
  assign new_n45046_ = ~new_n45042_ & new_n45045_;
  assign new_n45047_ = ~new_n44962_ & ~new_n45046_;
  assign new_n45048_ = \b[8]  & ~new_n44951_;
  assign new_n45049_ = ~new_n44949_ & new_n45048_;
  assign new_n45050_ = ~new_n44953_ & ~new_n45049_;
  assign new_n45051_ = ~new_n45047_ & new_n45050_;
  assign new_n45052_ = ~new_n44953_ & ~new_n45051_;
  assign new_n45053_ = \b[9]  & ~new_n44942_;
  assign new_n45054_ = ~new_n44940_ & new_n45053_;
  assign new_n45055_ = ~new_n44944_ & ~new_n45054_;
  assign new_n45056_ = ~new_n45052_ & new_n45055_;
  assign new_n45057_ = ~new_n44944_ & ~new_n45056_;
  assign new_n45058_ = \b[10]  & ~new_n44933_;
  assign new_n45059_ = ~new_n44931_ & new_n45058_;
  assign new_n45060_ = ~new_n44935_ & ~new_n45059_;
  assign new_n45061_ = ~new_n45057_ & new_n45060_;
  assign new_n45062_ = ~new_n44935_ & ~new_n45061_;
  assign new_n45063_ = \b[11]  & ~new_n44924_;
  assign new_n45064_ = ~new_n44922_ & new_n45063_;
  assign new_n45065_ = ~new_n44926_ & ~new_n45064_;
  assign new_n45066_ = ~new_n45062_ & new_n45065_;
  assign new_n45067_ = ~new_n44926_ & ~new_n45066_;
  assign new_n45068_ = \b[12]  & ~new_n44915_;
  assign new_n45069_ = ~new_n44913_ & new_n45068_;
  assign new_n45070_ = ~new_n44917_ & ~new_n45069_;
  assign new_n45071_ = ~new_n45067_ & new_n45070_;
  assign new_n45072_ = ~new_n44917_ & ~new_n45071_;
  assign new_n45073_ = \b[13]  & ~new_n44906_;
  assign new_n45074_ = ~new_n44904_ & new_n45073_;
  assign new_n45075_ = ~new_n44908_ & ~new_n45074_;
  assign new_n45076_ = ~new_n45072_ & new_n45075_;
  assign new_n45077_ = ~new_n44908_ & ~new_n45076_;
  assign new_n45078_ = \b[14]  & ~new_n44897_;
  assign new_n45079_ = ~new_n44895_ & new_n45078_;
  assign new_n45080_ = ~new_n44899_ & ~new_n45079_;
  assign new_n45081_ = ~new_n45077_ & new_n45080_;
  assign new_n45082_ = ~new_n44899_ & ~new_n45081_;
  assign new_n45083_ = \b[15]  & ~new_n44888_;
  assign new_n45084_ = ~new_n44886_ & new_n45083_;
  assign new_n45085_ = ~new_n44890_ & ~new_n45084_;
  assign new_n45086_ = ~new_n45082_ & new_n45085_;
  assign new_n45087_ = ~new_n44890_ & ~new_n45086_;
  assign new_n45088_ = \b[16]  & ~new_n44879_;
  assign new_n45089_ = ~new_n44877_ & new_n45088_;
  assign new_n45090_ = ~new_n44881_ & ~new_n45089_;
  assign new_n45091_ = ~new_n45087_ & new_n45090_;
  assign new_n45092_ = ~new_n44881_ & ~new_n45091_;
  assign new_n45093_ = \b[17]  & ~new_n44870_;
  assign new_n45094_ = ~new_n44868_ & new_n45093_;
  assign new_n45095_ = ~new_n44872_ & ~new_n45094_;
  assign new_n45096_ = ~new_n45092_ & new_n45095_;
  assign new_n45097_ = ~new_n44872_ & ~new_n45096_;
  assign new_n45098_ = \b[18]  & ~new_n44861_;
  assign new_n45099_ = ~new_n44859_ & new_n45098_;
  assign new_n45100_ = ~new_n44863_ & ~new_n45099_;
  assign new_n45101_ = ~new_n45097_ & new_n45100_;
  assign new_n45102_ = ~new_n44863_ & ~new_n45101_;
  assign new_n45103_ = \b[19]  & ~new_n44852_;
  assign new_n45104_ = ~new_n44850_ & new_n45103_;
  assign new_n45105_ = ~new_n44854_ & ~new_n45104_;
  assign new_n45106_ = ~new_n45102_ & new_n45105_;
  assign new_n45107_ = ~new_n44854_ & ~new_n45106_;
  assign new_n45108_ = \b[20]  & ~new_n44843_;
  assign new_n45109_ = ~new_n44841_ & new_n45108_;
  assign new_n45110_ = ~new_n44845_ & ~new_n45109_;
  assign new_n45111_ = ~new_n45107_ & new_n45110_;
  assign new_n45112_ = ~new_n44845_ & ~new_n45111_;
  assign new_n45113_ = \b[21]  & ~new_n44834_;
  assign new_n45114_ = ~new_n44832_ & new_n45113_;
  assign new_n45115_ = ~new_n44836_ & ~new_n45114_;
  assign new_n45116_ = ~new_n45112_ & new_n45115_;
  assign new_n45117_ = ~new_n44836_ & ~new_n45116_;
  assign new_n45118_ = \b[22]  & ~new_n44825_;
  assign new_n45119_ = ~new_n44823_ & new_n45118_;
  assign new_n45120_ = ~new_n44827_ & ~new_n45119_;
  assign new_n45121_ = ~new_n45117_ & new_n45120_;
  assign new_n45122_ = ~new_n44827_ & ~new_n45121_;
  assign new_n45123_ = \b[23]  & ~new_n44816_;
  assign new_n45124_ = ~new_n44814_ & new_n45123_;
  assign new_n45125_ = ~new_n44818_ & ~new_n45124_;
  assign new_n45126_ = ~new_n45122_ & new_n45125_;
  assign new_n45127_ = ~new_n44818_ & ~new_n45126_;
  assign new_n45128_ = \b[24]  & ~new_n44807_;
  assign new_n45129_ = ~new_n44805_ & new_n45128_;
  assign new_n45130_ = ~new_n44809_ & ~new_n45129_;
  assign new_n45131_ = ~new_n45127_ & new_n45130_;
  assign new_n45132_ = ~new_n44809_ & ~new_n45131_;
  assign new_n45133_ = \b[25]  & ~new_n44798_;
  assign new_n45134_ = ~new_n44796_ & new_n45133_;
  assign new_n45135_ = ~new_n44800_ & ~new_n45134_;
  assign new_n45136_ = ~new_n45132_ & new_n45135_;
  assign new_n45137_ = ~new_n44800_ & ~new_n45136_;
  assign new_n45138_ = \b[26]  & ~new_n44789_;
  assign new_n45139_ = ~new_n44787_ & new_n45138_;
  assign new_n45140_ = ~new_n44791_ & ~new_n45139_;
  assign new_n45141_ = ~new_n45137_ & new_n45140_;
  assign new_n45142_ = ~new_n44791_ & ~new_n45141_;
  assign new_n45143_ = \b[27]  & ~new_n44780_;
  assign new_n45144_ = ~new_n44778_ & new_n45143_;
  assign new_n45145_ = ~new_n44782_ & ~new_n45144_;
  assign new_n45146_ = ~new_n45142_ & new_n45145_;
  assign new_n45147_ = ~new_n44782_ & ~new_n45146_;
  assign new_n45148_ = \b[28]  & ~new_n44771_;
  assign new_n45149_ = ~new_n44769_ & new_n45148_;
  assign new_n45150_ = ~new_n44773_ & ~new_n45149_;
  assign new_n45151_ = ~new_n45147_ & new_n45150_;
  assign new_n45152_ = ~new_n44773_ & ~new_n45151_;
  assign new_n45153_ = \b[29]  & ~new_n44762_;
  assign new_n45154_ = ~new_n44760_ & new_n45153_;
  assign new_n45155_ = ~new_n44764_ & ~new_n45154_;
  assign new_n45156_ = ~new_n45152_ & new_n45155_;
  assign new_n45157_ = ~new_n44764_ & ~new_n45156_;
  assign new_n45158_ = \b[30]  & ~new_n44753_;
  assign new_n45159_ = ~new_n44751_ & new_n45158_;
  assign new_n45160_ = ~new_n44755_ & ~new_n45159_;
  assign new_n45161_ = ~new_n45157_ & new_n45160_;
  assign new_n45162_ = ~new_n44755_ & ~new_n45161_;
  assign new_n45163_ = \b[31]  & ~new_n44744_;
  assign new_n45164_ = ~new_n44742_ & new_n45163_;
  assign new_n45165_ = ~new_n44746_ & ~new_n45164_;
  assign new_n45166_ = ~new_n45162_ & new_n45165_;
  assign new_n45167_ = ~new_n44746_ & ~new_n45166_;
  assign new_n45168_ = \b[32]  & ~new_n44735_;
  assign new_n45169_ = ~new_n44733_ & new_n45168_;
  assign new_n45170_ = ~new_n44737_ & ~new_n45169_;
  assign new_n45171_ = ~new_n45167_ & new_n45170_;
  assign new_n45172_ = ~new_n44737_ & ~new_n45171_;
  assign new_n45173_ = \b[33]  & ~new_n44726_;
  assign new_n45174_ = ~new_n44724_ & new_n45173_;
  assign new_n45175_ = ~new_n44728_ & ~new_n45174_;
  assign new_n45176_ = ~new_n45172_ & new_n45175_;
  assign new_n45177_ = ~new_n44728_ & ~new_n45176_;
  assign new_n45178_ = \b[34]  & ~new_n44717_;
  assign new_n45179_ = ~new_n44715_ & new_n45178_;
  assign new_n45180_ = ~new_n44719_ & ~new_n45179_;
  assign new_n45181_ = ~new_n45177_ & new_n45180_;
  assign new_n45182_ = ~new_n44719_ & ~new_n45181_;
  assign new_n45183_ = \b[35]  & ~new_n44708_;
  assign new_n45184_ = ~new_n44706_ & new_n45183_;
  assign new_n45185_ = ~new_n44710_ & ~new_n45184_;
  assign new_n45186_ = ~new_n45182_ & new_n45185_;
  assign new_n45187_ = ~new_n44710_ & ~new_n45186_;
  assign new_n45188_ = \b[36]  & ~new_n44699_;
  assign new_n45189_ = ~new_n44697_ & new_n45188_;
  assign new_n45190_ = ~new_n44701_ & ~new_n45189_;
  assign new_n45191_ = ~new_n45187_ & new_n45190_;
  assign new_n45192_ = ~new_n44701_ & ~new_n45191_;
  assign new_n45193_ = \b[37]  & ~new_n44690_;
  assign new_n45194_ = ~new_n44688_ & new_n45193_;
  assign new_n45195_ = ~new_n44692_ & ~new_n45194_;
  assign new_n45196_ = ~new_n45192_ & new_n45195_;
  assign new_n45197_ = ~new_n44692_ & ~new_n45196_;
  assign new_n45198_ = \b[38]  & ~new_n44681_;
  assign new_n45199_ = ~new_n44679_ & new_n45198_;
  assign new_n45200_ = ~new_n44683_ & ~new_n45199_;
  assign new_n45201_ = ~new_n45197_ & new_n45200_;
  assign new_n45202_ = ~new_n44683_ & ~new_n45201_;
  assign new_n45203_ = \b[39]  & ~new_n44672_;
  assign new_n45204_ = ~new_n44670_ & new_n45203_;
  assign new_n45205_ = ~new_n44674_ & ~new_n45204_;
  assign new_n45206_ = ~new_n45202_ & new_n45205_;
  assign new_n45207_ = ~new_n44674_ & ~new_n45206_;
  assign new_n45208_ = \b[40]  & ~new_n44663_;
  assign new_n45209_ = ~new_n44661_ & new_n45208_;
  assign new_n45210_ = ~new_n44665_ & ~new_n45209_;
  assign new_n45211_ = ~new_n45207_ & new_n45210_;
  assign new_n45212_ = ~new_n44665_ & ~new_n45211_;
  assign new_n45213_ = \b[41]  & ~new_n44654_;
  assign new_n45214_ = ~new_n44652_ & new_n45213_;
  assign new_n45215_ = ~new_n44656_ & ~new_n45214_;
  assign new_n45216_ = ~new_n45212_ & new_n45215_;
  assign new_n45217_ = ~new_n44656_ & ~new_n45216_;
  assign new_n45218_ = \b[42]  & ~new_n44645_;
  assign new_n45219_ = ~new_n44643_ & new_n45218_;
  assign new_n45220_ = ~new_n44647_ & ~new_n45219_;
  assign new_n45221_ = ~new_n45217_ & new_n45220_;
  assign new_n45222_ = ~new_n44647_ & ~new_n45221_;
  assign new_n45223_ = \b[43]  & ~new_n44636_;
  assign new_n45224_ = ~new_n44634_ & new_n45223_;
  assign new_n45225_ = ~new_n44638_ & ~new_n45224_;
  assign new_n45226_ = ~new_n45222_ & new_n45225_;
  assign new_n45227_ = ~new_n44638_ & ~new_n45226_;
  assign new_n45228_ = \b[44]  & ~new_n44627_;
  assign new_n45229_ = ~new_n44625_ & new_n45228_;
  assign new_n45230_ = ~new_n44629_ & ~new_n45229_;
  assign new_n45231_ = ~new_n45227_ & new_n45230_;
  assign new_n45232_ = ~new_n44629_ & ~new_n45231_;
  assign new_n45233_ = \b[45]  & ~new_n44618_;
  assign new_n45234_ = ~new_n44616_ & new_n45233_;
  assign new_n45235_ = ~new_n44620_ & ~new_n45234_;
  assign new_n45236_ = ~new_n45232_ & new_n45235_;
  assign new_n45237_ = ~new_n44620_ & ~new_n45236_;
  assign new_n45238_ = \b[46]  & ~new_n44609_;
  assign new_n45239_ = ~new_n44607_ & new_n45238_;
  assign new_n45240_ = ~new_n44611_ & ~new_n45239_;
  assign new_n45241_ = ~new_n45237_ & new_n45240_;
  assign new_n45242_ = ~new_n44611_ & ~new_n45241_;
  assign new_n45243_ = \b[47]  & ~new_n44589_;
  assign new_n45244_ = ~new_n44587_ & new_n45243_;
  assign new_n45245_ = ~new_n44602_ & ~new_n45244_;
  assign new_n45246_ = ~new_n45242_ & new_n45245_;
  assign new_n45247_ = ~new_n44602_ & ~new_n45246_;
  assign new_n45248_ = \b[48]  & ~new_n44599_;
  assign new_n45249_ = ~new_n44597_ & new_n45248_;
  assign new_n45250_ = ~new_n44601_ & ~new_n45249_;
  assign new_n45251_ = ~new_n45247_ & new_n45250_;
  assign new_n45252_ = ~new_n44601_ & ~new_n45251_;
  assign new_n45253_ = new_n408_ & ~new_n45252_;
  assign new_n45254_ = ~new_n44590_ & ~new_n45253_;
  assign new_n45255_ = ~new_n44611_ & new_n45245_;
  assign new_n45256_ = ~new_n45241_ & new_n45255_;
  assign new_n45257_ = ~new_n45242_ & ~new_n45245_;
  assign new_n45258_ = ~new_n45256_ & ~new_n45257_;
  assign new_n45259_ = new_n408_ & ~new_n45258_;
  assign new_n45260_ = ~new_n45252_ & new_n45259_;
  assign new_n45261_ = ~new_n45254_ & ~new_n45260_;
  assign new_n45262_ = ~\b[48]  & ~new_n45261_;
  assign new_n45263_ = ~new_n44610_ & ~new_n45253_;
  assign new_n45264_ = ~new_n44620_ & new_n45240_;
  assign new_n45265_ = ~new_n45236_ & new_n45264_;
  assign new_n45266_ = ~new_n45237_ & ~new_n45240_;
  assign new_n45267_ = ~new_n45265_ & ~new_n45266_;
  assign new_n45268_ = new_n408_ & ~new_n45267_;
  assign new_n45269_ = ~new_n45252_ & new_n45268_;
  assign new_n45270_ = ~new_n45263_ & ~new_n45269_;
  assign new_n45271_ = ~\b[47]  & ~new_n45270_;
  assign new_n45272_ = ~new_n44619_ & ~new_n45253_;
  assign new_n45273_ = ~new_n44629_ & new_n45235_;
  assign new_n45274_ = ~new_n45231_ & new_n45273_;
  assign new_n45275_ = ~new_n45232_ & ~new_n45235_;
  assign new_n45276_ = ~new_n45274_ & ~new_n45275_;
  assign new_n45277_ = new_n408_ & ~new_n45276_;
  assign new_n45278_ = ~new_n45252_ & new_n45277_;
  assign new_n45279_ = ~new_n45272_ & ~new_n45278_;
  assign new_n45280_ = ~\b[46]  & ~new_n45279_;
  assign new_n45281_ = ~new_n44628_ & ~new_n45253_;
  assign new_n45282_ = ~new_n44638_ & new_n45230_;
  assign new_n45283_ = ~new_n45226_ & new_n45282_;
  assign new_n45284_ = ~new_n45227_ & ~new_n45230_;
  assign new_n45285_ = ~new_n45283_ & ~new_n45284_;
  assign new_n45286_ = new_n408_ & ~new_n45285_;
  assign new_n45287_ = ~new_n45252_ & new_n45286_;
  assign new_n45288_ = ~new_n45281_ & ~new_n45287_;
  assign new_n45289_ = ~\b[45]  & ~new_n45288_;
  assign new_n45290_ = ~new_n44637_ & ~new_n45253_;
  assign new_n45291_ = ~new_n44647_ & new_n45225_;
  assign new_n45292_ = ~new_n45221_ & new_n45291_;
  assign new_n45293_ = ~new_n45222_ & ~new_n45225_;
  assign new_n45294_ = ~new_n45292_ & ~new_n45293_;
  assign new_n45295_ = new_n408_ & ~new_n45294_;
  assign new_n45296_ = ~new_n45252_ & new_n45295_;
  assign new_n45297_ = ~new_n45290_ & ~new_n45296_;
  assign new_n45298_ = ~\b[44]  & ~new_n45297_;
  assign new_n45299_ = ~new_n44646_ & ~new_n45253_;
  assign new_n45300_ = ~new_n44656_ & new_n45220_;
  assign new_n45301_ = ~new_n45216_ & new_n45300_;
  assign new_n45302_ = ~new_n45217_ & ~new_n45220_;
  assign new_n45303_ = ~new_n45301_ & ~new_n45302_;
  assign new_n45304_ = new_n408_ & ~new_n45303_;
  assign new_n45305_ = ~new_n45252_ & new_n45304_;
  assign new_n45306_ = ~new_n45299_ & ~new_n45305_;
  assign new_n45307_ = ~\b[43]  & ~new_n45306_;
  assign new_n45308_ = ~new_n44655_ & ~new_n45253_;
  assign new_n45309_ = ~new_n44665_ & new_n45215_;
  assign new_n45310_ = ~new_n45211_ & new_n45309_;
  assign new_n45311_ = ~new_n45212_ & ~new_n45215_;
  assign new_n45312_ = ~new_n45310_ & ~new_n45311_;
  assign new_n45313_ = new_n408_ & ~new_n45312_;
  assign new_n45314_ = ~new_n45252_ & new_n45313_;
  assign new_n45315_ = ~new_n45308_ & ~new_n45314_;
  assign new_n45316_ = ~\b[42]  & ~new_n45315_;
  assign new_n45317_ = ~new_n44664_ & ~new_n45253_;
  assign new_n45318_ = ~new_n44674_ & new_n45210_;
  assign new_n45319_ = ~new_n45206_ & new_n45318_;
  assign new_n45320_ = ~new_n45207_ & ~new_n45210_;
  assign new_n45321_ = ~new_n45319_ & ~new_n45320_;
  assign new_n45322_ = new_n408_ & ~new_n45321_;
  assign new_n45323_ = ~new_n45252_ & new_n45322_;
  assign new_n45324_ = ~new_n45317_ & ~new_n45323_;
  assign new_n45325_ = ~\b[41]  & ~new_n45324_;
  assign new_n45326_ = ~new_n44673_ & ~new_n45253_;
  assign new_n45327_ = ~new_n44683_ & new_n45205_;
  assign new_n45328_ = ~new_n45201_ & new_n45327_;
  assign new_n45329_ = ~new_n45202_ & ~new_n45205_;
  assign new_n45330_ = ~new_n45328_ & ~new_n45329_;
  assign new_n45331_ = new_n408_ & ~new_n45330_;
  assign new_n45332_ = ~new_n45252_ & new_n45331_;
  assign new_n45333_ = ~new_n45326_ & ~new_n45332_;
  assign new_n45334_ = ~\b[40]  & ~new_n45333_;
  assign new_n45335_ = ~new_n44682_ & ~new_n45253_;
  assign new_n45336_ = ~new_n44692_ & new_n45200_;
  assign new_n45337_ = ~new_n45196_ & new_n45336_;
  assign new_n45338_ = ~new_n45197_ & ~new_n45200_;
  assign new_n45339_ = ~new_n45337_ & ~new_n45338_;
  assign new_n45340_ = new_n408_ & ~new_n45339_;
  assign new_n45341_ = ~new_n45252_ & new_n45340_;
  assign new_n45342_ = ~new_n45335_ & ~new_n45341_;
  assign new_n45343_ = ~\b[39]  & ~new_n45342_;
  assign new_n45344_ = ~new_n44691_ & ~new_n45253_;
  assign new_n45345_ = ~new_n44701_ & new_n45195_;
  assign new_n45346_ = ~new_n45191_ & new_n45345_;
  assign new_n45347_ = ~new_n45192_ & ~new_n45195_;
  assign new_n45348_ = ~new_n45346_ & ~new_n45347_;
  assign new_n45349_ = new_n408_ & ~new_n45348_;
  assign new_n45350_ = ~new_n45252_ & new_n45349_;
  assign new_n45351_ = ~new_n45344_ & ~new_n45350_;
  assign new_n45352_ = ~\b[38]  & ~new_n45351_;
  assign new_n45353_ = ~new_n44700_ & ~new_n45253_;
  assign new_n45354_ = ~new_n44710_ & new_n45190_;
  assign new_n45355_ = ~new_n45186_ & new_n45354_;
  assign new_n45356_ = ~new_n45187_ & ~new_n45190_;
  assign new_n45357_ = ~new_n45355_ & ~new_n45356_;
  assign new_n45358_ = new_n408_ & ~new_n45357_;
  assign new_n45359_ = ~new_n45252_ & new_n45358_;
  assign new_n45360_ = ~new_n45353_ & ~new_n45359_;
  assign new_n45361_ = ~\b[37]  & ~new_n45360_;
  assign new_n45362_ = ~new_n44709_ & ~new_n45253_;
  assign new_n45363_ = ~new_n44719_ & new_n45185_;
  assign new_n45364_ = ~new_n45181_ & new_n45363_;
  assign new_n45365_ = ~new_n45182_ & ~new_n45185_;
  assign new_n45366_ = ~new_n45364_ & ~new_n45365_;
  assign new_n45367_ = new_n408_ & ~new_n45366_;
  assign new_n45368_ = ~new_n45252_ & new_n45367_;
  assign new_n45369_ = ~new_n45362_ & ~new_n45368_;
  assign new_n45370_ = ~\b[36]  & ~new_n45369_;
  assign new_n45371_ = ~new_n44718_ & ~new_n45253_;
  assign new_n45372_ = ~new_n44728_ & new_n45180_;
  assign new_n45373_ = ~new_n45176_ & new_n45372_;
  assign new_n45374_ = ~new_n45177_ & ~new_n45180_;
  assign new_n45375_ = ~new_n45373_ & ~new_n45374_;
  assign new_n45376_ = new_n408_ & ~new_n45375_;
  assign new_n45377_ = ~new_n45252_ & new_n45376_;
  assign new_n45378_ = ~new_n45371_ & ~new_n45377_;
  assign new_n45379_ = ~\b[35]  & ~new_n45378_;
  assign new_n45380_ = ~new_n44727_ & ~new_n45253_;
  assign new_n45381_ = ~new_n44737_ & new_n45175_;
  assign new_n45382_ = ~new_n45171_ & new_n45381_;
  assign new_n45383_ = ~new_n45172_ & ~new_n45175_;
  assign new_n45384_ = ~new_n45382_ & ~new_n45383_;
  assign new_n45385_ = new_n408_ & ~new_n45384_;
  assign new_n45386_ = ~new_n45252_ & new_n45385_;
  assign new_n45387_ = ~new_n45380_ & ~new_n45386_;
  assign new_n45388_ = ~\b[34]  & ~new_n45387_;
  assign new_n45389_ = ~new_n44736_ & ~new_n45253_;
  assign new_n45390_ = ~new_n44746_ & new_n45170_;
  assign new_n45391_ = ~new_n45166_ & new_n45390_;
  assign new_n45392_ = ~new_n45167_ & ~new_n45170_;
  assign new_n45393_ = ~new_n45391_ & ~new_n45392_;
  assign new_n45394_ = new_n408_ & ~new_n45393_;
  assign new_n45395_ = ~new_n45252_ & new_n45394_;
  assign new_n45396_ = ~new_n45389_ & ~new_n45395_;
  assign new_n45397_ = ~\b[33]  & ~new_n45396_;
  assign new_n45398_ = ~new_n44745_ & ~new_n45253_;
  assign new_n45399_ = ~new_n44755_ & new_n45165_;
  assign new_n45400_ = ~new_n45161_ & new_n45399_;
  assign new_n45401_ = ~new_n45162_ & ~new_n45165_;
  assign new_n45402_ = ~new_n45400_ & ~new_n45401_;
  assign new_n45403_ = new_n408_ & ~new_n45402_;
  assign new_n45404_ = ~new_n45252_ & new_n45403_;
  assign new_n45405_ = ~new_n45398_ & ~new_n45404_;
  assign new_n45406_ = ~\b[32]  & ~new_n45405_;
  assign new_n45407_ = ~new_n44754_ & ~new_n45253_;
  assign new_n45408_ = ~new_n44764_ & new_n45160_;
  assign new_n45409_ = ~new_n45156_ & new_n45408_;
  assign new_n45410_ = ~new_n45157_ & ~new_n45160_;
  assign new_n45411_ = ~new_n45409_ & ~new_n45410_;
  assign new_n45412_ = new_n408_ & ~new_n45411_;
  assign new_n45413_ = ~new_n45252_ & new_n45412_;
  assign new_n45414_ = ~new_n45407_ & ~new_n45413_;
  assign new_n45415_ = ~\b[31]  & ~new_n45414_;
  assign new_n45416_ = ~new_n44763_ & ~new_n45253_;
  assign new_n45417_ = ~new_n44773_ & new_n45155_;
  assign new_n45418_ = ~new_n45151_ & new_n45417_;
  assign new_n45419_ = ~new_n45152_ & ~new_n45155_;
  assign new_n45420_ = ~new_n45418_ & ~new_n45419_;
  assign new_n45421_ = new_n408_ & ~new_n45420_;
  assign new_n45422_ = ~new_n45252_ & new_n45421_;
  assign new_n45423_ = ~new_n45416_ & ~new_n45422_;
  assign new_n45424_ = ~\b[30]  & ~new_n45423_;
  assign new_n45425_ = ~new_n44772_ & ~new_n45253_;
  assign new_n45426_ = ~new_n44782_ & new_n45150_;
  assign new_n45427_ = ~new_n45146_ & new_n45426_;
  assign new_n45428_ = ~new_n45147_ & ~new_n45150_;
  assign new_n45429_ = ~new_n45427_ & ~new_n45428_;
  assign new_n45430_ = new_n408_ & ~new_n45429_;
  assign new_n45431_ = ~new_n45252_ & new_n45430_;
  assign new_n45432_ = ~new_n45425_ & ~new_n45431_;
  assign new_n45433_ = ~\b[29]  & ~new_n45432_;
  assign new_n45434_ = ~new_n44781_ & ~new_n45253_;
  assign new_n45435_ = ~new_n44791_ & new_n45145_;
  assign new_n45436_ = ~new_n45141_ & new_n45435_;
  assign new_n45437_ = ~new_n45142_ & ~new_n45145_;
  assign new_n45438_ = ~new_n45436_ & ~new_n45437_;
  assign new_n45439_ = new_n408_ & ~new_n45438_;
  assign new_n45440_ = ~new_n45252_ & new_n45439_;
  assign new_n45441_ = ~new_n45434_ & ~new_n45440_;
  assign new_n45442_ = ~\b[28]  & ~new_n45441_;
  assign new_n45443_ = ~new_n44790_ & ~new_n45253_;
  assign new_n45444_ = ~new_n44800_ & new_n45140_;
  assign new_n45445_ = ~new_n45136_ & new_n45444_;
  assign new_n45446_ = ~new_n45137_ & ~new_n45140_;
  assign new_n45447_ = ~new_n45445_ & ~new_n45446_;
  assign new_n45448_ = new_n408_ & ~new_n45447_;
  assign new_n45449_ = ~new_n45252_ & new_n45448_;
  assign new_n45450_ = ~new_n45443_ & ~new_n45449_;
  assign new_n45451_ = ~\b[27]  & ~new_n45450_;
  assign new_n45452_ = ~new_n44799_ & ~new_n45253_;
  assign new_n45453_ = ~new_n44809_ & new_n45135_;
  assign new_n45454_ = ~new_n45131_ & new_n45453_;
  assign new_n45455_ = ~new_n45132_ & ~new_n45135_;
  assign new_n45456_ = ~new_n45454_ & ~new_n45455_;
  assign new_n45457_ = new_n408_ & ~new_n45456_;
  assign new_n45458_ = ~new_n45252_ & new_n45457_;
  assign new_n45459_ = ~new_n45452_ & ~new_n45458_;
  assign new_n45460_ = ~\b[26]  & ~new_n45459_;
  assign new_n45461_ = ~new_n44808_ & ~new_n45253_;
  assign new_n45462_ = ~new_n44818_ & new_n45130_;
  assign new_n45463_ = ~new_n45126_ & new_n45462_;
  assign new_n45464_ = ~new_n45127_ & ~new_n45130_;
  assign new_n45465_ = ~new_n45463_ & ~new_n45464_;
  assign new_n45466_ = new_n408_ & ~new_n45465_;
  assign new_n45467_ = ~new_n45252_ & new_n45466_;
  assign new_n45468_ = ~new_n45461_ & ~new_n45467_;
  assign new_n45469_ = ~\b[25]  & ~new_n45468_;
  assign new_n45470_ = ~new_n44817_ & ~new_n45253_;
  assign new_n45471_ = ~new_n44827_ & new_n45125_;
  assign new_n45472_ = ~new_n45121_ & new_n45471_;
  assign new_n45473_ = ~new_n45122_ & ~new_n45125_;
  assign new_n45474_ = ~new_n45472_ & ~new_n45473_;
  assign new_n45475_ = new_n408_ & ~new_n45474_;
  assign new_n45476_ = ~new_n45252_ & new_n45475_;
  assign new_n45477_ = ~new_n45470_ & ~new_n45476_;
  assign new_n45478_ = ~\b[24]  & ~new_n45477_;
  assign new_n45479_ = ~new_n44826_ & ~new_n45253_;
  assign new_n45480_ = ~new_n44836_ & new_n45120_;
  assign new_n45481_ = ~new_n45116_ & new_n45480_;
  assign new_n45482_ = ~new_n45117_ & ~new_n45120_;
  assign new_n45483_ = ~new_n45481_ & ~new_n45482_;
  assign new_n45484_ = new_n408_ & ~new_n45483_;
  assign new_n45485_ = ~new_n45252_ & new_n45484_;
  assign new_n45486_ = ~new_n45479_ & ~new_n45485_;
  assign new_n45487_ = ~\b[23]  & ~new_n45486_;
  assign new_n45488_ = ~new_n44835_ & ~new_n45253_;
  assign new_n45489_ = ~new_n44845_ & new_n45115_;
  assign new_n45490_ = ~new_n45111_ & new_n45489_;
  assign new_n45491_ = ~new_n45112_ & ~new_n45115_;
  assign new_n45492_ = ~new_n45490_ & ~new_n45491_;
  assign new_n45493_ = new_n408_ & ~new_n45492_;
  assign new_n45494_ = ~new_n45252_ & new_n45493_;
  assign new_n45495_ = ~new_n45488_ & ~new_n45494_;
  assign new_n45496_ = ~\b[22]  & ~new_n45495_;
  assign new_n45497_ = ~new_n44844_ & ~new_n45253_;
  assign new_n45498_ = ~new_n44854_ & new_n45110_;
  assign new_n45499_ = ~new_n45106_ & new_n45498_;
  assign new_n45500_ = ~new_n45107_ & ~new_n45110_;
  assign new_n45501_ = ~new_n45499_ & ~new_n45500_;
  assign new_n45502_ = new_n408_ & ~new_n45501_;
  assign new_n45503_ = ~new_n45252_ & new_n45502_;
  assign new_n45504_ = ~new_n45497_ & ~new_n45503_;
  assign new_n45505_ = ~\b[21]  & ~new_n45504_;
  assign new_n45506_ = ~new_n44853_ & ~new_n45253_;
  assign new_n45507_ = ~new_n44863_ & new_n45105_;
  assign new_n45508_ = ~new_n45101_ & new_n45507_;
  assign new_n45509_ = ~new_n45102_ & ~new_n45105_;
  assign new_n45510_ = ~new_n45508_ & ~new_n45509_;
  assign new_n45511_ = new_n408_ & ~new_n45510_;
  assign new_n45512_ = ~new_n45252_ & new_n45511_;
  assign new_n45513_ = ~new_n45506_ & ~new_n45512_;
  assign new_n45514_ = ~\b[20]  & ~new_n45513_;
  assign new_n45515_ = ~new_n44862_ & ~new_n45253_;
  assign new_n45516_ = ~new_n44872_ & new_n45100_;
  assign new_n45517_ = ~new_n45096_ & new_n45516_;
  assign new_n45518_ = ~new_n45097_ & ~new_n45100_;
  assign new_n45519_ = ~new_n45517_ & ~new_n45518_;
  assign new_n45520_ = new_n408_ & ~new_n45519_;
  assign new_n45521_ = ~new_n45252_ & new_n45520_;
  assign new_n45522_ = ~new_n45515_ & ~new_n45521_;
  assign new_n45523_ = ~\b[19]  & ~new_n45522_;
  assign new_n45524_ = ~new_n44871_ & ~new_n45253_;
  assign new_n45525_ = ~new_n44881_ & new_n45095_;
  assign new_n45526_ = ~new_n45091_ & new_n45525_;
  assign new_n45527_ = ~new_n45092_ & ~new_n45095_;
  assign new_n45528_ = ~new_n45526_ & ~new_n45527_;
  assign new_n45529_ = new_n408_ & ~new_n45528_;
  assign new_n45530_ = ~new_n45252_ & new_n45529_;
  assign new_n45531_ = ~new_n45524_ & ~new_n45530_;
  assign new_n45532_ = ~\b[18]  & ~new_n45531_;
  assign new_n45533_ = ~new_n44880_ & ~new_n45253_;
  assign new_n45534_ = ~new_n44890_ & new_n45090_;
  assign new_n45535_ = ~new_n45086_ & new_n45534_;
  assign new_n45536_ = ~new_n45087_ & ~new_n45090_;
  assign new_n45537_ = ~new_n45535_ & ~new_n45536_;
  assign new_n45538_ = new_n408_ & ~new_n45537_;
  assign new_n45539_ = ~new_n45252_ & new_n45538_;
  assign new_n45540_ = ~new_n45533_ & ~new_n45539_;
  assign new_n45541_ = ~\b[17]  & ~new_n45540_;
  assign new_n45542_ = ~new_n44889_ & ~new_n45253_;
  assign new_n45543_ = ~new_n44899_ & new_n45085_;
  assign new_n45544_ = ~new_n45081_ & new_n45543_;
  assign new_n45545_ = ~new_n45082_ & ~new_n45085_;
  assign new_n45546_ = ~new_n45544_ & ~new_n45545_;
  assign new_n45547_ = new_n408_ & ~new_n45546_;
  assign new_n45548_ = ~new_n45252_ & new_n45547_;
  assign new_n45549_ = ~new_n45542_ & ~new_n45548_;
  assign new_n45550_ = ~\b[16]  & ~new_n45549_;
  assign new_n45551_ = ~new_n44898_ & ~new_n45253_;
  assign new_n45552_ = ~new_n44908_ & new_n45080_;
  assign new_n45553_ = ~new_n45076_ & new_n45552_;
  assign new_n45554_ = ~new_n45077_ & ~new_n45080_;
  assign new_n45555_ = ~new_n45553_ & ~new_n45554_;
  assign new_n45556_ = new_n408_ & ~new_n45555_;
  assign new_n45557_ = ~new_n45252_ & new_n45556_;
  assign new_n45558_ = ~new_n45551_ & ~new_n45557_;
  assign new_n45559_ = ~\b[15]  & ~new_n45558_;
  assign new_n45560_ = ~new_n44907_ & ~new_n45253_;
  assign new_n45561_ = ~new_n44917_ & new_n45075_;
  assign new_n45562_ = ~new_n45071_ & new_n45561_;
  assign new_n45563_ = ~new_n45072_ & ~new_n45075_;
  assign new_n45564_ = ~new_n45562_ & ~new_n45563_;
  assign new_n45565_ = new_n408_ & ~new_n45564_;
  assign new_n45566_ = ~new_n45252_ & new_n45565_;
  assign new_n45567_ = ~new_n45560_ & ~new_n45566_;
  assign new_n45568_ = ~\b[14]  & ~new_n45567_;
  assign new_n45569_ = ~new_n44916_ & ~new_n45253_;
  assign new_n45570_ = ~new_n44926_ & new_n45070_;
  assign new_n45571_ = ~new_n45066_ & new_n45570_;
  assign new_n45572_ = ~new_n45067_ & ~new_n45070_;
  assign new_n45573_ = ~new_n45571_ & ~new_n45572_;
  assign new_n45574_ = new_n408_ & ~new_n45573_;
  assign new_n45575_ = ~new_n45252_ & new_n45574_;
  assign new_n45576_ = ~new_n45569_ & ~new_n45575_;
  assign new_n45577_ = ~\b[13]  & ~new_n45576_;
  assign new_n45578_ = ~new_n44925_ & ~new_n45253_;
  assign new_n45579_ = ~new_n44935_ & new_n45065_;
  assign new_n45580_ = ~new_n45061_ & new_n45579_;
  assign new_n45581_ = ~new_n45062_ & ~new_n45065_;
  assign new_n45582_ = ~new_n45580_ & ~new_n45581_;
  assign new_n45583_ = new_n408_ & ~new_n45582_;
  assign new_n45584_ = ~new_n45252_ & new_n45583_;
  assign new_n45585_ = ~new_n45578_ & ~new_n45584_;
  assign new_n45586_ = ~\b[12]  & ~new_n45585_;
  assign new_n45587_ = ~new_n44934_ & ~new_n45253_;
  assign new_n45588_ = ~new_n44944_ & new_n45060_;
  assign new_n45589_ = ~new_n45056_ & new_n45588_;
  assign new_n45590_ = ~new_n45057_ & ~new_n45060_;
  assign new_n45591_ = ~new_n45589_ & ~new_n45590_;
  assign new_n45592_ = new_n408_ & ~new_n45591_;
  assign new_n45593_ = ~new_n45252_ & new_n45592_;
  assign new_n45594_ = ~new_n45587_ & ~new_n45593_;
  assign new_n45595_ = ~\b[11]  & ~new_n45594_;
  assign new_n45596_ = ~new_n44943_ & ~new_n45253_;
  assign new_n45597_ = ~new_n44953_ & new_n45055_;
  assign new_n45598_ = ~new_n45051_ & new_n45597_;
  assign new_n45599_ = ~new_n45052_ & ~new_n45055_;
  assign new_n45600_ = ~new_n45598_ & ~new_n45599_;
  assign new_n45601_ = new_n408_ & ~new_n45600_;
  assign new_n45602_ = ~new_n45252_ & new_n45601_;
  assign new_n45603_ = ~new_n45596_ & ~new_n45602_;
  assign new_n45604_ = ~\b[10]  & ~new_n45603_;
  assign new_n45605_ = ~new_n44952_ & ~new_n45253_;
  assign new_n45606_ = ~new_n44962_ & new_n45050_;
  assign new_n45607_ = ~new_n45046_ & new_n45606_;
  assign new_n45608_ = ~new_n45047_ & ~new_n45050_;
  assign new_n45609_ = ~new_n45607_ & ~new_n45608_;
  assign new_n45610_ = new_n408_ & ~new_n45609_;
  assign new_n45611_ = ~new_n45252_ & new_n45610_;
  assign new_n45612_ = ~new_n45605_ & ~new_n45611_;
  assign new_n45613_ = ~\b[9]  & ~new_n45612_;
  assign new_n45614_ = ~new_n44961_ & ~new_n45253_;
  assign new_n45615_ = ~new_n44971_ & new_n45045_;
  assign new_n45616_ = ~new_n45041_ & new_n45615_;
  assign new_n45617_ = ~new_n45042_ & ~new_n45045_;
  assign new_n45618_ = ~new_n45616_ & ~new_n45617_;
  assign new_n45619_ = new_n408_ & ~new_n45618_;
  assign new_n45620_ = ~new_n45252_ & new_n45619_;
  assign new_n45621_ = ~new_n45614_ & ~new_n45620_;
  assign new_n45622_ = ~\b[8]  & ~new_n45621_;
  assign new_n45623_ = ~new_n44970_ & ~new_n45253_;
  assign new_n45624_ = ~new_n44980_ & new_n45040_;
  assign new_n45625_ = ~new_n45036_ & new_n45624_;
  assign new_n45626_ = ~new_n45037_ & ~new_n45040_;
  assign new_n45627_ = ~new_n45625_ & ~new_n45626_;
  assign new_n45628_ = new_n408_ & ~new_n45627_;
  assign new_n45629_ = ~new_n45252_ & new_n45628_;
  assign new_n45630_ = ~new_n45623_ & ~new_n45629_;
  assign new_n45631_ = ~\b[7]  & ~new_n45630_;
  assign new_n45632_ = ~new_n44979_ & ~new_n45253_;
  assign new_n45633_ = ~new_n44989_ & new_n45035_;
  assign new_n45634_ = ~new_n45031_ & new_n45633_;
  assign new_n45635_ = ~new_n45032_ & ~new_n45035_;
  assign new_n45636_ = ~new_n45634_ & ~new_n45635_;
  assign new_n45637_ = new_n408_ & ~new_n45636_;
  assign new_n45638_ = ~new_n45252_ & new_n45637_;
  assign new_n45639_ = ~new_n45632_ & ~new_n45638_;
  assign new_n45640_ = ~\b[6]  & ~new_n45639_;
  assign new_n45641_ = ~new_n44988_ & ~new_n45253_;
  assign new_n45642_ = ~new_n44998_ & new_n45030_;
  assign new_n45643_ = ~new_n45026_ & new_n45642_;
  assign new_n45644_ = ~new_n45027_ & ~new_n45030_;
  assign new_n45645_ = ~new_n45643_ & ~new_n45644_;
  assign new_n45646_ = new_n408_ & ~new_n45645_;
  assign new_n45647_ = ~new_n45252_ & new_n45646_;
  assign new_n45648_ = ~new_n45641_ & ~new_n45647_;
  assign new_n45649_ = ~\b[5]  & ~new_n45648_;
  assign new_n45650_ = ~new_n44997_ & ~new_n45253_;
  assign new_n45651_ = ~new_n45006_ & new_n45025_;
  assign new_n45652_ = ~new_n45021_ & new_n45651_;
  assign new_n45653_ = ~new_n45022_ & ~new_n45025_;
  assign new_n45654_ = ~new_n45652_ & ~new_n45653_;
  assign new_n45655_ = new_n408_ & ~new_n45654_;
  assign new_n45656_ = ~new_n45252_ & new_n45655_;
  assign new_n45657_ = ~new_n45650_ & ~new_n45656_;
  assign new_n45658_ = ~\b[4]  & ~new_n45657_;
  assign new_n45659_ = ~new_n45005_ & ~new_n45253_;
  assign new_n45660_ = ~new_n45016_ & new_n45020_;
  assign new_n45661_ = ~new_n45015_ & new_n45660_;
  assign new_n45662_ = ~new_n45017_ & ~new_n45020_;
  assign new_n45663_ = ~new_n45661_ & ~new_n45662_;
  assign new_n45664_ = new_n408_ & ~new_n45663_;
  assign new_n45665_ = ~new_n45252_ & new_n45664_;
  assign new_n45666_ = ~new_n45659_ & ~new_n45665_;
  assign new_n45667_ = ~\b[3]  & ~new_n45666_;
  assign new_n45668_ = ~new_n45010_ & ~new_n45253_;
  assign new_n45669_ = new_n16956_ & ~new_n45013_;
  assign new_n45670_ = ~new_n45011_ & new_n45669_;
  assign new_n45671_ = new_n408_ & ~new_n45670_;
  assign new_n45672_ = ~new_n45015_ & new_n45671_;
  assign new_n45673_ = ~new_n45252_ & new_n45672_;
  assign new_n45674_ = ~new_n45668_ & ~new_n45673_;
  assign new_n45675_ = ~\b[2]  & ~new_n45674_;
  assign new_n45676_ = new_n17621_ & ~new_n45252_;
  assign new_n45677_ = \a[15]  & ~new_n45676_;
  assign new_n45678_ = new_n17625_ & ~new_n45252_;
  assign new_n45679_ = ~new_n45677_ & ~new_n45678_;
  assign new_n45680_ = \b[1]  & ~new_n45679_;
  assign new_n45681_ = ~\b[1]  & ~new_n45678_;
  assign new_n45682_ = ~new_n45677_ & new_n45681_;
  assign new_n45683_ = ~new_n45680_ & ~new_n45682_;
  assign new_n45684_ = ~new_n17632_ & ~new_n45683_;
  assign new_n45685_ = ~\b[1]  & ~new_n45679_;
  assign new_n45686_ = ~new_n45684_ & ~new_n45685_;
  assign new_n45687_ = \b[2]  & ~new_n45673_;
  assign new_n45688_ = ~new_n45668_ & new_n45687_;
  assign new_n45689_ = ~new_n45675_ & ~new_n45688_;
  assign new_n45690_ = ~new_n45686_ & new_n45689_;
  assign new_n45691_ = ~new_n45675_ & ~new_n45690_;
  assign new_n45692_ = \b[3]  & ~new_n45665_;
  assign new_n45693_ = ~new_n45659_ & new_n45692_;
  assign new_n45694_ = ~new_n45667_ & ~new_n45693_;
  assign new_n45695_ = ~new_n45691_ & new_n45694_;
  assign new_n45696_ = ~new_n45667_ & ~new_n45695_;
  assign new_n45697_ = \b[4]  & ~new_n45656_;
  assign new_n45698_ = ~new_n45650_ & new_n45697_;
  assign new_n45699_ = ~new_n45658_ & ~new_n45698_;
  assign new_n45700_ = ~new_n45696_ & new_n45699_;
  assign new_n45701_ = ~new_n45658_ & ~new_n45700_;
  assign new_n45702_ = \b[5]  & ~new_n45647_;
  assign new_n45703_ = ~new_n45641_ & new_n45702_;
  assign new_n45704_ = ~new_n45649_ & ~new_n45703_;
  assign new_n45705_ = ~new_n45701_ & new_n45704_;
  assign new_n45706_ = ~new_n45649_ & ~new_n45705_;
  assign new_n45707_ = \b[6]  & ~new_n45638_;
  assign new_n45708_ = ~new_n45632_ & new_n45707_;
  assign new_n45709_ = ~new_n45640_ & ~new_n45708_;
  assign new_n45710_ = ~new_n45706_ & new_n45709_;
  assign new_n45711_ = ~new_n45640_ & ~new_n45710_;
  assign new_n45712_ = \b[7]  & ~new_n45629_;
  assign new_n45713_ = ~new_n45623_ & new_n45712_;
  assign new_n45714_ = ~new_n45631_ & ~new_n45713_;
  assign new_n45715_ = ~new_n45711_ & new_n45714_;
  assign new_n45716_ = ~new_n45631_ & ~new_n45715_;
  assign new_n45717_ = \b[8]  & ~new_n45620_;
  assign new_n45718_ = ~new_n45614_ & new_n45717_;
  assign new_n45719_ = ~new_n45622_ & ~new_n45718_;
  assign new_n45720_ = ~new_n45716_ & new_n45719_;
  assign new_n45721_ = ~new_n45622_ & ~new_n45720_;
  assign new_n45722_ = \b[9]  & ~new_n45611_;
  assign new_n45723_ = ~new_n45605_ & new_n45722_;
  assign new_n45724_ = ~new_n45613_ & ~new_n45723_;
  assign new_n45725_ = ~new_n45721_ & new_n45724_;
  assign new_n45726_ = ~new_n45613_ & ~new_n45725_;
  assign new_n45727_ = \b[10]  & ~new_n45602_;
  assign new_n45728_ = ~new_n45596_ & new_n45727_;
  assign new_n45729_ = ~new_n45604_ & ~new_n45728_;
  assign new_n45730_ = ~new_n45726_ & new_n45729_;
  assign new_n45731_ = ~new_n45604_ & ~new_n45730_;
  assign new_n45732_ = \b[11]  & ~new_n45593_;
  assign new_n45733_ = ~new_n45587_ & new_n45732_;
  assign new_n45734_ = ~new_n45595_ & ~new_n45733_;
  assign new_n45735_ = ~new_n45731_ & new_n45734_;
  assign new_n45736_ = ~new_n45595_ & ~new_n45735_;
  assign new_n45737_ = \b[12]  & ~new_n45584_;
  assign new_n45738_ = ~new_n45578_ & new_n45737_;
  assign new_n45739_ = ~new_n45586_ & ~new_n45738_;
  assign new_n45740_ = ~new_n45736_ & new_n45739_;
  assign new_n45741_ = ~new_n45586_ & ~new_n45740_;
  assign new_n45742_ = \b[13]  & ~new_n45575_;
  assign new_n45743_ = ~new_n45569_ & new_n45742_;
  assign new_n45744_ = ~new_n45577_ & ~new_n45743_;
  assign new_n45745_ = ~new_n45741_ & new_n45744_;
  assign new_n45746_ = ~new_n45577_ & ~new_n45745_;
  assign new_n45747_ = \b[14]  & ~new_n45566_;
  assign new_n45748_ = ~new_n45560_ & new_n45747_;
  assign new_n45749_ = ~new_n45568_ & ~new_n45748_;
  assign new_n45750_ = ~new_n45746_ & new_n45749_;
  assign new_n45751_ = ~new_n45568_ & ~new_n45750_;
  assign new_n45752_ = \b[15]  & ~new_n45557_;
  assign new_n45753_ = ~new_n45551_ & new_n45752_;
  assign new_n45754_ = ~new_n45559_ & ~new_n45753_;
  assign new_n45755_ = ~new_n45751_ & new_n45754_;
  assign new_n45756_ = ~new_n45559_ & ~new_n45755_;
  assign new_n45757_ = \b[16]  & ~new_n45548_;
  assign new_n45758_ = ~new_n45542_ & new_n45757_;
  assign new_n45759_ = ~new_n45550_ & ~new_n45758_;
  assign new_n45760_ = ~new_n45756_ & new_n45759_;
  assign new_n45761_ = ~new_n45550_ & ~new_n45760_;
  assign new_n45762_ = \b[17]  & ~new_n45539_;
  assign new_n45763_ = ~new_n45533_ & new_n45762_;
  assign new_n45764_ = ~new_n45541_ & ~new_n45763_;
  assign new_n45765_ = ~new_n45761_ & new_n45764_;
  assign new_n45766_ = ~new_n45541_ & ~new_n45765_;
  assign new_n45767_ = \b[18]  & ~new_n45530_;
  assign new_n45768_ = ~new_n45524_ & new_n45767_;
  assign new_n45769_ = ~new_n45532_ & ~new_n45768_;
  assign new_n45770_ = ~new_n45766_ & new_n45769_;
  assign new_n45771_ = ~new_n45532_ & ~new_n45770_;
  assign new_n45772_ = \b[19]  & ~new_n45521_;
  assign new_n45773_ = ~new_n45515_ & new_n45772_;
  assign new_n45774_ = ~new_n45523_ & ~new_n45773_;
  assign new_n45775_ = ~new_n45771_ & new_n45774_;
  assign new_n45776_ = ~new_n45523_ & ~new_n45775_;
  assign new_n45777_ = \b[20]  & ~new_n45512_;
  assign new_n45778_ = ~new_n45506_ & new_n45777_;
  assign new_n45779_ = ~new_n45514_ & ~new_n45778_;
  assign new_n45780_ = ~new_n45776_ & new_n45779_;
  assign new_n45781_ = ~new_n45514_ & ~new_n45780_;
  assign new_n45782_ = \b[21]  & ~new_n45503_;
  assign new_n45783_ = ~new_n45497_ & new_n45782_;
  assign new_n45784_ = ~new_n45505_ & ~new_n45783_;
  assign new_n45785_ = ~new_n45781_ & new_n45784_;
  assign new_n45786_ = ~new_n45505_ & ~new_n45785_;
  assign new_n45787_ = \b[22]  & ~new_n45494_;
  assign new_n45788_ = ~new_n45488_ & new_n45787_;
  assign new_n45789_ = ~new_n45496_ & ~new_n45788_;
  assign new_n45790_ = ~new_n45786_ & new_n45789_;
  assign new_n45791_ = ~new_n45496_ & ~new_n45790_;
  assign new_n45792_ = \b[23]  & ~new_n45485_;
  assign new_n45793_ = ~new_n45479_ & new_n45792_;
  assign new_n45794_ = ~new_n45487_ & ~new_n45793_;
  assign new_n45795_ = ~new_n45791_ & new_n45794_;
  assign new_n45796_ = ~new_n45487_ & ~new_n45795_;
  assign new_n45797_ = \b[24]  & ~new_n45476_;
  assign new_n45798_ = ~new_n45470_ & new_n45797_;
  assign new_n45799_ = ~new_n45478_ & ~new_n45798_;
  assign new_n45800_ = ~new_n45796_ & new_n45799_;
  assign new_n45801_ = ~new_n45478_ & ~new_n45800_;
  assign new_n45802_ = \b[25]  & ~new_n45467_;
  assign new_n45803_ = ~new_n45461_ & new_n45802_;
  assign new_n45804_ = ~new_n45469_ & ~new_n45803_;
  assign new_n45805_ = ~new_n45801_ & new_n45804_;
  assign new_n45806_ = ~new_n45469_ & ~new_n45805_;
  assign new_n45807_ = \b[26]  & ~new_n45458_;
  assign new_n45808_ = ~new_n45452_ & new_n45807_;
  assign new_n45809_ = ~new_n45460_ & ~new_n45808_;
  assign new_n45810_ = ~new_n45806_ & new_n45809_;
  assign new_n45811_ = ~new_n45460_ & ~new_n45810_;
  assign new_n45812_ = \b[27]  & ~new_n45449_;
  assign new_n45813_ = ~new_n45443_ & new_n45812_;
  assign new_n45814_ = ~new_n45451_ & ~new_n45813_;
  assign new_n45815_ = ~new_n45811_ & new_n45814_;
  assign new_n45816_ = ~new_n45451_ & ~new_n45815_;
  assign new_n45817_ = \b[28]  & ~new_n45440_;
  assign new_n45818_ = ~new_n45434_ & new_n45817_;
  assign new_n45819_ = ~new_n45442_ & ~new_n45818_;
  assign new_n45820_ = ~new_n45816_ & new_n45819_;
  assign new_n45821_ = ~new_n45442_ & ~new_n45820_;
  assign new_n45822_ = \b[29]  & ~new_n45431_;
  assign new_n45823_ = ~new_n45425_ & new_n45822_;
  assign new_n45824_ = ~new_n45433_ & ~new_n45823_;
  assign new_n45825_ = ~new_n45821_ & new_n45824_;
  assign new_n45826_ = ~new_n45433_ & ~new_n45825_;
  assign new_n45827_ = \b[30]  & ~new_n45422_;
  assign new_n45828_ = ~new_n45416_ & new_n45827_;
  assign new_n45829_ = ~new_n45424_ & ~new_n45828_;
  assign new_n45830_ = ~new_n45826_ & new_n45829_;
  assign new_n45831_ = ~new_n45424_ & ~new_n45830_;
  assign new_n45832_ = \b[31]  & ~new_n45413_;
  assign new_n45833_ = ~new_n45407_ & new_n45832_;
  assign new_n45834_ = ~new_n45415_ & ~new_n45833_;
  assign new_n45835_ = ~new_n45831_ & new_n45834_;
  assign new_n45836_ = ~new_n45415_ & ~new_n45835_;
  assign new_n45837_ = \b[32]  & ~new_n45404_;
  assign new_n45838_ = ~new_n45398_ & new_n45837_;
  assign new_n45839_ = ~new_n45406_ & ~new_n45838_;
  assign new_n45840_ = ~new_n45836_ & new_n45839_;
  assign new_n45841_ = ~new_n45406_ & ~new_n45840_;
  assign new_n45842_ = \b[33]  & ~new_n45395_;
  assign new_n45843_ = ~new_n45389_ & new_n45842_;
  assign new_n45844_ = ~new_n45397_ & ~new_n45843_;
  assign new_n45845_ = ~new_n45841_ & new_n45844_;
  assign new_n45846_ = ~new_n45397_ & ~new_n45845_;
  assign new_n45847_ = \b[34]  & ~new_n45386_;
  assign new_n45848_ = ~new_n45380_ & new_n45847_;
  assign new_n45849_ = ~new_n45388_ & ~new_n45848_;
  assign new_n45850_ = ~new_n45846_ & new_n45849_;
  assign new_n45851_ = ~new_n45388_ & ~new_n45850_;
  assign new_n45852_ = \b[35]  & ~new_n45377_;
  assign new_n45853_ = ~new_n45371_ & new_n45852_;
  assign new_n45854_ = ~new_n45379_ & ~new_n45853_;
  assign new_n45855_ = ~new_n45851_ & new_n45854_;
  assign new_n45856_ = ~new_n45379_ & ~new_n45855_;
  assign new_n45857_ = \b[36]  & ~new_n45368_;
  assign new_n45858_ = ~new_n45362_ & new_n45857_;
  assign new_n45859_ = ~new_n45370_ & ~new_n45858_;
  assign new_n45860_ = ~new_n45856_ & new_n45859_;
  assign new_n45861_ = ~new_n45370_ & ~new_n45860_;
  assign new_n45862_ = \b[37]  & ~new_n45359_;
  assign new_n45863_ = ~new_n45353_ & new_n45862_;
  assign new_n45864_ = ~new_n45361_ & ~new_n45863_;
  assign new_n45865_ = ~new_n45861_ & new_n45864_;
  assign new_n45866_ = ~new_n45361_ & ~new_n45865_;
  assign new_n45867_ = \b[38]  & ~new_n45350_;
  assign new_n45868_ = ~new_n45344_ & new_n45867_;
  assign new_n45869_ = ~new_n45352_ & ~new_n45868_;
  assign new_n45870_ = ~new_n45866_ & new_n45869_;
  assign new_n45871_ = ~new_n45352_ & ~new_n45870_;
  assign new_n45872_ = \b[39]  & ~new_n45341_;
  assign new_n45873_ = ~new_n45335_ & new_n45872_;
  assign new_n45874_ = ~new_n45343_ & ~new_n45873_;
  assign new_n45875_ = ~new_n45871_ & new_n45874_;
  assign new_n45876_ = ~new_n45343_ & ~new_n45875_;
  assign new_n45877_ = \b[40]  & ~new_n45332_;
  assign new_n45878_ = ~new_n45326_ & new_n45877_;
  assign new_n45879_ = ~new_n45334_ & ~new_n45878_;
  assign new_n45880_ = ~new_n45876_ & new_n45879_;
  assign new_n45881_ = ~new_n45334_ & ~new_n45880_;
  assign new_n45882_ = \b[41]  & ~new_n45323_;
  assign new_n45883_ = ~new_n45317_ & new_n45882_;
  assign new_n45884_ = ~new_n45325_ & ~new_n45883_;
  assign new_n45885_ = ~new_n45881_ & new_n45884_;
  assign new_n45886_ = ~new_n45325_ & ~new_n45885_;
  assign new_n45887_ = \b[42]  & ~new_n45314_;
  assign new_n45888_ = ~new_n45308_ & new_n45887_;
  assign new_n45889_ = ~new_n45316_ & ~new_n45888_;
  assign new_n45890_ = ~new_n45886_ & new_n45889_;
  assign new_n45891_ = ~new_n45316_ & ~new_n45890_;
  assign new_n45892_ = \b[43]  & ~new_n45305_;
  assign new_n45893_ = ~new_n45299_ & new_n45892_;
  assign new_n45894_ = ~new_n45307_ & ~new_n45893_;
  assign new_n45895_ = ~new_n45891_ & new_n45894_;
  assign new_n45896_ = ~new_n45307_ & ~new_n45895_;
  assign new_n45897_ = \b[44]  & ~new_n45296_;
  assign new_n45898_ = ~new_n45290_ & new_n45897_;
  assign new_n45899_ = ~new_n45298_ & ~new_n45898_;
  assign new_n45900_ = ~new_n45896_ & new_n45899_;
  assign new_n45901_ = ~new_n45298_ & ~new_n45900_;
  assign new_n45902_ = \b[45]  & ~new_n45287_;
  assign new_n45903_ = ~new_n45281_ & new_n45902_;
  assign new_n45904_ = ~new_n45289_ & ~new_n45903_;
  assign new_n45905_ = ~new_n45901_ & new_n45904_;
  assign new_n45906_ = ~new_n45289_ & ~new_n45905_;
  assign new_n45907_ = \b[46]  & ~new_n45278_;
  assign new_n45908_ = ~new_n45272_ & new_n45907_;
  assign new_n45909_ = ~new_n45280_ & ~new_n45908_;
  assign new_n45910_ = ~new_n45906_ & new_n45909_;
  assign new_n45911_ = ~new_n45280_ & ~new_n45910_;
  assign new_n45912_ = \b[47]  & ~new_n45269_;
  assign new_n45913_ = ~new_n45263_ & new_n45912_;
  assign new_n45914_ = ~new_n45271_ & ~new_n45913_;
  assign new_n45915_ = ~new_n45911_ & new_n45914_;
  assign new_n45916_ = ~new_n45271_ & ~new_n45915_;
  assign new_n45917_ = \b[48]  & ~new_n45260_;
  assign new_n45918_ = ~new_n45254_ & new_n45917_;
  assign new_n45919_ = ~new_n45262_ & ~new_n45918_;
  assign new_n45920_ = ~new_n45916_ & new_n45919_;
  assign new_n45921_ = ~new_n45262_ & ~new_n45920_;
  assign new_n45922_ = ~new_n44600_ & ~new_n45253_;
  assign new_n45923_ = ~new_n44602_ & new_n45250_;
  assign new_n45924_ = ~new_n45246_ & new_n45923_;
  assign new_n45925_ = ~new_n45247_ & ~new_n45250_;
  assign new_n45926_ = ~new_n45924_ & ~new_n45925_;
  assign new_n45927_ = new_n45253_ & ~new_n45926_;
  assign new_n45928_ = ~new_n45922_ & ~new_n45927_;
  assign new_n45929_ = ~\b[49]  & ~new_n45928_;
  assign new_n45930_ = \b[49]  & ~new_n45922_;
  assign new_n45931_ = ~new_n45927_ & new_n45930_;
  assign new_n45932_ = new_n17882_ & ~new_n45931_;
  assign new_n45933_ = ~new_n45929_ & new_n45932_;
  assign new_n45934_ = ~new_n45921_ & new_n45933_;
  assign new_n45935_ = new_n408_ & ~new_n45928_;
  assign new_n45936_ = ~new_n45934_ & ~new_n45935_;
  assign new_n45937_ = ~new_n45271_ & new_n45919_;
  assign new_n45938_ = ~new_n45915_ & new_n45937_;
  assign new_n45939_ = ~new_n45916_ & ~new_n45919_;
  assign new_n45940_ = ~new_n45938_ & ~new_n45939_;
  assign new_n45941_ = ~new_n45936_ & ~new_n45940_;
  assign new_n45942_ = ~new_n45261_ & ~new_n45935_;
  assign new_n45943_ = ~new_n45934_ & new_n45942_;
  assign new_n45944_ = ~new_n45941_ & ~new_n45943_;
  assign new_n45945_ = ~\b[49]  & ~new_n45944_;
  assign new_n45946_ = ~new_n45280_ & new_n45914_;
  assign new_n45947_ = ~new_n45910_ & new_n45946_;
  assign new_n45948_ = ~new_n45911_ & ~new_n45914_;
  assign new_n45949_ = ~new_n45947_ & ~new_n45948_;
  assign new_n45950_ = ~new_n45936_ & ~new_n45949_;
  assign new_n45951_ = ~new_n45270_ & ~new_n45935_;
  assign new_n45952_ = ~new_n45934_ & new_n45951_;
  assign new_n45953_ = ~new_n45950_ & ~new_n45952_;
  assign new_n45954_ = ~\b[48]  & ~new_n45953_;
  assign new_n45955_ = ~new_n45289_ & new_n45909_;
  assign new_n45956_ = ~new_n45905_ & new_n45955_;
  assign new_n45957_ = ~new_n45906_ & ~new_n45909_;
  assign new_n45958_ = ~new_n45956_ & ~new_n45957_;
  assign new_n45959_ = ~new_n45936_ & ~new_n45958_;
  assign new_n45960_ = ~new_n45279_ & ~new_n45935_;
  assign new_n45961_ = ~new_n45934_ & new_n45960_;
  assign new_n45962_ = ~new_n45959_ & ~new_n45961_;
  assign new_n45963_ = ~\b[47]  & ~new_n45962_;
  assign new_n45964_ = ~new_n45298_ & new_n45904_;
  assign new_n45965_ = ~new_n45900_ & new_n45964_;
  assign new_n45966_ = ~new_n45901_ & ~new_n45904_;
  assign new_n45967_ = ~new_n45965_ & ~new_n45966_;
  assign new_n45968_ = ~new_n45936_ & ~new_n45967_;
  assign new_n45969_ = ~new_n45288_ & ~new_n45935_;
  assign new_n45970_ = ~new_n45934_ & new_n45969_;
  assign new_n45971_ = ~new_n45968_ & ~new_n45970_;
  assign new_n45972_ = ~\b[46]  & ~new_n45971_;
  assign new_n45973_ = ~new_n45307_ & new_n45899_;
  assign new_n45974_ = ~new_n45895_ & new_n45973_;
  assign new_n45975_ = ~new_n45896_ & ~new_n45899_;
  assign new_n45976_ = ~new_n45974_ & ~new_n45975_;
  assign new_n45977_ = ~new_n45936_ & ~new_n45976_;
  assign new_n45978_ = ~new_n45297_ & ~new_n45935_;
  assign new_n45979_ = ~new_n45934_ & new_n45978_;
  assign new_n45980_ = ~new_n45977_ & ~new_n45979_;
  assign new_n45981_ = ~\b[45]  & ~new_n45980_;
  assign new_n45982_ = ~new_n45316_ & new_n45894_;
  assign new_n45983_ = ~new_n45890_ & new_n45982_;
  assign new_n45984_ = ~new_n45891_ & ~new_n45894_;
  assign new_n45985_ = ~new_n45983_ & ~new_n45984_;
  assign new_n45986_ = ~new_n45936_ & ~new_n45985_;
  assign new_n45987_ = ~new_n45306_ & ~new_n45935_;
  assign new_n45988_ = ~new_n45934_ & new_n45987_;
  assign new_n45989_ = ~new_n45986_ & ~new_n45988_;
  assign new_n45990_ = ~\b[44]  & ~new_n45989_;
  assign new_n45991_ = ~new_n45325_ & new_n45889_;
  assign new_n45992_ = ~new_n45885_ & new_n45991_;
  assign new_n45993_ = ~new_n45886_ & ~new_n45889_;
  assign new_n45994_ = ~new_n45992_ & ~new_n45993_;
  assign new_n45995_ = ~new_n45936_ & ~new_n45994_;
  assign new_n45996_ = ~new_n45315_ & ~new_n45935_;
  assign new_n45997_ = ~new_n45934_ & new_n45996_;
  assign new_n45998_ = ~new_n45995_ & ~new_n45997_;
  assign new_n45999_ = ~\b[43]  & ~new_n45998_;
  assign new_n46000_ = ~new_n45334_ & new_n45884_;
  assign new_n46001_ = ~new_n45880_ & new_n46000_;
  assign new_n46002_ = ~new_n45881_ & ~new_n45884_;
  assign new_n46003_ = ~new_n46001_ & ~new_n46002_;
  assign new_n46004_ = ~new_n45936_ & ~new_n46003_;
  assign new_n46005_ = ~new_n45324_ & ~new_n45935_;
  assign new_n46006_ = ~new_n45934_ & new_n46005_;
  assign new_n46007_ = ~new_n46004_ & ~new_n46006_;
  assign new_n46008_ = ~\b[42]  & ~new_n46007_;
  assign new_n46009_ = ~new_n45343_ & new_n45879_;
  assign new_n46010_ = ~new_n45875_ & new_n46009_;
  assign new_n46011_ = ~new_n45876_ & ~new_n45879_;
  assign new_n46012_ = ~new_n46010_ & ~new_n46011_;
  assign new_n46013_ = ~new_n45936_ & ~new_n46012_;
  assign new_n46014_ = ~new_n45333_ & ~new_n45935_;
  assign new_n46015_ = ~new_n45934_ & new_n46014_;
  assign new_n46016_ = ~new_n46013_ & ~new_n46015_;
  assign new_n46017_ = ~\b[41]  & ~new_n46016_;
  assign new_n46018_ = ~new_n45352_ & new_n45874_;
  assign new_n46019_ = ~new_n45870_ & new_n46018_;
  assign new_n46020_ = ~new_n45871_ & ~new_n45874_;
  assign new_n46021_ = ~new_n46019_ & ~new_n46020_;
  assign new_n46022_ = ~new_n45936_ & ~new_n46021_;
  assign new_n46023_ = ~new_n45342_ & ~new_n45935_;
  assign new_n46024_ = ~new_n45934_ & new_n46023_;
  assign new_n46025_ = ~new_n46022_ & ~new_n46024_;
  assign new_n46026_ = ~\b[40]  & ~new_n46025_;
  assign new_n46027_ = ~new_n45361_ & new_n45869_;
  assign new_n46028_ = ~new_n45865_ & new_n46027_;
  assign new_n46029_ = ~new_n45866_ & ~new_n45869_;
  assign new_n46030_ = ~new_n46028_ & ~new_n46029_;
  assign new_n46031_ = ~new_n45936_ & ~new_n46030_;
  assign new_n46032_ = ~new_n45351_ & ~new_n45935_;
  assign new_n46033_ = ~new_n45934_ & new_n46032_;
  assign new_n46034_ = ~new_n46031_ & ~new_n46033_;
  assign new_n46035_ = ~\b[39]  & ~new_n46034_;
  assign new_n46036_ = ~new_n45370_ & new_n45864_;
  assign new_n46037_ = ~new_n45860_ & new_n46036_;
  assign new_n46038_ = ~new_n45861_ & ~new_n45864_;
  assign new_n46039_ = ~new_n46037_ & ~new_n46038_;
  assign new_n46040_ = ~new_n45936_ & ~new_n46039_;
  assign new_n46041_ = ~new_n45360_ & ~new_n45935_;
  assign new_n46042_ = ~new_n45934_ & new_n46041_;
  assign new_n46043_ = ~new_n46040_ & ~new_n46042_;
  assign new_n46044_ = ~\b[38]  & ~new_n46043_;
  assign new_n46045_ = ~new_n45379_ & new_n45859_;
  assign new_n46046_ = ~new_n45855_ & new_n46045_;
  assign new_n46047_ = ~new_n45856_ & ~new_n45859_;
  assign new_n46048_ = ~new_n46046_ & ~new_n46047_;
  assign new_n46049_ = ~new_n45936_ & ~new_n46048_;
  assign new_n46050_ = ~new_n45369_ & ~new_n45935_;
  assign new_n46051_ = ~new_n45934_ & new_n46050_;
  assign new_n46052_ = ~new_n46049_ & ~new_n46051_;
  assign new_n46053_ = ~\b[37]  & ~new_n46052_;
  assign new_n46054_ = ~new_n45388_ & new_n45854_;
  assign new_n46055_ = ~new_n45850_ & new_n46054_;
  assign new_n46056_ = ~new_n45851_ & ~new_n45854_;
  assign new_n46057_ = ~new_n46055_ & ~new_n46056_;
  assign new_n46058_ = ~new_n45936_ & ~new_n46057_;
  assign new_n46059_ = ~new_n45378_ & ~new_n45935_;
  assign new_n46060_ = ~new_n45934_ & new_n46059_;
  assign new_n46061_ = ~new_n46058_ & ~new_n46060_;
  assign new_n46062_ = ~\b[36]  & ~new_n46061_;
  assign new_n46063_ = ~new_n45397_ & new_n45849_;
  assign new_n46064_ = ~new_n45845_ & new_n46063_;
  assign new_n46065_ = ~new_n45846_ & ~new_n45849_;
  assign new_n46066_ = ~new_n46064_ & ~new_n46065_;
  assign new_n46067_ = ~new_n45936_ & ~new_n46066_;
  assign new_n46068_ = ~new_n45387_ & ~new_n45935_;
  assign new_n46069_ = ~new_n45934_ & new_n46068_;
  assign new_n46070_ = ~new_n46067_ & ~new_n46069_;
  assign new_n46071_ = ~\b[35]  & ~new_n46070_;
  assign new_n46072_ = ~new_n45406_ & new_n45844_;
  assign new_n46073_ = ~new_n45840_ & new_n46072_;
  assign new_n46074_ = ~new_n45841_ & ~new_n45844_;
  assign new_n46075_ = ~new_n46073_ & ~new_n46074_;
  assign new_n46076_ = ~new_n45936_ & ~new_n46075_;
  assign new_n46077_ = ~new_n45396_ & ~new_n45935_;
  assign new_n46078_ = ~new_n45934_ & new_n46077_;
  assign new_n46079_ = ~new_n46076_ & ~new_n46078_;
  assign new_n46080_ = ~\b[34]  & ~new_n46079_;
  assign new_n46081_ = ~new_n45415_ & new_n45839_;
  assign new_n46082_ = ~new_n45835_ & new_n46081_;
  assign new_n46083_ = ~new_n45836_ & ~new_n45839_;
  assign new_n46084_ = ~new_n46082_ & ~new_n46083_;
  assign new_n46085_ = ~new_n45936_ & ~new_n46084_;
  assign new_n46086_ = ~new_n45405_ & ~new_n45935_;
  assign new_n46087_ = ~new_n45934_ & new_n46086_;
  assign new_n46088_ = ~new_n46085_ & ~new_n46087_;
  assign new_n46089_ = ~\b[33]  & ~new_n46088_;
  assign new_n46090_ = ~new_n45424_ & new_n45834_;
  assign new_n46091_ = ~new_n45830_ & new_n46090_;
  assign new_n46092_ = ~new_n45831_ & ~new_n45834_;
  assign new_n46093_ = ~new_n46091_ & ~new_n46092_;
  assign new_n46094_ = ~new_n45936_ & ~new_n46093_;
  assign new_n46095_ = ~new_n45414_ & ~new_n45935_;
  assign new_n46096_ = ~new_n45934_ & new_n46095_;
  assign new_n46097_ = ~new_n46094_ & ~new_n46096_;
  assign new_n46098_ = ~\b[32]  & ~new_n46097_;
  assign new_n46099_ = ~new_n45433_ & new_n45829_;
  assign new_n46100_ = ~new_n45825_ & new_n46099_;
  assign new_n46101_ = ~new_n45826_ & ~new_n45829_;
  assign new_n46102_ = ~new_n46100_ & ~new_n46101_;
  assign new_n46103_ = ~new_n45936_ & ~new_n46102_;
  assign new_n46104_ = ~new_n45423_ & ~new_n45935_;
  assign new_n46105_ = ~new_n45934_ & new_n46104_;
  assign new_n46106_ = ~new_n46103_ & ~new_n46105_;
  assign new_n46107_ = ~\b[31]  & ~new_n46106_;
  assign new_n46108_ = ~new_n45442_ & new_n45824_;
  assign new_n46109_ = ~new_n45820_ & new_n46108_;
  assign new_n46110_ = ~new_n45821_ & ~new_n45824_;
  assign new_n46111_ = ~new_n46109_ & ~new_n46110_;
  assign new_n46112_ = ~new_n45936_ & ~new_n46111_;
  assign new_n46113_ = ~new_n45432_ & ~new_n45935_;
  assign new_n46114_ = ~new_n45934_ & new_n46113_;
  assign new_n46115_ = ~new_n46112_ & ~new_n46114_;
  assign new_n46116_ = ~\b[30]  & ~new_n46115_;
  assign new_n46117_ = ~new_n45451_ & new_n45819_;
  assign new_n46118_ = ~new_n45815_ & new_n46117_;
  assign new_n46119_ = ~new_n45816_ & ~new_n45819_;
  assign new_n46120_ = ~new_n46118_ & ~new_n46119_;
  assign new_n46121_ = ~new_n45936_ & ~new_n46120_;
  assign new_n46122_ = ~new_n45441_ & ~new_n45935_;
  assign new_n46123_ = ~new_n45934_ & new_n46122_;
  assign new_n46124_ = ~new_n46121_ & ~new_n46123_;
  assign new_n46125_ = ~\b[29]  & ~new_n46124_;
  assign new_n46126_ = ~new_n45460_ & new_n45814_;
  assign new_n46127_ = ~new_n45810_ & new_n46126_;
  assign new_n46128_ = ~new_n45811_ & ~new_n45814_;
  assign new_n46129_ = ~new_n46127_ & ~new_n46128_;
  assign new_n46130_ = ~new_n45936_ & ~new_n46129_;
  assign new_n46131_ = ~new_n45450_ & ~new_n45935_;
  assign new_n46132_ = ~new_n45934_ & new_n46131_;
  assign new_n46133_ = ~new_n46130_ & ~new_n46132_;
  assign new_n46134_ = ~\b[28]  & ~new_n46133_;
  assign new_n46135_ = ~new_n45469_ & new_n45809_;
  assign new_n46136_ = ~new_n45805_ & new_n46135_;
  assign new_n46137_ = ~new_n45806_ & ~new_n45809_;
  assign new_n46138_ = ~new_n46136_ & ~new_n46137_;
  assign new_n46139_ = ~new_n45936_ & ~new_n46138_;
  assign new_n46140_ = ~new_n45459_ & ~new_n45935_;
  assign new_n46141_ = ~new_n45934_ & new_n46140_;
  assign new_n46142_ = ~new_n46139_ & ~new_n46141_;
  assign new_n46143_ = ~\b[27]  & ~new_n46142_;
  assign new_n46144_ = ~new_n45478_ & new_n45804_;
  assign new_n46145_ = ~new_n45800_ & new_n46144_;
  assign new_n46146_ = ~new_n45801_ & ~new_n45804_;
  assign new_n46147_ = ~new_n46145_ & ~new_n46146_;
  assign new_n46148_ = ~new_n45936_ & ~new_n46147_;
  assign new_n46149_ = ~new_n45468_ & ~new_n45935_;
  assign new_n46150_ = ~new_n45934_ & new_n46149_;
  assign new_n46151_ = ~new_n46148_ & ~new_n46150_;
  assign new_n46152_ = ~\b[26]  & ~new_n46151_;
  assign new_n46153_ = ~new_n45487_ & new_n45799_;
  assign new_n46154_ = ~new_n45795_ & new_n46153_;
  assign new_n46155_ = ~new_n45796_ & ~new_n45799_;
  assign new_n46156_ = ~new_n46154_ & ~new_n46155_;
  assign new_n46157_ = ~new_n45936_ & ~new_n46156_;
  assign new_n46158_ = ~new_n45477_ & ~new_n45935_;
  assign new_n46159_ = ~new_n45934_ & new_n46158_;
  assign new_n46160_ = ~new_n46157_ & ~new_n46159_;
  assign new_n46161_ = ~\b[25]  & ~new_n46160_;
  assign new_n46162_ = ~new_n45496_ & new_n45794_;
  assign new_n46163_ = ~new_n45790_ & new_n46162_;
  assign new_n46164_ = ~new_n45791_ & ~new_n45794_;
  assign new_n46165_ = ~new_n46163_ & ~new_n46164_;
  assign new_n46166_ = ~new_n45936_ & ~new_n46165_;
  assign new_n46167_ = ~new_n45486_ & ~new_n45935_;
  assign new_n46168_ = ~new_n45934_ & new_n46167_;
  assign new_n46169_ = ~new_n46166_ & ~new_n46168_;
  assign new_n46170_ = ~\b[24]  & ~new_n46169_;
  assign new_n46171_ = ~new_n45505_ & new_n45789_;
  assign new_n46172_ = ~new_n45785_ & new_n46171_;
  assign new_n46173_ = ~new_n45786_ & ~new_n45789_;
  assign new_n46174_ = ~new_n46172_ & ~new_n46173_;
  assign new_n46175_ = ~new_n45936_ & ~new_n46174_;
  assign new_n46176_ = ~new_n45495_ & ~new_n45935_;
  assign new_n46177_ = ~new_n45934_ & new_n46176_;
  assign new_n46178_ = ~new_n46175_ & ~new_n46177_;
  assign new_n46179_ = ~\b[23]  & ~new_n46178_;
  assign new_n46180_ = ~new_n45514_ & new_n45784_;
  assign new_n46181_ = ~new_n45780_ & new_n46180_;
  assign new_n46182_ = ~new_n45781_ & ~new_n45784_;
  assign new_n46183_ = ~new_n46181_ & ~new_n46182_;
  assign new_n46184_ = ~new_n45936_ & ~new_n46183_;
  assign new_n46185_ = ~new_n45504_ & ~new_n45935_;
  assign new_n46186_ = ~new_n45934_ & new_n46185_;
  assign new_n46187_ = ~new_n46184_ & ~new_n46186_;
  assign new_n46188_ = ~\b[22]  & ~new_n46187_;
  assign new_n46189_ = ~new_n45523_ & new_n45779_;
  assign new_n46190_ = ~new_n45775_ & new_n46189_;
  assign new_n46191_ = ~new_n45776_ & ~new_n45779_;
  assign new_n46192_ = ~new_n46190_ & ~new_n46191_;
  assign new_n46193_ = ~new_n45936_ & ~new_n46192_;
  assign new_n46194_ = ~new_n45513_ & ~new_n45935_;
  assign new_n46195_ = ~new_n45934_ & new_n46194_;
  assign new_n46196_ = ~new_n46193_ & ~new_n46195_;
  assign new_n46197_ = ~\b[21]  & ~new_n46196_;
  assign new_n46198_ = ~new_n45532_ & new_n45774_;
  assign new_n46199_ = ~new_n45770_ & new_n46198_;
  assign new_n46200_ = ~new_n45771_ & ~new_n45774_;
  assign new_n46201_ = ~new_n46199_ & ~new_n46200_;
  assign new_n46202_ = ~new_n45936_ & ~new_n46201_;
  assign new_n46203_ = ~new_n45522_ & ~new_n45935_;
  assign new_n46204_ = ~new_n45934_ & new_n46203_;
  assign new_n46205_ = ~new_n46202_ & ~new_n46204_;
  assign new_n46206_ = ~\b[20]  & ~new_n46205_;
  assign new_n46207_ = ~new_n45541_ & new_n45769_;
  assign new_n46208_ = ~new_n45765_ & new_n46207_;
  assign new_n46209_ = ~new_n45766_ & ~new_n45769_;
  assign new_n46210_ = ~new_n46208_ & ~new_n46209_;
  assign new_n46211_ = ~new_n45936_ & ~new_n46210_;
  assign new_n46212_ = ~new_n45531_ & ~new_n45935_;
  assign new_n46213_ = ~new_n45934_ & new_n46212_;
  assign new_n46214_ = ~new_n46211_ & ~new_n46213_;
  assign new_n46215_ = ~\b[19]  & ~new_n46214_;
  assign new_n46216_ = ~new_n45550_ & new_n45764_;
  assign new_n46217_ = ~new_n45760_ & new_n46216_;
  assign new_n46218_ = ~new_n45761_ & ~new_n45764_;
  assign new_n46219_ = ~new_n46217_ & ~new_n46218_;
  assign new_n46220_ = ~new_n45936_ & ~new_n46219_;
  assign new_n46221_ = ~new_n45540_ & ~new_n45935_;
  assign new_n46222_ = ~new_n45934_ & new_n46221_;
  assign new_n46223_ = ~new_n46220_ & ~new_n46222_;
  assign new_n46224_ = ~\b[18]  & ~new_n46223_;
  assign new_n46225_ = ~new_n45559_ & new_n45759_;
  assign new_n46226_ = ~new_n45755_ & new_n46225_;
  assign new_n46227_ = ~new_n45756_ & ~new_n45759_;
  assign new_n46228_ = ~new_n46226_ & ~new_n46227_;
  assign new_n46229_ = ~new_n45936_ & ~new_n46228_;
  assign new_n46230_ = ~new_n45549_ & ~new_n45935_;
  assign new_n46231_ = ~new_n45934_ & new_n46230_;
  assign new_n46232_ = ~new_n46229_ & ~new_n46231_;
  assign new_n46233_ = ~\b[17]  & ~new_n46232_;
  assign new_n46234_ = ~new_n45568_ & new_n45754_;
  assign new_n46235_ = ~new_n45750_ & new_n46234_;
  assign new_n46236_ = ~new_n45751_ & ~new_n45754_;
  assign new_n46237_ = ~new_n46235_ & ~new_n46236_;
  assign new_n46238_ = ~new_n45936_ & ~new_n46237_;
  assign new_n46239_ = ~new_n45558_ & ~new_n45935_;
  assign new_n46240_ = ~new_n45934_ & new_n46239_;
  assign new_n46241_ = ~new_n46238_ & ~new_n46240_;
  assign new_n46242_ = ~\b[16]  & ~new_n46241_;
  assign new_n46243_ = ~new_n45577_ & new_n45749_;
  assign new_n46244_ = ~new_n45745_ & new_n46243_;
  assign new_n46245_ = ~new_n45746_ & ~new_n45749_;
  assign new_n46246_ = ~new_n46244_ & ~new_n46245_;
  assign new_n46247_ = ~new_n45936_ & ~new_n46246_;
  assign new_n46248_ = ~new_n45567_ & ~new_n45935_;
  assign new_n46249_ = ~new_n45934_ & new_n46248_;
  assign new_n46250_ = ~new_n46247_ & ~new_n46249_;
  assign new_n46251_ = ~\b[15]  & ~new_n46250_;
  assign new_n46252_ = ~new_n45586_ & new_n45744_;
  assign new_n46253_ = ~new_n45740_ & new_n46252_;
  assign new_n46254_ = ~new_n45741_ & ~new_n45744_;
  assign new_n46255_ = ~new_n46253_ & ~new_n46254_;
  assign new_n46256_ = ~new_n45936_ & ~new_n46255_;
  assign new_n46257_ = ~new_n45576_ & ~new_n45935_;
  assign new_n46258_ = ~new_n45934_ & new_n46257_;
  assign new_n46259_ = ~new_n46256_ & ~new_n46258_;
  assign new_n46260_ = ~\b[14]  & ~new_n46259_;
  assign new_n46261_ = ~new_n45595_ & new_n45739_;
  assign new_n46262_ = ~new_n45735_ & new_n46261_;
  assign new_n46263_ = ~new_n45736_ & ~new_n45739_;
  assign new_n46264_ = ~new_n46262_ & ~new_n46263_;
  assign new_n46265_ = ~new_n45936_ & ~new_n46264_;
  assign new_n46266_ = ~new_n45585_ & ~new_n45935_;
  assign new_n46267_ = ~new_n45934_ & new_n46266_;
  assign new_n46268_ = ~new_n46265_ & ~new_n46267_;
  assign new_n46269_ = ~\b[13]  & ~new_n46268_;
  assign new_n46270_ = ~new_n45604_ & new_n45734_;
  assign new_n46271_ = ~new_n45730_ & new_n46270_;
  assign new_n46272_ = ~new_n45731_ & ~new_n45734_;
  assign new_n46273_ = ~new_n46271_ & ~new_n46272_;
  assign new_n46274_ = ~new_n45936_ & ~new_n46273_;
  assign new_n46275_ = ~new_n45594_ & ~new_n45935_;
  assign new_n46276_ = ~new_n45934_ & new_n46275_;
  assign new_n46277_ = ~new_n46274_ & ~new_n46276_;
  assign new_n46278_ = ~\b[12]  & ~new_n46277_;
  assign new_n46279_ = ~new_n45613_ & new_n45729_;
  assign new_n46280_ = ~new_n45725_ & new_n46279_;
  assign new_n46281_ = ~new_n45726_ & ~new_n45729_;
  assign new_n46282_ = ~new_n46280_ & ~new_n46281_;
  assign new_n46283_ = ~new_n45936_ & ~new_n46282_;
  assign new_n46284_ = ~new_n45603_ & ~new_n45935_;
  assign new_n46285_ = ~new_n45934_ & new_n46284_;
  assign new_n46286_ = ~new_n46283_ & ~new_n46285_;
  assign new_n46287_ = ~\b[11]  & ~new_n46286_;
  assign new_n46288_ = ~new_n45622_ & new_n45724_;
  assign new_n46289_ = ~new_n45720_ & new_n46288_;
  assign new_n46290_ = ~new_n45721_ & ~new_n45724_;
  assign new_n46291_ = ~new_n46289_ & ~new_n46290_;
  assign new_n46292_ = ~new_n45936_ & ~new_n46291_;
  assign new_n46293_ = ~new_n45612_ & ~new_n45935_;
  assign new_n46294_ = ~new_n45934_ & new_n46293_;
  assign new_n46295_ = ~new_n46292_ & ~new_n46294_;
  assign new_n46296_ = ~\b[10]  & ~new_n46295_;
  assign new_n46297_ = ~new_n45631_ & new_n45719_;
  assign new_n46298_ = ~new_n45715_ & new_n46297_;
  assign new_n46299_ = ~new_n45716_ & ~new_n45719_;
  assign new_n46300_ = ~new_n46298_ & ~new_n46299_;
  assign new_n46301_ = ~new_n45936_ & ~new_n46300_;
  assign new_n46302_ = ~new_n45621_ & ~new_n45935_;
  assign new_n46303_ = ~new_n45934_ & new_n46302_;
  assign new_n46304_ = ~new_n46301_ & ~new_n46303_;
  assign new_n46305_ = ~\b[9]  & ~new_n46304_;
  assign new_n46306_ = ~new_n45640_ & new_n45714_;
  assign new_n46307_ = ~new_n45710_ & new_n46306_;
  assign new_n46308_ = ~new_n45711_ & ~new_n45714_;
  assign new_n46309_ = ~new_n46307_ & ~new_n46308_;
  assign new_n46310_ = ~new_n45936_ & ~new_n46309_;
  assign new_n46311_ = ~new_n45630_ & ~new_n45935_;
  assign new_n46312_ = ~new_n45934_ & new_n46311_;
  assign new_n46313_ = ~new_n46310_ & ~new_n46312_;
  assign new_n46314_ = ~\b[8]  & ~new_n46313_;
  assign new_n46315_ = ~new_n45649_ & new_n45709_;
  assign new_n46316_ = ~new_n45705_ & new_n46315_;
  assign new_n46317_ = ~new_n45706_ & ~new_n45709_;
  assign new_n46318_ = ~new_n46316_ & ~new_n46317_;
  assign new_n46319_ = ~new_n45936_ & ~new_n46318_;
  assign new_n46320_ = ~new_n45639_ & ~new_n45935_;
  assign new_n46321_ = ~new_n45934_ & new_n46320_;
  assign new_n46322_ = ~new_n46319_ & ~new_n46321_;
  assign new_n46323_ = ~\b[7]  & ~new_n46322_;
  assign new_n46324_ = ~new_n45658_ & new_n45704_;
  assign new_n46325_ = ~new_n45700_ & new_n46324_;
  assign new_n46326_ = ~new_n45701_ & ~new_n45704_;
  assign new_n46327_ = ~new_n46325_ & ~new_n46326_;
  assign new_n46328_ = ~new_n45936_ & ~new_n46327_;
  assign new_n46329_ = ~new_n45648_ & ~new_n45935_;
  assign new_n46330_ = ~new_n45934_ & new_n46329_;
  assign new_n46331_ = ~new_n46328_ & ~new_n46330_;
  assign new_n46332_ = ~\b[6]  & ~new_n46331_;
  assign new_n46333_ = ~new_n45667_ & new_n45699_;
  assign new_n46334_ = ~new_n45695_ & new_n46333_;
  assign new_n46335_ = ~new_n45696_ & ~new_n45699_;
  assign new_n46336_ = ~new_n46334_ & ~new_n46335_;
  assign new_n46337_ = ~new_n45936_ & ~new_n46336_;
  assign new_n46338_ = ~new_n45657_ & ~new_n45935_;
  assign new_n46339_ = ~new_n45934_ & new_n46338_;
  assign new_n46340_ = ~new_n46337_ & ~new_n46339_;
  assign new_n46341_ = ~\b[5]  & ~new_n46340_;
  assign new_n46342_ = ~new_n45675_ & new_n45694_;
  assign new_n46343_ = ~new_n45690_ & new_n46342_;
  assign new_n46344_ = ~new_n45691_ & ~new_n45694_;
  assign new_n46345_ = ~new_n46343_ & ~new_n46344_;
  assign new_n46346_ = ~new_n45936_ & ~new_n46345_;
  assign new_n46347_ = ~new_n45666_ & ~new_n45935_;
  assign new_n46348_ = ~new_n45934_ & new_n46347_;
  assign new_n46349_ = ~new_n46346_ & ~new_n46348_;
  assign new_n46350_ = ~\b[4]  & ~new_n46349_;
  assign new_n46351_ = ~new_n45685_ & new_n45689_;
  assign new_n46352_ = ~new_n45684_ & new_n46351_;
  assign new_n46353_ = ~new_n45686_ & ~new_n45689_;
  assign new_n46354_ = ~new_n46352_ & ~new_n46353_;
  assign new_n46355_ = ~new_n45936_ & ~new_n46354_;
  assign new_n46356_ = ~new_n45674_ & ~new_n45935_;
  assign new_n46357_ = ~new_n45934_ & new_n46356_;
  assign new_n46358_ = ~new_n46355_ & ~new_n46357_;
  assign new_n46359_ = ~\b[3]  & ~new_n46358_;
  assign new_n46360_ = new_n17632_ & ~new_n45682_;
  assign new_n46361_ = ~new_n45680_ & new_n46360_;
  assign new_n46362_ = ~new_n45684_ & ~new_n46361_;
  assign new_n46363_ = ~new_n45936_ & new_n46362_;
  assign new_n46364_ = ~new_n45679_ & ~new_n45935_;
  assign new_n46365_ = ~new_n45934_ & new_n46364_;
  assign new_n46366_ = ~new_n46363_ & ~new_n46365_;
  assign new_n46367_ = ~\b[2]  & ~new_n46366_;
  assign new_n46368_ = \b[0]  & ~new_n45936_;
  assign new_n46369_ = \a[14]  & ~new_n46368_;
  assign new_n46370_ = new_n17632_ & ~new_n45936_;
  assign new_n46371_ = ~new_n46369_ & ~new_n46370_;
  assign new_n46372_ = \b[1]  & ~new_n46371_;
  assign new_n46373_ = ~\b[1]  & ~new_n46370_;
  assign new_n46374_ = ~new_n46369_ & new_n46373_;
  assign new_n46375_ = ~new_n46372_ & ~new_n46374_;
  assign new_n46376_ = ~new_n18327_ & ~new_n46375_;
  assign new_n46377_ = ~\b[1]  & ~new_n46371_;
  assign new_n46378_ = ~new_n46376_ & ~new_n46377_;
  assign new_n46379_ = \b[2]  & ~new_n46365_;
  assign new_n46380_ = ~new_n46363_ & new_n46379_;
  assign new_n46381_ = ~new_n46367_ & ~new_n46380_;
  assign new_n46382_ = ~new_n46378_ & new_n46381_;
  assign new_n46383_ = ~new_n46367_ & ~new_n46382_;
  assign new_n46384_ = \b[3]  & ~new_n46357_;
  assign new_n46385_ = ~new_n46355_ & new_n46384_;
  assign new_n46386_ = ~new_n46359_ & ~new_n46385_;
  assign new_n46387_ = ~new_n46383_ & new_n46386_;
  assign new_n46388_ = ~new_n46359_ & ~new_n46387_;
  assign new_n46389_ = \b[4]  & ~new_n46348_;
  assign new_n46390_ = ~new_n46346_ & new_n46389_;
  assign new_n46391_ = ~new_n46350_ & ~new_n46390_;
  assign new_n46392_ = ~new_n46388_ & new_n46391_;
  assign new_n46393_ = ~new_n46350_ & ~new_n46392_;
  assign new_n46394_ = \b[5]  & ~new_n46339_;
  assign new_n46395_ = ~new_n46337_ & new_n46394_;
  assign new_n46396_ = ~new_n46341_ & ~new_n46395_;
  assign new_n46397_ = ~new_n46393_ & new_n46396_;
  assign new_n46398_ = ~new_n46341_ & ~new_n46397_;
  assign new_n46399_ = \b[6]  & ~new_n46330_;
  assign new_n46400_ = ~new_n46328_ & new_n46399_;
  assign new_n46401_ = ~new_n46332_ & ~new_n46400_;
  assign new_n46402_ = ~new_n46398_ & new_n46401_;
  assign new_n46403_ = ~new_n46332_ & ~new_n46402_;
  assign new_n46404_ = \b[7]  & ~new_n46321_;
  assign new_n46405_ = ~new_n46319_ & new_n46404_;
  assign new_n46406_ = ~new_n46323_ & ~new_n46405_;
  assign new_n46407_ = ~new_n46403_ & new_n46406_;
  assign new_n46408_ = ~new_n46323_ & ~new_n46407_;
  assign new_n46409_ = \b[8]  & ~new_n46312_;
  assign new_n46410_ = ~new_n46310_ & new_n46409_;
  assign new_n46411_ = ~new_n46314_ & ~new_n46410_;
  assign new_n46412_ = ~new_n46408_ & new_n46411_;
  assign new_n46413_ = ~new_n46314_ & ~new_n46412_;
  assign new_n46414_ = \b[9]  & ~new_n46303_;
  assign new_n46415_ = ~new_n46301_ & new_n46414_;
  assign new_n46416_ = ~new_n46305_ & ~new_n46415_;
  assign new_n46417_ = ~new_n46413_ & new_n46416_;
  assign new_n46418_ = ~new_n46305_ & ~new_n46417_;
  assign new_n46419_ = \b[10]  & ~new_n46294_;
  assign new_n46420_ = ~new_n46292_ & new_n46419_;
  assign new_n46421_ = ~new_n46296_ & ~new_n46420_;
  assign new_n46422_ = ~new_n46418_ & new_n46421_;
  assign new_n46423_ = ~new_n46296_ & ~new_n46422_;
  assign new_n46424_ = \b[11]  & ~new_n46285_;
  assign new_n46425_ = ~new_n46283_ & new_n46424_;
  assign new_n46426_ = ~new_n46287_ & ~new_n46425_;
  assign new_n46427_ = ~new_n46423_ & new_n46426_;
  assign new_n46428_ = ~new_n46287_ & ~new_n46427_;
  assign new_n46429_ = \b[12]  & ~new_n46276_;
  assign new_n46430_ = ~new_n46274_ & new_n46429_;
  assign new_n46431_ = ~new_n46278_ & ~new_n46430_;
  assign new_n46432_ = ~new_n46428_ & new_n46431_;
  assign new_n46433_ = ~new_n46278_ & ~new_n46432_;
  assign new_n46434_ = \b[13]  & ~new_n46267_;
  assign new_n46435_ = ~new_n46265_ & new_n46434_;
  assign new_n46436_ = ~new_n46269_ & ~new_n46435_;
  assign new_n46437_ = ~new_n46433_ & new_n46436_;
  assign new_n46438_ = ~new_n46269_ & ~new_n46437_;
  assign new_n46439_ = \b[14]  & ~new_n46258_;
  assign new_n46440_ = ~new_n46256_ & new_n46439_;
  assign new_n46441_ = ~new_n46260_ & ~new_n46440_;
  assign new_n46442_ = ~new_n46438_ & new_n46441_;
  assign new_n46443_ = ~new_n46260_ & ~new_n46442_;
  assign new_n46444_ = \b[15]  & ~new_n46249_;
  assign new_n46445_ = ~new_n46247_ & new_n46444_;
  assign new_n46446_ = ~new_n46251_ & ~new_n46445_;
  assign new_n46447_ = ~new_n46443_ & new_n46446_;
  assign new_n46448_ = ~new_n46251_ & ~new_n46447_;
  assign new_n46449_ = \b[16]  & ~new_n46240_;
  assign new_n46450_ = ~new_n46238_ & new_n46449_;
  assign new_n46451_ = ~new_n46242_ & ~new_n46450_;
  assign new_n46452_ = ~new_n46448_ & new_n46451_;
  assign new_n46453_ = ~new_n46242_ & ~new_n46452_;
  assign new_n46454_ = \b[17]  & ~new_n46231_;
  assign new_n46455_ = ~new_n46229_ & new_n46454_;
  assign new_n46456_ = ~new_n46233_ & ~new_n46455_;
  assign new_n46457_ = ~new_n46453_ & new_n46456_;
  assign new_n46458_ = ~new_n46233_ & ~new_n46457_;
  assign new_n46459_ = \b[18]  & ~new_n46222_;
  assign new_n46460_ = ~new_n46220_ & new_n46459_;
  assign new_n46461_ = ~new_n46224_ & ~new_n46460_;
  assign new_n46462_ = ~new_n46458_ & new_n46461_;
  assign new_n46463_ = ~new_n46224_ & ~new_n46462_;
  assign new_n46464_ = \b[19]  & ~new_n46213_;
  assign new_n46465_ = ~new_n46211_ & new_n46464_;
  assign new_n46466_ = ~new_n46215_ & ~new_n46465_;
  assign new_n46467_ = ~new_n46463_ & new_n46466_;
  assign new_n46468_ = ~new_n46215_ & ~new_n46467_;
  assign new_n46469_ = \b[20]  & ~new_n46204_;
  assign new_n46470_ = ~new_n46202_ & new_n46469_;
  assign new_n46471_ = ~new_n46206_ & ~new_n46470_;
  assign new_n46472_ = ~new_n46468_ & new_n46471_;
  assign new_n46473_ = ~new_n46206_ & ~new_n46472_;
  assign new_n46474_ = \b[21]  & ~new_n46195_;
  assign new_n46475_ = ~new_n46193_ & new_n46474_;
  assign new_n46476_ = ~new_n46197_ & ~new_n46475_;
  assign new_n46477_ = ~new_n46473_ & new_n46476_;
  assign new_n46478_ = ~new_n46197_ & ~new_n46477_;
  assign new_n46479_ = \b[22]  & ~new_n46186_;
  assign new_n46480_ = ~new_n46184_ & new_n46479_;
  assign new_n46481_ = ~new_n46188_ & ~new_n46480_;
  assign new_n46482_ = ~new_n46478_ & new_n46481_;
  assign new_n46483_ = ~new_n46188_ & ~new_n46482_;
  assign new_n46484_ = \b[23]  & ~new_n46177_;
  assign new_n46485_ = ~new_n46175_ & new_n46484_;
  assign new_n46486_ = ~new_n46179_ & ~new_n46485_;
  assign new_n46487_ = ~new_n46483_ & new_n46486_;
  assign new_n46488_ = ~new_n46179_ & ~new_n46487_;
  assign new_n46489_ = \b[24]  & ~new_n46168_;
  assign new_n46490_ = ~new_n46166_ & new_n46489_;
  assign new_n46491_ = ~new_n46170_ & ~new_n46490_;
  assign new_n46492_ = ~new_n46488_ & new_n46491_;
  assign new_n46493_ = ~new_n46170_ & ~new_n46492_;
  assign new_n46494_ = \b[25]  & ~new_n46159_;
  assign new_n46495_ = ~new_n46157_ & new_n46494_;
  assign new_n46496_ = ~new_n46161_ & ~new_n46495_;
  assign new_n46497_ = ~new_n46493_ & new_n46496_;
  assign new_n46498_ = ~new_n46161_ & ~new_n46497_;
  assign new_n46499_ = \b[26]  & ~new_n46150_;
  assign new_n46500_ = ~new_n46148_ & new_n46499_;
  assign new_n46501_ = ~new_n46152_ & ~new_n46500_;
  assign new_n46502_ = ~new_n46498_ & new_n46501_;
  assign new_n46503_ = ~new_n46152_ & ~new_n46502_;
  assign new_n46504_ = \b[27]  & ~new_n46141_;
  assign new_n46505_ = ~new_n46139_ & new_n46504_;
  assign new_n46506_ = ~new_n46143_ & ~new_n46505_;
  assign new_n46507_ = ~new_n46503_ & new_n46506_;
  assign new_n46508_ = ~new_n46143_ & ~new_n46507_;
  assign new_n46509_ = \b[28]  & ~new_n46132_;
  assign new_n46510_ = ~new_n46130_ & new_n46509_;
  assign new_n46511_ = ~new_n46134_ & ~new_n46510_;
  assign new_n46512_ = ~new_n46508_ & new_n46511_;
  assign new_n46513_ = ~new_n46134_ & ~new_n46512_;
  assign new_n46514_ = \b[29]  & ~new_n46123_;
  assign new_n46515_ = ~new_n46121_ & new_n46514_;
  assign new_n46516_ = ~new_n46125_ & ~new_n46515_;
  assign new_n46517_ = ~new_n46513_ & new_n46516_;
  assign new_n46518_ = ~new_n46125_ & ~new_n46517_;
  assign new_n46519_ = \b[30]  & ~new_n46114_;
  assign new_n46520_ = ~new_n46112_ & new_n46519_;
  assign new_n46521_ = ~new_n46116_ & ~new_n46520_;
  assign new_n46522_ = ~new_n46518_ & new_n46521_;
  assign new_n46523_ = ~new_n46116_ & ~new_n46522_;
  assign new_n46524_ = \b[31]  & ~new_n46105_;
  assign new_n46525_ = ~new_n46103_ & new_n46524_;
  assign new_n46526_ = ~new_n46107_ & ~new_n46525_;
  assign new_n46527_ = ~new_n46523_ & new_n46526_;
  assign new_n46528_ = ~new_n46107_ & ~new_n46527_;
  assign new_n46529_ = \b[32]  & ~new_n46096_;
  assign new_n46530_ = ~new_n46094_ & new_n46529_;
  assign new_n46531_ = ~new_n46098_ & ~new_n46530_;
  assign new_n46532_ = ~new_n46528_ & new_n46531_;
  assign new_n46533_ = ~new_n46098_ & ~new_n46532_;
  assign new_n46534_ = \b[33]  & ~new_n46087_;
  assign new_n46535_ = ~new_n46085_ & new_n46534_;
  assign new_n46536_ = ~new_n46089_ & ~new_n46535_;
  assign new_n46537_ = ~new_n46533_ & new_n46536_;
  assign new_n46538_ = ~new_n46089_ & ~new_n46537_;
  assign new_n46539_ = \b[34]  & ~new_n46078_;
  assign new_n46540_ = ~new_n46076_ & new_n46539_;
  assign new_n46541_ = ~new_n46080_ & ~new_n46540_;
  assign new_n46542_ = ~new_n46538_ & new_n46541_;
  assign new_n46543_ = ~new_n46080_ & ~new_n46542_;
  assign new_n46544_ = \b[35]  & ~new_n46069_;
  assign new_n46545_ = ~new_n46067_ & new_n46544_;
  assign new_n46546_ = ~new_n46071_ & ~new_n46545_;
  assign new_n46547_ = ~new_n46543_ & new_n46546_;
  assign new_n46548_ = ~new_n46071_ & ~new_n46547_;
  assign new_n46549_ = \b[36]  & ~new_n46060_;
  assign new_n46550_ = ~new_n46058_ & new_n46549_;
  assign new_n46551_ = ~new_n46062_ & ~new_n46550_;
  assign new_n46552_ = ~new_n46548_ & new_n46551_;
  assign new_n46553_ = ~new_n46062_ & ~new_n46552_;
  assign new_n46554_ = \b[37]  & ~new_n46051_;
  assign new_n46555_ = ~new_n46049_ & new_n46554_;
  assign new_n46556_ = ~new_n46053_ & ~new_n46555_;
  assign new_n46557_ = ~new_n46553_ & new_n46556_;
  assign new_n46558_ = ~new_n46053_ & ~new_n46557_;
  assign new_n46559_ = \b[38]  & ~new_n46042_;
  assign new_n46560_ = ~new_n46040_ & new_n46559_;
  assign new_n46561_ = ~new_n46044_ & ~new_n46560_;
  assign new_n46562_ = ~new_n46558_ & new_n46561_;
  assign new_n46563_ = ~new_n46044_ & ~new_n46562_;
  assign new_n46564_ = \b[39]  & ~new_n46033_;
  assign new_n46565_ = ~new_n46031_ & new_n46564_;
  assign new_n46566_ = ~new_n46035_ & ~new_n46565_;
  assign new_n46567_ = ~new_n46563_ & new_n46566_;
  assign new_n46568_ = ~new_n46035_ & ~new_n46567_;
  assign new_n46569_ = \b[40]  & ~new_n46024_;
  assign new_n46570_ = ~new_n46022_ & new_n46569_;
  assign new_n46571_ = ~new_n46026_ & ~new_n46570_;
  assign new_n46572_ = ~new_n46568_ & new_n46571_;
  assign new_n46573_ = ~new_n46026_ & ~new_n46572_;
  assign new_n46574_ = \b[41]  & ~new_n46015_;
  assign new_n46575_ = ~new_n46013_ & new_n46574_;
  assign new_n46576_ = ~new_n46017_ & ~new_n46575_;
  assign new_n46577_ = ~new_n46573_ & new_n46576_;
  assign new_n46578_ = ~new_n46017_ & ~new_n46577_;
  assign new_n46579_ = \b[42]  & ~new_n46006_;
  assign new_n46580_ = ~new_n46004_ & new_n46579_;
  assign new_n46581_ = ~new_n46008_ & ~new_n46580_;
  assign new_n46582_ = ~new_n46578_ & new_n46581_;
  assign new_n46583_ = ~new_n46008_ & ~new_n46582_;
  assign new_n46584_ = \b[43]  & ~new_n45997_;
  assign new_n46585_ = ~new_n45995_ & new_n46584_;
  assign new_n46586_ = ~new_n45999_ & ~new_n46585_;
  assign new_n46587_ = ~new_n46583_ & new_n46586_;
  assign new_n46588_ = ~new_n45999_ & ~new_n46587_;
  assign new_n46589_ = \b[44]  & ~new_n45988_;
  assign new_n46590_ = ~new_n45986_ & new_n46589_;
  assign new_n46591_ = ~new_n45990_ & ~new_n46590_;
  assign new_n46592_ = ~new_n46588_ & new_n46591_;
  assign new_n46593_ = ~new_n45990_ & ~new_n46592_;
  assign new_n46594_ = \b[45]  & ~new_n45979_;
  assign new_n46595_ = ~new_n45977_ & new_n46594_;
  assign new_n46596_ = ~new_n45981_ & ~new_n46595_;
  assign new_n46597_ = ~new_n46593_ & new_n46596_;
  assign new_n46598_ = ~new_n45981_ & ~new_n46597_;
  assign new_n46599_ = \b[46]  & ~new_n45970_;
  assign new_n46600_ = ~new_n45968_ & new_n46599_;
  assign new_n46601_ = ~new_n45972_ & ~new_n46600_;
  assign new_n46602_ = ~new_n46598_ & new_n46601_;
  assign new_n46603_ = ~new_n45972_ & ~new_n46602_;
  assign new_n46604_ = \b[47]  & ~new_n45961_;
  assign new_n46605_ = ~new_n45959_ & new_n46604_;
  assign new_n46606_ = ~new_n45963_ & ~new_n46605_;
  assign new_n46607_ = ~new_n46603_ & new_n46606_;
  assign new_n46608_ = ~new_n45963_ & ~new_n46607_;
  assign new_n46609_ = \b[48]  & ~new_n45952_;
  assign new_n46610_ = ~new_n45950_ & new_n46609_;
  assign new_n46611_ = ~new_n45954_ & ~new_n46610_;
  assign new_n46612_ = ~new_n46608_ & new_n46611_;
  assign new_n46613_ = ~new_n45954_ & ~new_n46612_;
  assign new_n46614_ = \b[49]  & ~new_n45943_;
  assign new_n46615_ = ~new_n45941_ & new_n46614_;
  assign new_n46616_ = ~new_n45945_ & ~new_n46615_;
  assign new_n46617_ = ~new_n46613_ & new_n46616_;
  assign new_n46618_ = ~new_n45945_ & ~new_n46617_;
  assign new_n46619_ = ~new_n45262_ & ~new_n45931_;
  assign new_n46620_ = ~new_n45929_ & new_n46619_;
  assign new_n46621_ = ~new_n45920_ & new_n46620_;
  assign new_n46622_ = ~new_n45929_ & ~new_n45931_;
  assign new_n46623_ = ~new_n45921_ & ~new_n46622_;
  assign new_n46624_ = ~new_n46621_ & ~new_n46623_;
  assign new_n46625_ = ~new_n45936_ & ~new_n46624_;
  assign new_n46626_ = ~new_n45928_ & ~new_n45935_;
  assign new_n46627_ = ~new_n45934_ & new_n46626_;
  assign new_n46628_ = ~new_n46625_ & ~new_n46627_;
  assign new_n46629_ = ~\b[50]  & ~new_n46628_;
  assign new_n46630_ = \b[50]  & ~new_n46627_;
  assign new_n46631_ = ~new_n46625_ & new_n46630_;
  assign new_n46632_ = new_n18585_ & ~new_n46631_;
  assign new_n46633_ = ~new_n46629_ & new_n46632_;
  assign new_n46634_ = ~new_n46618_ & new_n46633_;
  assign new_n46635_ = new_n17882_ & ~new_n46628_;
  assign new_n46636_ = ~new_n46634_ & ~new_n46635_;
  assign new_n46637_ = ~new_n45954_ & new_n46616_;
  assign new_n46638_ = ~new_n46612_ & new_n46637_;
  assign new_n46639_ = ~new_n46613_ & ~new_n46616_;
  assign new_n46640_ = ~new_n46638_ & ~new_n46639_;
  assign new_n46641_ = ~new_n46636_ & ~new_n46640_;
  assign new_n46642_ = ~new_n45944_ & ~new_n46635_;
  assign new_n46643_ = ~new_n46634_ & new_n46642_;
  assign new_n46644_ = ~new_n46641_ & ~new_n46643_;
  assign new_n46645_ = ~new_n45945_ & ~new_n46631_;
  assign new_n46646_ = ~new_n46629_ & new_n46645_;
  assign new_n46647_ = ~new_n46617_ & new_n46646_;
  assign new_n46648_ = ~new_n46629_ & ~new_n46631_;
  assign new_n46649_ = ~new_n46618_ & ~new_n46648_;
  assign new_n46650_ = ~new_n46647_ & ~new_n46649_;
  assign new_n46651_ = ~new_n46636_ & ~new_n46650_;
  assign new_n46652_ = ~new_n46628_ & ~new_n46635_;
  assign new_n46653_ = ~new_n46634_ & new_n46652_;
  assign new_n46654_ = ~new_n46651_ & ~new_n46653_;
  assign new_n46655_ = ~\b[51]  & ~new_n46654_;
  assign new_n46656_ = ~\b[50]  & ~new_n46644_;
  assign new_n46657_ = ~new_n45963_ & new_n46611_;
  assign new_n46658_ = ~new_n46607_ & new_n46657_;
  assign new_n46659_ = ~new_n46608_ & ~new_n46611_;
  assign new_n46660_ = ~new_n46658_ & ~new_n46659_;
  assign new_n46661_ = ~new_n46636_ & ~new_n46660_;
  assign new_n46662_ = ~new_n45953_ & ~new_n46635_;
  assign new_n46663_ = ~new_n46634_ & new_n46662_;
  assign new_n46664_ = ~new_n46661_ & ~new_n46663_;
  assign new_n46665_ = ~\b[49]  & ~new_n46664_;
  assign new_n46666_ = ~new_n45972_ & new_n46606_;
  assign new_n46667_ = ~new_n46602_ & new_n46666_;
  assign new_n46668_ = ~new_n46603_ & ~new_n46606_;
  assign new_n46669_ = ~new_n46667_ & ~new_n46668_;
  assign new_n46670_ = ~new_n46636_ & ~new_n46669_;
  assign new_n46671_ = ~new_n45962_ & ~new_n46635_;
  assign new_n46672_ = ~new_n46634_ & new_n46671_;
  assign new_n46673_ = ~new_n46670_ & ~new_n46672_;
  assign new_n46674_ = ~\b[48]  & ~new_n46673_;
  assign new_n46675_ = ~new_n45981_ & new_n46601_;
  assign new_n46676_ = ~new_n46597_ & new_n46675_;
  assign new_n46677_ = ~new_n46598_ & ~new_n46601_;
  assign new_n46678_ = ~new_n46676_ & ~new_n46677_;
  assign new_n46679_ = ~new_n46636_ & ~new_n46678_;
  assign new_n46680_ = ~new_n45971_ & ~new_n46635_;
  assign new_n46681_ = ~new_n46634_ & new_n46680_;
  assign new_n46682_ = ~new_n46679_ & ~new_n46681_;
  assign new_n46683_ = ~\b[47]  & ~new_n46682_;
  assign new_n46684_ = ~new_n45990_ & new_n46596_;
  assign new_n46685_ = ~new_n46592_ & new_n46684_;
  assign new_n46686_ = ~new_n46593_ & ~new_n46596_;
  assign new_n46687_ = ~new_n46685_ & ~new_n46686_;
  assign new_n46688_ = ~new_n46636_ & ~new_n46687_;
  assign new_n46689_ = ~new_n45980_ & ~new_n46635_;
  assign new_n46690_ = ~new_n46634_ & new_n46689_;
  assign new_n46691_ = ~new_n46688_ & ~new_n46690_;
  assign new_n46692_ = ~\b[46]  & ~new_n46691_;
  assign new_n46693_ = ~new_n45999_ & new_n46591_;
  assign new_n46694_ = ~new_n46587_ & new_n46693_;
  assign new_n46695_ = ~new_n46588_ & ~new_n46591_;
  assign new_n46696_ = ~new_n46694_ & ~new_n46695_;
  assign new_n46697_ = ~new_n46636_ & ~new_n46696_;
  assign new_n46698_ = ~new_n45989_ & ~new_n46635_;
  assign new_n46699_ = ~new_n46634_ & new_n46698_;
  assign new_n46700_ = ~new_n46697_ & ~new_n46699_;
  assign new_n46701_ = ~\b[45]  & ~new_n46700_;
  assign new_n46702_ = ~new_n46008_ & new_n46586_;
  assign new_n46703_ = ~new_n46582_ & new_n46702_;
  assign new_n46704_ = ~new_n46583_ & ~new_n46586_;
  assign new_n46705_ = ~new_n46703_ & ~new_n46704_;
  assign new_n46706_ = ~new_n46636_ & ~new_n46705_;
  assign new_n46707_ = ~new_n45998_ & ~new_n46635_;
  assign new_n46708_ = ~new_n46634_ & new_n46707_;
  assign new_n46709_ = ~new_n46706_ & ~new_n46708_;
  assign new_n46710_ = ~\b[44]  & ~new_n46709_;
  assign new_n46711_ = ~new_n46017_ & new_n46581_;
  assign new_n46712_ = ~new_n46577_ & new_n46711_;
  assign new_n46713_ = ~new_n46578_ & ~new_n46581_;
  assign new_n46714_ = ~new_n46712_ & ~new_n46713_;
  assign new_n46715_ = ~new_n46636_ & ~new_n46714_;
  assign new_n46716_ = ~new_n46007_ & ~new_n46635_;
  assign new_n46717_ = ~new_n46634_ & new_n46716_;
  assign new_n46718_ = ~new_n46715_ & ~new_n46717_;
  assign new_n46719_ = ~\b[43]  & ~new_n46718_;
  assign new_n46720_ = ~new_n46026_ & new_n46576_;
  assign new_n46721_ = ~new_n46572_ & new_n46720_;
  assign new_n46722_ = ~new_n46573_ & ~new_n46576_;
  assign new_n46723_ = ~new_n46721_ & ~new_n46722_;
  assign new_n46724_ = ~new_n46636_ & ~new_n46723_;
  assign new_n46725_ = ~new_n46016_ & ~new_n46635_;
  assign new_n46726_ = ~new_n46634_ & new_n46725_;
  assign new_n46727_ = ~new_n46724_ & ~new_n46726_;
  assign new_n46728_ = ~\b[42]  & ~new_n46727_;
  assign new_n46729_ = ~new_n46035_ & new_n46571_;
  assign new_n46730_ = ~new_n46567_ & new_n46729_;
  assign new_n46731_ = ~new_n46568_ & ~new_n46571_;
  assign new_n46732_ = ~new_n46730_ & ~new_n46731_;
  assign new_n46733_ = ~new_n46636_ & ~new_n46732_;
  assign new_n46734_ = ~new_n46025_ & ~new_n46635_;
  assign new_n46735_ = ~new_n46634_ & new_n46734_;
  assign new_n46736_ = ~new_n46733_ & ~new_n46735_;
  assign new_n46737_ = ~\b[41]  & ~new_n46736_;
  assign new_n46738_ = ~new_n46044_ & new_n46566_;
  assign new_n46739_ = ~new_n46562_ & new_n46738_;
  assign new_n46740_ = ~new_n46563_ & ~new_n46566_;
  assign new_n46741_ = ~new_n46739_ & ~new_n46740_;
  assign new_n46742_ = ~new_n46636_ & ~new_n46741_;
  assign new_n46743_ = ~new_n46034_ & ~new_n46635_;
  assign new_n46744_ = ~new_n46634_ & new_n46743_;
  assign new_n46745_ = ~new_n46742_ & ~new_n46744_;
  assign new_n46746_ = ~\b[40]  & ~new_n46745_;
  assign new_n46747_ = ~new_n46053_ & new_n46561_;
  assign new_n46748_ = ~new_n46557_ & new_n46747_;
  assign new_n46749_ = ~new_n46558_ & ~new_n46561_;
  assign new_n46750_ = ~new_n46748_ & ~new_n46749_;
  assign new_n46751_ = ~new_n46636_ & ~new_n46750_;
  assign new_n46752_ = ~new_n46043_ & ~new_n46635_;
  assign new_n46753_ = ~new_n46634_ & new_n46752_;
  assign new_n46754_ = ~new_n46751_ & ~new_n46753_;
  assign new_n46755_ = ~\b[39]  & ~new_n46754_;
  assign new_n46756_ = ~new_n46062_ & new_n46556_;
  assign new_n46757_ = ~new_n46552_ & new_n46756_;
  assign new_n46758_ = ~new_n46553_ & ~new_n46556_;
  assign new_n46759_ = ~new_n46757_ & ~new_n46758_;
  assign new_n46760_ = ~new_n46636_ & ~new_n46759_;
  assign new_n46761_ = ~new_n46052_ & ~new_n46635_;
  assign new_n46762_ = ~new_n46634_ & new_n46761_;
  assign new_n46763_ = ~new_n46760_ & ~new_n46762_;
  assign new_n46764_ = ~\b[38]  & ~new_n46763_;
  assign new_n46765_ = ~new_n46071_ & new_n46551_;
  assign new_n46766_ = ~new_n46547_ & new_n46765_;
  assign new_n46767_ = ~new_n46548_ & ~new_n46551_;
  assign new_n46768_ = ~new_n46766_ & ~new_n46767_;
  assign new_n46769_ = ~new_n46636_ & ~new_n46768_;
  assign new_n46770_ = ~new_n46061_ & ~new_n46635_;
  assign new_n46771_ = ~new_n46634_ & new_n46770_;
  assign new_n46772_ = ~new_n46769_ & ~new_n46771_;
  assign new_n46773_ = ~\b[37]  & ~new_n46772_;
  assign new_n46774_ = ~new_n46080_ & new_n46546_;
  assign new_n46775_ = ~new_n46542_ & new_n46774_;
  assign new_n46776_ = ~new_n46543_ & ~new_n46546_;
  assign new_n46777_ = ~new_n46775_ & ~new_n46776_;
  assign new_n46778_ = ~new_n46636_ & ~new_n46777_;
  assign new_n46779_ = ~new_n46070_ & ~new_n46635_;
  assign new_n46780_ = ~new_n46634_ & new_n46779_;
  assign new_n46781_ = ~new_n46778_ & ~new_n46780_;
  assign new_n46782_ = ~\b[36]  & ~new_n46781_;
  assign new_n46783_ = ~new_n46089_ & new_n46541_;
  assign new_n46784_ = ~new_n46537_ & new_n46783_;
  assign new_n46785_ = ~new_n46538_ & ~new_n46541_;
  assign new_n46786_ = ~new_n46784_ & ~new_n46785_;
  assign new_n46787_ = ~new_n46636_ & ~new_n46786_;
  assign new_n46788_ = ~new_n46079_ & ~new_n46635_;
  assign new_n46789_ = ~new_n46634_ & new_n46788_;
  assign new_n46790_ = ~new_n46787_ & ~new_n46789_;
  assign new_n46791_ = ~\b[35]  & ~new_n46790_;
  assign new_n46792_ = ~new_n46098_ & new_n46536_;
  assign new_n46793_ = ~new_n46532_ & new_n46792_;
  assign new_n46794_ = ~new_n46533_ & ~new_n46536_;
  assign new_n46795_ = ~new_n46793_ & ~new_n46794_;
  assign new_n46796_ = ~new_n46636_ & ~new_n46795_;
  assign new_n46797_ = ~new_n46088_ & ~new_n46635_;
  assign new_n46798_ = ~new_n46634_ & new_n46797_;
  assign new_n46799_ = ~new_n46796_ & ~new_n46798_;
  assign new_n46800_ = ~\b[34]  & ~new_n46799_;
  assign new_n46801_ = ~new_n46107_ & new_n46531_;
  assign new_n46802_ = ~new_n46527_ & new_n46801_;
  assign new_n46803_ = ~new_n46528_ & ~new_n46531_;
  assign new_n46804_ = ~new_n46802_ & ~new_n46803_;
  assign new_n46805_ = ~new_n46636_ & ~new_n46804_;
  assign new_n46806_ = ~new_n46097_ & ~new_n46635_;
  assign new_n46807_ = ~new_n46634_ & new_n46806_;
  assign new_n46808_ = ~new_n46805_ & ~new_n46807_;
  assign new_n46809_ = ~\b[33]  & ~new_n46808_;
  assign new_n46810_ = ~new_n46116_ & new_n46526_;
  assign new_n46811_ = ~new_n46522_ & new_n46810_;
  assign new_n46812_ = ~new_n46523_ & ~new_n46526_;
  assign new_n46813_ = ~new_n46811_ & ~new_n46812_;
  assign new_n46814_ = ~new_n46636_ & ~new_n46813_;
  assign new_n46815_ = ~new_n46106_ & ~new_n46635_;
  assign new_n46816_ = ~new_n46634_ & new_n46815_;
  assign new_n46817_ = ~new_n46814_ & ~new_n46816_;
  assign new_n46818_ = ~\b[32]  & ~new_n46817_;
  assign new_n46819_ = ~new_n46125_ & new_n46521_;
  assign new_n46820_ = ~new_n46517_ & new_n46819_;
  assign new_n46821_ = ~new_n46518_ & ~new_n46521_;
  assign new_n46822_ = ~new_n46820_ & ~new_n46821_;
  assign new_n46823_ = ~new_n46636_ & ~new_n46822_;
  assign new_n46824_ = ~new_n46115_ & ~new_n46635_;
  assign new_n46825_ = ~new_n46634_ & new_n46824_;
  assign new_n46826_ = ~new_n46823_ & ~new_n46825_;
  assign new_n46827_ = ~\b[31]  & ~new_n46826_;
  assign new_n46828_ = ~new_n46134_ & new_n46516_;
  assign new_n46829_ = ~new_n46512_ & new_n46828_;
  assign new_n46830_ = ~new_n46513_ & ~new_n46516_;
  assign new_n46831_ = ~new_n46829_ & ~new_n46830_;
  assign new_n46832_ = ~new_n46636_ & ~new_n46831_;
  assign new_n46833_ = ~new_n46124_ & ~new_n46635_;
  assign new_n46834_ = ~new_n46634_ & new_n46833_;
  assign new_n46835_ = ~new_n46832_ & ~new_n46834_;
  assign new_n46836_ = ~\b[30]  & ~new_n46835_;
  assign new_n46837_ = ~new_n46143_ & new_n46511_;
  assign new_n46838_ = ~new_n46507_ & new_n46837_;
  assign new_n46839_ = ~new_n46508_ & ~new_n46511_;
  assign new_n46840_ = ~new_n46838_ & ~new_n46839_;
  assign new_n46841_ = ~new_n46636_ & ~new_n46840_;
  assign new_n46842_ = ~new_n46133_ & ~new_n46635_;
  assign new_n46843_ = ~new_n46634_ & new_n46842_;
  assign new_n46844_ = ~new_n46841_ & ~new_n46843_;
  assign new_n46845_ = ~\b[29]  & ~new_n46844_;
  assign new_n46846_ = ~new_n46152_ & new_n46506_;
  assign new_n46847_ = ~new_n46502_ & new_n46846_;
  assign new_n46848_ = ~new_n46503_ & ~new_n46506_;
  assign new_n46849_ = ~new_n46847_ & ~new_n46848_;
  assign new_n46850_ = ~new_n46636_ & ~new_n46849_;
  assign new_n46851_ = ~new_n46142_ & ~new_n46635_;
  assign new_n46852_ = ~new_n46634_ & new_n46851_;
  assign new_n46853_ = ~new_n46850_ & ~new_n46852_;
  assign new_n46854_ = ~\b[28]  & ~new_n46853_;
  assign new_n46855_ = ~new_n46161_ & new_n46501_;
  assign new_n46856_ = ~new_n46497_ & new_n46855_;
  assign new_n46857_ = ~new_n46498_ & ~new_n46501_;
  assign new_n46858_ = ~new_n46856_ & ~new_n46857_;
  assign new_n46859_ = ~new_n46636_ & ~new_n46858_;
  assign new_n46860_ = ~new_n46151_ & ~new_n46635_;
  assign new_n46861_ = ~new_n46634_ & new_n46860_;
  assign new_n46862_ = ~new_n46859_ & ~new_n46861_;
  assign new_n46863_ = ~\b[27]  & ~new_n46862_;
  assign new_n46864_ = ~new_n46170_ & new_n46496_;
  assign new_n46865_ = ~new_n46492_ & new_n46864_;
  assign new_n46866_ = ~new_n46493_ & ~new_n46496_;
  assign new_n46867_ = ~new_n46865_ & ~new_n46866_;
  assign new_n46868_ = ~new_n46636_ & ~new_n46867_;
  assign new_n46869_ = ~new_n46160_ & ~new_n46635_;
  assign new_n46870_ = ~new_n46634_ & new_n46869_;
  assign new_n46871_ = ~new_n46868_ & ~new_n46870_;
  assign new_n46872_ = ~\b[26]  & ~new_n46871_;
  assign new_n46873_ = ~new_n46179_ & new_n46491_;
  assign new_n46874_ = ~new_n46487_ & new_n46873_;
  assign new_n46875_ = ~new_n46488_ & ~new_n46491_;
  assign new_n46876_ = ~new_n46874_ & ~new_n46875_;
  assign new_n46877_ = ~new_n46636_ & ~new_n46876_;
  assign new_n46878_ = ~new_n46169_ & ~new_n46635_;
  assign new_n46879_ = ~new_n46634_ & new_n46878_;
  assign new_n46880_ = ~new_n46877_ & ~new_n46879_;
  assign new_n46881_ = ~\b[25]  & ~new_n46880_;
  assign new_n46882_ = ~new_n46188_ & new_n46486_;
  assign new_n46883_ = ~new_n46482_ & new_n46882_;
  assign new_n46884_ = ~new_n46483_ & ~new_n46486_;
  assign new_n46885_ = ~new_n46883_ & ~new_n46884_;
  assign new_n46886_ = ~new_n46636_ & ~new_n46885_;
  assign new_n46887_ = ~new_n46178_ & ~new_n46635_;
  assign new_n46888_ = ~new_n46634_ & new_n46887_;
  assign new_n46889_ = ~new_n46886_ & ~new_n46888_;
  assign new_n46890_ = ~\b[24]  & ~new_n46889_;
  assign new_n46891_ = ~new_n46197_ & new_n46481_;
  assign new_n46892_ = ~new_n46477_ & new_n46891_;
  assign new_n46893_ = ~new_n46478_ & ~new_n46481_;
  assign new_n46894_ = ~new_n46892_ & ~new_n46893_;
  assign new_n46895_ = ~new_n46636_ & ~new_n46894_;
  assign new_n46896_ = ~new_n46187_ & ~new_n46635_;
  assign new_n46897_ = ~new_n46634_ & new_n46896_;
  assign new_n46898_ = ~new_n46895_ & ~new_n46897_;
  assign new_n46899_ = ~\b[23]  & ~new_n46898_;
  assign new_n46900_ = ~new_n46206_ & new_n46476_;
  assign new_n46901_ = ~new_n46472_ & new_n46900_;
  assign new_n46902_ = ~new_n46473_ & ~new_n46476_;
  assign new_n46903_ = ~new_n46901_ & ~new_n46902_;
  assign new_n46904_ = ~new_n46636_ & ~new_n46903_;
  assign new_n46905_ = ~new_n46196_ & ~new_n46635_;
  assign new_n46906_ = ~new_n46634_ & new_n46905_;
  assign new_n46907_ = ~new_n46904_ & ~new_n46906_;
  assign new_n46908_ = ~\b[22]  & ~new_n46907_;
  assign new_n46909_ = ~new_n46215_ & new_n46471_;
  assign new_n46910_ = ~new_n46467_ & new_n46909_;
  assign new_n46911_ = ~new_n46468_ & ~new_n46471_;
  assign new_n46912_ = ~new_n46910_ & ~new_n46911_;
  assign new_n46913_ = ~new_n46636_ & ~new_n46912_;
  assign new_n46914_ = ~new_n46205_ & ~new_n46635_;
  assign new_n46915_ = ~new_n46634_ & new_n46914_;
  assign new_n46916_ = ~new_n46913_ & ~new_n46915_;
  assign new_n46917_ = ~\b[21]  & ~new_n46916_;
  assign new_n46918_ = ~new_n46224_ & new_n46466_;
  assign new_n46919_ = ~new_n46462_ & new_n46918_;
  assign new_n46920_ = ~new_n46463_ & ~new_n46466_;
  assign new_n46921_ = ~new_n46919_ & ~new_n46920_;
  assign new_n46922_ = ~new_n46636_ & ~new_n46921_;
  assign new_n46923_ = ~new_n46214_ & ~new_n46635_;
  assign new_n46924_ = ~new_n46634_ & new_n46923_;
  assign new_n46925_ = ~new_n46922_ & ~new_n46924_;
  assign new_n46926_ = ~\b[20]  & ~new_n46925_;
  assign new_n46927_ = ~new_n46233_ & new_n46461_;
  assign new_n46928_ = ~new_n46457_ & new_n46927_;
  assign new_n46929_ = ~new_n46458_ & ~new_n46461_;
  assign new_n46930_ = ~new_n46928_ & ~new_n46929_;
  assign new_n46931_ = ~new_n46636_ & ~new_n46930_;
  assign new_n46932_ = ~new_n46223_ & ~new_n46635_;
  assign new_n46933_ = ~new_n46634_ & new_n46932_;
  assign new_n46934_ = ~new_n46931_ & ~new_n46933_;
  assign new_n46935_ = ~\b[19]  & ~new_n46934_;
  assign new_n46936_ = ~new_n46242_ & new_n46456_;
  assign new_n46937_ = ~new_n46452_ & new_n46936_;
  assign new_n46938_ = ~new_n46453_ & ~new_n46456_;
  assign new_n46939_ = ~new_n46937_ & ~new_n46938_;
  assign new_n46940_ = ~new_n46636_ & ~new_n46939_;
  assign new_n46941_ = ~new_n46232_ & ~new_n46635_;
  assign new_n46942_ = ~new_n46634_ & new_n46941_;
  assign new_n46943_ = ~new_n46940_ & ~new_n46942_;
  assign new_n46944_ = ~\b[18]  & ~new_n46943_;
  assign new_n46945_ = ~new_n46251_ & new_n46451_;
  assign new_n46946_ = ~new_n46447_ & new_n46945_;
  assign new_n46947_ = ~new_n46448_ & ~new_n46451_;
  assign new_n46948_ = ~new_n46946_ & ~new_n46947_;
  assign new_n46949_ = ~new_n46636_ & ~new_n46948_;
  assign new_n46950_ = ~new_n46241_ & ~new_n46635_;
  assign new_n46951_ = ~new_n46634_ & new_n46950_;
  assign new_n46952_ = ~new_n46949_ & ~new_n46951_;
  assign new_n46953_ = ~\b[17]  & ~new_n46952_;
  assign new_n46954_ = ~new_n46260_ & new_n46446_;
  assign new_n46955_ = ~new_n46442_ & new_n46954_;
  assign new_n46956_ = ~new_n46443_ & ~new_n46446_;
  assign new_n46957_ = ~new_n46955_ & ~new_n46956_;
  assign new_n46958_ = ~new_n46636_ & ~new_n46957_;
  assign new_n46959_ = ~new_n46250_ & ~new_n46635_;
  assign new_n46960_ = ~new_n46634_ & new_n46959_;
  assign new_n46961_ = ~new_n46958_ & ~new_n46960_;
  assign new_n46962_ = ~\b[16]  & ~new_n46961_;
  assign new_n46963_ = ~new_n46269_ & new_n46441_;
  assign new_n46964_ = ~new_n46437_ & new_n46963_;
  assign new_n46965_ = ~new_n46438_ & ~new_n46441_;
  assign new_n46966_ = ~new_n46964_ & ~new_n46965_;
  assign new_n46967_ = ~new_n46636_ & ~new_n46966_;
  assign new_n46968_ = ~new_n46259_ & ~new_n46635_;
  assign new_n46969_ = ~new_n46634_ & new_n46968_;
  assign new_n46970_ = ~new_n46967_ & ~new_n46969_;
  assign new_n46971_ = ~\b[15]  & ~new_n46970_;
  assign new_n46972_ = ~new_n46278_ & new_n46436_;
  assign new_n46973_ = ~new_n46432_ & new_n46972_;
  assign new_n46974_ = ~new_n46433_ & ~new_n46436_;
  assign new_n46975_ = ~new_n46973_ & ~new_n46974_;
  assign new_n46976_ = ~new_n46636_ & ~new_n46975_;
  assign new_n46977_ = ~new_n46268_ & ~new_n46635_;
  assign new_n46978_ = ~new_n46634_ & new_n46977_;
  assign new_n46979_ = ~new_n46976_ & ~new_n46978_;
  assign new_n46980_ = ~\b[14]  & ~new_n46979_;
  assign new_n46981_ = ~new_n46287_ & new_n46431_;
  assign new_n46982_ = ~new_n46427_ & new_n46981_;
  assign new_n46983_ = ~new_n46428_ & ~new_n46431_;
  assign new_n46984_ = ~new_n46982_ & ~new_n46983_;
  assign new_n46985_ = ~new_n46636_ & ~new_n46984_;
  assign new_n46986_ = ~new_n46277_ & ~new_n46635_;
  assign new_n46987_ = ~new_n46634_ & new_n46986_;
  assign new_n46988_ = ~new_n46985_ & ~new_n46987_;
  assign new_n46989_ = ~\b[13]  & ~new_n46988_;
  assign new_n46990_ = ~new_n46296_ & new_n46426_;
  assign new_n46991_ = ~new_n46422_ & new_n46990_;
  assign new_n46992_ = ~new_n46423_ & ~new_n46426_;
  assign new_n46993_ = ~new_n46991_ & ~new_n46992_;
  assign new_n46994_ = ~new_n46636_ & ~new_n46993_;
  assign new_n46995_ = ~new_n46286_ & ~new_n46635_;
  assign new_n46996_ = ~new_n46634_ & new_n46995_;
  assign new_n46997_ = ~new_n46994_ & ~new_n46996_;
  assign new_n46998_ = ~\b[12]  & ~new_n46997_;
  assign new_n46999_ = ~new_n46305_ & new_n46421_;
  assign new_n47000_ = ~new_n46417_ & new_n46999_;
  assign new_n47001_ = ~new_n46418_ & ~new_n46421_;
  assign new_n47002_ = ~new_n47000_ & ~new_n47001_;
  assign new_n47003_ = ~new_n46636_ & ~new_n47002_;
  assign new_n47004_ = ~new_n46295_ & ~new_n46635_;
  assign new_n47005_ = ~new_n46634_ & new_n47004_;
  assign new_n47006_ = ~new_n47003_ & ~new_n47005_;
  assign new_n47007_ = ~\b[11]  & ~new_n47006_;
  assign new_n47008_ = ~new_n46314_ & new_n46416_;
  assign new_n47009_ = ~new_n46412_ & new_n47008_;
  assign new_n47010_ = ~new_n46413_ & ~new_n46416_;
  assign new_n47011_ = ~new_n47009_ & ~new_n47010_;
  assign new_n47012_ = ~new_n46636_ & ~new_n47011_;
  assign new_n47013_ = ~new_n46304_ & ~new_n46635_;
  assign new_n47014_ = ~new_n46634_ & new_n47013_;
  assign new_n47015_ = ~new_n47012_ & ~new_n47014_;
  assign new_n47016_ = ~\b[10]  & ~new_n47015_;
  assign new_n47017_ = ~new_n46323_ & new_n46411_;
  assign new_n47018_ = ~new_n46407_ & new_n47017_;
  assign new_n47019_ = ~new_n46408_ & ~new_n46411_;
  assign new_n47020_ = ~new_n47018_ & ~new_n47019_;
  assign new_n47021_ = ~new_n46636_ & ~new_n47020_;
  assign new_n47022_ = ~new_n46313_ & ~new_n46635_;
  assign new_n47023_ = ~new_n46634_ & new_n47022_;
  assign new_n47024_ = ~new_n47021_ & ~new_n47023_;
  assign new_n47025_ = ~\b[9]  & ~new_n47024_;
  assign new_n47026_ = ~new_n46332_ & new_n46406_;
  assign new_n47027_ = ~new_n46402_ & new_n47026_;
  assign new_n47028_ = ~new_n46403_ & ~new_n46406_;
  assign new_n47029_ = ~new_n47027_ & ~new_n47028_;
  assign new_n47030_ = ~new_n46636_ & ~new_n47029_;
  assign new_n47031_ = ~new_n46322_ & ~new_n46635_;
  assign new_n47032_ = ~new_n46634_ & new_n47031_;
  assign new_n47033_ = ~new_n47030_ & ~new_n47032_;
  assign new_n47034_ = ~\b[8]  & ~new_n47033_;
  assign new_n47035_ = ~new_n46341_ & new_n46401_;
  assign new_n47036_ = ~new_n46397_ & new_n47035_;
  assign new_n47037_ = ~new_n46398_ & ~new_n46401_;
  assign new_n47038_ = ~new_n47036_ & ~new_n47037_;
  assign new_n47039_ = ~new_n46636_ & ~new_n47038_;
  assign new_n47040_ = ~new_n46331_ & ~new_n46635_;
  assign new_n47041_ = ~new_n46634_ & new_n47040_;
  assign new_n47042_ = ~new_n47039_ & ~new_n47041_;
  assign new_n47043_ = ~\b[7]  & ~new_n47042_;
  assign new_n47044_ = ~new_n46350_ & new_n46396_;
  assign new_n47045_ = ~new_n46392_ & new_n47044_;
  assign new_n47046_ = ~new_n46393_ & ~new_n46396_;
  assign new_n47047_ = ~new_n47045_ & ~new_n47046_;
  assign new_n47048_ = ~new_n46636_ & ~new_n47047_;
  assign new_n47049_ = ~new_n46340_ & ~new_n46635_;
  assign new_n47050_ = ~new_n46634_ & new_n47049_;
  assign new_n47051_ = ~new_n47048_ & ~new_n47050_;
  assign new_n47052_ = ~\b[6]  & ~new_n47051_;
  assign new_n47053_ = ~new_n46359_ & new_n46391_;
  assign new_n47054_ = ~new_n46387_ & new_n47053_;
  assign new_n47055_ = ~new_n46388_ & ~new_n46391_;
  assign new_n47056_ = ~new_n47054_ & ~new_n47055_;
  assign new_n47057_ = ~new_n46636_ & ~new_n47056_;
  assign new_n47058_ = ~new_n46349_ & ~new_n46635_;
  assign new_n47059_ = ~new_n46634_ & new_n47058_;
  assign new_n47060_ = ~new_n47057_ & ~new_n47059_;
  assign new_n47061_ = ~\b[5]  & ~new_n47060_;
  assign new_n47062_ = ~new_n46367_ & new_n46386_;
  assign new_n47063_ = ~new_n46382_ & new_n47062_;
  assign new_n47064_ = ~new_n46383_ & ~new_n46386_;
  assign new_n47065_ = ~new_n47063_ & ~new_n47064_;
  assign new_n47066_ = ~new_n46636_ & ~new_n47065_;
  assign new_n47067_ = ~new_n46358_ & ~new_n46635_;
  assign new_n47068_ = ~new_n46634_ & new_n47067_;
  assign new_n47069_ = ~new_n47066_ & ~new_n47068_;
  assign new_n47070_ = ~\b[4]  & ~new_n47069_;
  assign new_n47071_ = ~new_n46377_ & new_n46381_;
  assign new_n47072_ = ~new_n46376_ & new_n47071_;
  assign new_n47073_ = ~new_n46378_ & ~new_n46381_;
  assign new_n47074_ = ~new_n47072_ & ~new_n47073_;
  assign new_n47075_ = ~new_n46636_ & ~new_n47074_;
  assign new_n47076_ = ~new_n46366_ & ~new_n46635_;
  assign new_n47077_ = ~new_n46634_ & new_n47076_;
  assign new_n47078_ = ~new_n47075_ & ~new_n47077_;
  assign new_n47079_ = ~\b[3]  & ~new_n47078_;
  assign new_n47080_ = new_n18327_ & ~new_n46374_;
  assign new_n47081_ = ~new_n46372_ & new_n47080_;
  assign new_n47082_ = ~new_n46376_ & ~new_n47081_;
  assign new_n47083_ = ~new_n46636_ & new_n47082_;
  assign new_n47084_ = ~new_n46371_ & ~new_n46635_;
  assign new_n47085_ = ~new_n46634_ & new_n47084_;
  assign new_n47086_ = ~new_n47083_ & ~new_n47085_;
  assign new_n47087_ = ~\b[2]  & ~new_n47086_;
  assign new_n47088_ = \b[0]  & ~new_n46636_;
  assign new_n47089_ = \a[13]  & ~new_n47088_;
  assign new_n47090_ = new_n18327_ & ~new_n46636_;
  assign new_n47091_ = ~new_n47089_ & ~new_n47090_;
  assign new_n47092_ = \b[1]  & ~new_n47091_;
  assign new_n47093_ = ~\b[1]  & ~new_n47090_;
  assign new_n47094_ = ~new_n47089_ & new_n47093_;
  assign new_n47095_ = ~new_n47092_ & ~new_n47094_;
  assign new_n47096_ = ~new_n19050_ & ~new_n47095_;
  assign new_n47097_ = ~\b[1]  & ~new_n47091_;
  assign new_n47098_ = ~new_n47096_ & ~new_n47097_;
  assign new_n47099_ = \b[2]  & ~new_n47085_;
  assign new_n47100_ = ~new_n47083_ & new_n47099_;
  assign new_n47101_ = ~new_n47087_ & ~new_n47100_;
  assign new_n47102_ = ~new_n47098_ & new_n47101_;
  assign new_n47103_ = ~new_n47087_ & ~new_n47102_;
  assign new_n47104_ = \b[3]  & ~new_n47077_;
  assign new_n47105_ = ~new_n47075_ & new_n47104_;
  assign new_n47106_ = ~new_n47079_ & ~new_n47105_;
  assign new_n47107_ = ~new_n47103_ & new_n47106_;
  assign new_n47108_ = ~new_n47079_ & ~new_n47107_;
  assign new_n47109_ = \b[4]  & ~new_n47068_;
  assign new_n47110_ = ~new_n47066_ & new_n47109_;
  assign new_n47111_ = ~new_n47070_ & ~new_n47110_;
  assign new_n47112_ = ~new_n47108_ & new_n47111_;
  assign new_n47113_ = ~new_n47070_ & ~new_n47112_;
  assign new_n47114_ = \b[5]  & ~new_n47059_;
  assign new_n47115_ = ~new_n47057_ & new_n47114_;
  assign new_n47116_ = ~new_n47061_ & ~new_n47115_;
  assign new_n47117_ = ~new_n47113_ & new_n47116_;
  assign new_n47118_ = ~new_n47061_ & ~new_n47117_;
  assign new_n47119_ = \b[6]  & ~new_n47050_;
  assign new_n47120_ = ~new_n47048_ & new_n47119_;
  assign new_n47121_ = ~new_n47052_ & ~new_n47120_;
  assign new_n47122_ = ~new_n47118_ & new_n47121_;
  assign new_n47123_ = ~new_n47052_ & ~new_n47122_;
  assign new_n47124_ = \b[7]  & ~new_n47041_;
  assign new_n47125_ = ~new_n47039_ & new_n47124_;
  assign new_n47126_ = ~new_n47043_ & ~new_n47125_;
  assign new_n47127_ = ~new_n47123_ & new_n47126_;
  assign new_n47128_ = ~new_n47043_ & ~new_n47127_;
  assign new_n47129_ = \b[8]  & ~new_n47032_;
  assign new_n47130_ = ~new_n47030_ & new_n47129_;
  assign new_n47131_ = ~new_n47034_ & ~new_n47130_;
  assign new_n47132_ = ~new_n47128_ & new_n47131_;
  assign new_n47133_ = ~new_n47034_ & ~new_n47132_;
  assign new_n47134_ = \b[9]  & ~new_n47023_;
  assign new_n47135_ = ~new_n47021_ & new_n47134_;
  assign new_n47136_ = ~new_n47025_ & ~new_n47135_;
  assign new_n47137_ = ~new_n47133_ & new_n47136_;
  assign new_n47138_ = ~new_n47025_ & ~new_n47137_;
  assign new_n47139_ = \b[10]  & ~new_n47014_;
  assign new_n47140_ = ~new_n47012_ & new_n47139_;
  assign new_n47141_ = ~new_n47016_ & ~new_n47140_;
  assign new_n47142_ = ~new_n47138_ & new_n47141_;
  assign new_n47143_ = ~new_n47016_ & ~new_n47142_;
  assign new_n47144_ = \b[11]  & ~new_n47005_;
  assign new_n47145_ = ~new_n47003_ & new_n47144_;
  assign new_n47146_ = ~new_n47007_ & ~new_n47145_;
  assign new_n47147_ = ~new_n47143_ & new_n47146_;
  assign new_n47148_ = ~new_n47007_ & ~new_n47147_;
  assign new_n47149_ = \b[12]  & ~new_n46996_;
  assign new_n47150_ = ~new_n46994_ & new_n47149_;
  assign new_n47151_ = ~new_n46998_ & ~new_n47150_;
  assign new_n47152_ = ~new_n47148_ & new_n47151_;
  assign new_n47153_ = ~new_n46998_ & ~new_n47152_;
  assign new_n47154_ = \b[13]  & ~new_n46987_;
  assign new_n47155_ = ~new_n46985_ & new_n47154_;
  assign new_n47156_ = ~new_n46989_ & ~new_n47155_;
  assign new_n47157_ = ~new_n47153_ & new_n47156_;
  assign new_n47158_ = ~new_n46989_ & ~new_n47157_;
  assign new_n47159_ = \b[14]  & ~new_n46978_;
  assign new_n47160_ = ~new_n46976_ & new_n47159_;
  assign new_n47161_ = ~new_n46980_ & ~new_n47160_;
  assign new_n47162_ = ~new_n47158_ & new_n47161_;
  assign new_n47163_ = ~new_n46980_ & ~new_n47162_;
  assign new_n47164_ = \b[15]  & ~new_n46969_;
  assign new_n47165_ = ~new_n46967_ & new_n47164_;
  assign new_n47166_ = ~new_n46971_ & ~new_n47165_;
  assign new_n47167_ = ~new_n47163_ & new_n47166_;
  assign new_n47168_ = ~new_n46971_ & ~new_n47167_;
  assign new_n47169_ = \b[16]  & ~new_n46960_;
  assign new_n47170_ = ~new_n46958_ & new_n47169_;
  assign new_n47171_ = ~new_n46962_ & ~new_n47170_;
  assign new_n47172_ = ~new_n47168_ & new_n47171_;
  assign new_n47173_ = ~new_n46962_ & ~new_n47172_;
  assign new_n47174_ = \b[17]  & ~new_n46951_;
  assign new_n47175_ = ~new_n46949_ & new_n47174_;
  assign new_n47176_ = ~new_n46953_ & ~new_n47175_;
  assign new_n47177_ = ~new_n47173_ & new_n47176_;
  assign new_n47178_ = ~new_n46953_ & ~new_n47177_;
  assign new_n47179_ = \b[18]  & ~new_n46942_;
  assign new_n47180_ = ~new_n46940_ & new_n47179_;
  assign new_n47181_ = ~new_n46944_ & ~new_n47180_;
  assign new_n47182_ = ~new_n47178_ & new_n47181_;
  assign new_n47183_ = ~new_n46944_ & ~new_n47182_;
  assign new_n47184_ = \b[19]  & ~new_n46933_;
  assign new_n47185_ = ~new_n46931_ & new_n47184_;
  assign new_n47186_ = ~new_n46935_ & ~new_n47185_;
  assign new_n47187_ = ~new_n47183_ & new_n47186_;
  assign new_n47188_ = ~new_n46935_ & ~new_n47187_;
  assign new_n47189_ = \b[20]  & ~new_n46924_;
  assign new_n47190_ = ~new_n46922_ & new_n47189_;
  assign new_n47191_ = ~new_n46926_ & ~new_n47190_;
  assign new_n47192_ = ~new_n47188_ & new_n47191_;
  assign new_n47193_ = ~new_n46926_ & ~new_n47192_;
  assign new_n47194_ = \b[21]  & ~new_n46915_;
  assign new_n47195_ = ~new_n46913_ & new_n47194_;
  assign new_n47196_ = ~new_n46917_ & ~new_n47195_;
  assign new_n47197_ = ~new_n47193_ & new_n47196_;
  assign new_n47198_ = ~new_n46917_ & ~new_n47197_;
  assign new_n47199_ = \b[22]  & ~new_n46906_;
  assign new_n47200_ = ~new_n46904_ & new_n47199_;
  assign new_n47201_ = ~new_n46908_ & ~new_n47200_;
  assign new_n47202_ = ~new_n47198_ & new_n47201_;
  assign new_n47203_ = ~new_n46908_ & ~new_n47202_;
  assign new_n47204_ = \b[23]  & ~new_n46897_;
  assign new_n47205_ = ~new_n46895_ & new_n47204_;
  assign new_n47206_ = ~new_n46899_ & ~new_n47205_;
  assign new_n47207_ = ~new_n47203_ & new_n47206_;
  assign new_n47208_ = ~new_n46899_ & ~new_n47207_;
  assign new_n47209_ = \b[24]  & ~new_n46888_;
  assign new_n47210_ = ~new_n46886_ & new_n47209_;
  assign new_n47211_ = ~new_n46890_ & ~new_n47210_;
  assign new_n47212_ = ~new_n47208_ & new_n47211_;
  assign new_n47213_ = ~new_n46890_ & ~new_n47212_;
  assign new_n47214_ = \b[25]  & ~new_n46879_;
  assign new_n47215_ = ~new_n46877_ & new_n47214_;
  assign new_n47216_ = ~new_n46881_ & ~new_n47215_;
  assign new_n47217_ = ~new_n47213_ & new_n47216_;
  assign new_n47218_ = ~new_n46881_ & ~new_n47217_;
  assign new_n47219_ = \b[26]  & ~new_n46870_;
  assign new_n47220_ = ~new_n46868_ & new_n47219_;
  assign new_n47221_ = ~new_n46872_ & ~new_n47220_;
  assign new_n47222_ = ~new_n47218_ & new_n47221_;
  assign new_n47223_ = ~new_n46872_ & ~new_n47222_;
  assign new_n47224_ = \b[27]  & ~new_n46861_;
  assign new_n47225_ = ~new_n46859_ & new_n47224_;
  assign new_n47226_ = ~new_n46863_ & ~new_n47225_;
  assign new_n47227_ = ~new_n47223_ & new_n47226_;
  assign new_n47228_ = ~new_n46863_ & ~new_n47227_;
  assign new_n47229_ = \b[28]  & ~new_n46852_;
  assign new_n47230_ = ~new_n46850_ & new_n47229_;
  assign new_n47231_ = ~new_n46854_ & ~new_n47230_;
  assign new_n47232_ = ~new_n47228_ & new_n47231_;
  assign new_n47233_ = ~new_n46854_ & ~new_n47232_;
  assign new_n47234_ = \b[29]  & ~new_n46843_;
  assign new_n47235_ = ~new_n46841_ & new_n47234_;
  assign new_n47236_ = ~new_n46845_ & ~new_n47235_;
  assign new_n47237_ = ~new_n47233_ & new_n47236_;
  assign new_n47238_ = ~new_n46845_ & ~new_n47237_;
  assign new_n47239_ = \b[30]  & ~new_n46834_;
  assign new_n47240_ = ~new_n46832_ & new_n47239_;
  assign new_n47241_ = ~new_n46836_ & ~new_n47240_;
  assign new_n47242_ = ~new_n47238_ & new_n47241_;
  assign new_n47243_ = ~new_n46836_ & ~new_n47242_;
  assign new_n47244_ = \b[31]  & ~new_n46825_;
  assign new_n47245_ = ~new_n46823_ & new_n47244_;
  assign new_n47246_ = ~new_n46827_ & ~new_n47245_;
  assign new_n47247_ = ~new_n47243_ & new_n47246_;
  assign new_n47248_ = ~new_n46827_ & ~new_n47247_;
  assign new_n47249_ = \b[32]  & ~new_n46816_;
  assign new_n47250_ = ~new_n46814_ & new_n47249_;
  assign new_n47251_ = ~new_n46818_ & ~new_n47250_;
  assign new_n47252_ = ~new_n47248_ & new_n47251_;
  assign new_n47253_ = ~new_n46818_ & ~new_n47252_;
  assign new_n47254_ = \b[33]  & ~new_n46807_;
  assign new_n47255_ = ~new_n46805_ & new_n47254_;
  assign new_n47256_ = ~new_n46809_ & ~new_n47255_;
  assign new_n47257_ = ~new_n47253_ & new_n47256_;
  assign new_n47258_ = ~new_n46809_ & ~new_n47257_;
  assign new_n47259_ = \b[34]  & ~new_n46798_;
  assign new_n47260_ = ~new_n46796_ & new_n47259_;
  assign new_n47261_ = ~new_n46800_ & ~new_n47260_;
  assign new_n47262_ = ~new_n47258_ & new_n47261_;
  assign new_n47263_ = ~new_n46800_ & ~new_n47262_;
  assign new_n47264_ = \b[35]  & ~new_n46789_;
  assign new_n47265_ = ~new_n46787_ & new_n47264_;
  assign new_n47266_ = ~new_n46791_ & ~new_n47265_;
  assign new_n47267_ = ~new_n47263_ & new_n47266_;
  assign new_n47268_ = ~new_n46791_ & ~new_n47267_;
  assign new_n47269_ = \b[36]  & ~new_n46780_;
  assign new_n47270_ = ~new_n46778_ & new_n47269_;
  assign new_n47271_ = ~new_n46782_ & ~new_n47270_;
  assign new_n47272_ = ~new_n47268_ & new_n47271_;
  assign new_n47273_ = ~new_n46782_ & ~new_n47272_;
  assign new_n47274_ = \b[37]  & ~new_n46771_;
  assign new_n47275_ = ~new_n46769_ & new_n47274_;
  assign new_n47276_ = ~new_n46773_ & ~new_n47275_;
  assign new_n47277_ = ~new_n47273_ & new_n47276_;
  assign new_n47278_ = ~new_n46773_ & ~new_n47277_;
  assign new_n47279_ = \b[38]  & ~new_n46762_;
  assign new_n47280_ = ~new_n46760_ & new_n47279_;
  assign new_n47281_ = ~new_n46764_ & ~new_n47280_;
  assign new_n47282_ = ~new_n47278_ & new_n47281_;
  assign new_n47283_ = ~new_n46764_ & ~new_n47282_;
  assign new_n47284_ = \b[39]  & ~new_n46753_;
  assign new_n47285_ = ~new_n46751_ & new_n47284_;
  assign new_n47286_ = ~new_n46755_ & ~new_n47285_;
  assign new_n47287_ = ~new_n47283_ & new_n47286_;
  assign new_n47288_ = ~new_n46755_ & ~new_n47287_;
  assign new_n47289_ = \b[40]  & ~new_n46744_;
  assign new_n47290_ = ~new_n46742_ & new_n47289_;
  assign new_n47291_ = ~new_n46746_ & ~new_n47290_;
  assign new_n47292_ = ~new_n47288_ & new_n47291_;
  assign new_n47293_ = ~new_n46746_ & ~new_n47292_;
  assign new_n47294_ = \b[41]  & ~new_n46735_;
  assign new_n47295_ = ~new_n46733_ & new_n47294_;
  assign new_n47296_ = ~new_n46737_ & ~new_n47295_;
  assign new_n47297_ = ~new_n47293_ & new_n47296_;
  assign new_n47298_ = ~new_n46737_ & ~new_n47297_;
  assign new_n47299_ = \b[42]  & ~new_n46726_;
  assign new_n47300_ = ~new_n46724_ & new_n47299_;
  assign new_n47301_ = ~new_n46728_ & ~new_n47300_;
  assign new_n47302_ = ~new_n47298_ & new_n47301_;
  assign new_n47303_ = ~new_n46728_ & ~new_n47302_;
  assign new_n47304_ = \b[43]  & ~new_n46717_;
  assign new_n47305_ = ~new_n46715_ & new_n47304_;
  assign new_n47306_ = ~new_n46719_ & ~new_n47305_;
  assign new_n47307_ = ~new_n47303_ & new_n47306_;
  assign new_n47308_ = ~new_n46719_ & ~new_n47307_;
  assign new_n47309_ = \b[44]  & ~new_n46708_;
  assign new_n47310_ = ~new_n46706_ & new_n47309_;
  assign new_n47311_ = ~new_n46710_ & ~new_n47310_;
  assign new_n47312_ = ~new_n47308_ & new_n47311_;
  assign new_n47313_ = ~new_n46710_ & ~new_n47312_;
  assign new_n47314_ = \b[45]  & ~new_n46699_;
  assign new_n47315_ = ~new_n46697_ & new_n47314_;
  assign new_n47316_ = ~new_n46701_ & ~new_n47315_;
  assign new_n47317_ = ~new_n47313_ & new_n47316_;
  assign new_n47318_ = ~new_n46701_ & ~new_n47317_;
  assign new_n47319_ = \b[46]  & ~new_n46690_;
  assign new_n47320_ = ~new_n46688_ & new_n47319_;
  assign new_n47321_ = ~new_n46692_ & ~new_n47320_;
  assign new_n47322_ = ~new_n47318_ & new_n47321_;
  assign new_n47323_ = ~new_n46692_ & ~new_n47322_;
  assign new_n47324_ = \b[47]  & ~new_n46681_;
  assign new_n47325_ = ~new_n46679_ & new_n47324_;
  assign new_n47326_ = ~new_n46683_ & ~new_n47325_;
  assign new_n47327_ = ~new_n47323_ & new_n47326_;
  assign new_n47328_ = ~new_n46683_ & ~new_n47327_;
  assign new_n47329_ = \b[48]  & ~new_n46672_;
  assign new_n47330_ = ~new_n46670_ & new_n47329_;
  assign new_n47331_ = ~new_n46674_ & ~new_n47330_;
  assign new_n47332_ = ~new_n47328_ & new_n47331_;
  assign new_n47333_ = ~new_n46674_ & ~new_n47332_;
  assign new_n47334_ = \b[49]  & ~new_n46663_;
  assign new_n47335_ = ~new_n46661_ & new_n47334_;
  assign new_n47336_ = ~new_n46665_ & ~new_n47335_;
  assign new_n47337_ = ~new_n47333_ & new_n47336_;
  assign new_n47338_ = ~new_n46665_ & ~new_n47337_;
  assign new_n47339_ = \b[50]  & ~new_n46643_;
  assign new_n47340_ = ~new_n46641_ & new_n47339_;
  assign new_n47341_ = ~new_n46656_ & ~new_n47340_;
  assign new_n47342_ = ~new_n47338_ & new_n47341_;
  assign new_n47343_ = ~new_n46656_ & ~new_n47342_;
  assign new_n47344_ = \b[51]  & ~new_n46653_;
  assign new_n47345_ = ~new_n46651_ & new_n47344_;
  assign new_n47346_ = ~new_n46655_ & ~new_n47345_;
  assign new_n47347_ = ~new_n47343_ & new_n47346_;
  assign new_n47348_ = ~new_n46655_ & ~new_n47347_;
  assign new_n47349_ = new_n288_ & ~new_n47348_;
  assign new_n47350_ = ~new_n46644_ & ~new_n47349_;
  assign new_n47351_ = ~new_n46665_ & new_n47341_;
  assign new_n47352_ = ~new_n47337_ & new_n47351_;
  assign new_n47353_ = ~new_n47338_ & ~new_n47341_;
  assign new_n47354_ = ~new_n47352_ & ~new_n47353_;
  assign new_n47355_ = new_n288_ & ~new_n47354_;
  assign new_n47356_ = ~new_n47348_ & new_n47355_;
  assign new_n47357_ = ~new_n47350_ & ~new_n47356_;
  assign new_n47358_ = ~\b[51]  & ~new_n47357_;
  assign new_n47359_ = ~new_n46664_ & ~new_n47349_;
  assign new_n47360_ = ~new_n46674_ & new_n47336_;
  assign new_n47361_ = ~new_n47332_ & new_n47360_;
  assign new_n47362_ = ~new_n47333_ & ~new_n47336_;
  assign new_n47363_ = ~new_n47361_ & ~new_n47362_;
  assign new_n47364_ = new_n288_ & ~new_n47363_;
  assign new_n47365_ = ~new_n47348_ & new_n47364_;
  assign new_n47366_ = ~new_n47359_ & ~new_n47365_;
  assign new_n47367_ = ~\b[50]  & ~new_n47366_;
  assign new_n47368_ = ~new_n46673_ & ~new_n47349_;
  assign new_n47369_ = ~new_n46683_ & new_n47331_;
  assign new_n47370_ = ~new_n47327_ & new_n47369_;
  assign new_n47371_ = ~new_n47328_ & ~new_n47331_;
  assign new_n47372_ = ~new_n47370_ & ~new_n47371_;
  assign new_n47373_ = new_n288_ & ~new_n47372_;
  assign new_n47374_ = ~new_n47348_ & new_n47373_;
  assign new_n47375_ = ~new_n47368_ & ~new_n47374_;
  assign new_n47376_ = ~\b[49]  & ~new_n47375_;
  assign new_n47377_ = ~new_n46682_ & ~new_n47349_;
  assign new_n47378_ = ~new_n46692_ & new_n47326_;
  assign new_n47379_ = ~new_n47322_ & new_n47378_;
  assign new_n47380_ = ~new_n47323_ & ~new_n47326_;
  assign new_n47381_ = ~new_n47379_ & ~new_n47380_;
  assign new_n47382_ = new_n288_ & ~new_n47381_;
  assign new_n47383_ = ~new_n47348_ & new_n47382_;
  assign new_n47384_ = ~new_n47377_ & ~new_n47383_;
  assign new_n47385_ = ~\b[48]  & ~new_n47384_;
  assign new_n47386_ = ~new_n46691_ & ~new_n47349_;
  assign new_n47387_ = ~new_n46701_ & new_n47321_;
  assign new_n47388_ = ~new_n47317_ & new_n47387_;
  assign new_n47389_ = ~new_n47318_ & ~new_n47321_;
  assign new_n47390_ = ~new_n47388_ & ~new_n47389_;
  assign new_n47391_ = new_n288_ & ~new_n47390_;
  assign new_n47392_ = ~new_n47348_ & new_n47391_;
  assign new_n47393_ = ~new_n47386_ & ~new_n47392_;
  assign new_n47394_ = ~\b[47]  & ~new_n47393_;
  assign new_n47395_ = ~new_n46700_ & ~new_n47349_;
  assign new_n47396_ = ~new_n46710_ & new_n47316_;
  assign new_n47397_ = ~new_n47312_ & new_n47396_;
  assign new_n47398_ = ~new_n47313_ & ~new_n47316_;
  assign new_n47399_ = ~new_n47397_ & ~new_n47398_;
  assign new_n47400_ = new_n288_ & ~new_n47399_;
  assign new_n47401_ = ~new_n47348_ & new_n47400_;
  assign new_n47402_ = ~new_n47395_ & ~new_n47401_;
  assign new_n47403_ = ~\b[46]  & ~new_n47402_;
  assign new_n47404_ = ~new_n46709_ & ~new_n47349_;
  assign new_n47405_ = ~new_n46719_ & new_n47311_;
  assign new_n47406_ = ~new_n47307_ & new_n47405_;
  assign new_n47407_ = ~new_n47308_ & ~new_n47311_;
  assign new_n47408_ = ~new_n47406_ & ~new_n47407_;
  assign new_n47409_ = new_n288_ & ~new_n47408_;
  assign new_n47410_ = ~new_n47348_ & new_n47409_;
  assign new_n47411_ = ~new_n47404_ & ~new_n47410_;
  assign new_n47412_ = ~\b[45]  & ~new_n47411_;
  assign new_n47413_ = ~new_n46718_ & ~new_n47349_;
  assign new_n47414_ = ~new_n46728_ & new_n47306_;
  assign new_n47415_ = ~new_n47302_ & new_n47414_;
  assign new_n47416_ = ~new_n47303_ & ~new_n47306_;
  assign new_n47417_ = ~new_n47415_ & ~new_n47416_;
  assign new_n47418_ = new_n288_ & ~new_n47417_;
  assign new_n47419_ = ~new_n47348_ & new_n47418_;
  assign new_n47420_ = ~new_n47413_ & ~new_n47419_;
  assign new_n47421_ = ~\b[44]  & ~new_n47420_;
  assign new_n47422_ = ~new_n46727_ & ~new_n47349_;
  assign new_n47423_ = ~new_n46737_ & new_n47301_;
  assign new_n47424_ = ~new_n47297_ & new_n47423_;
  assign new_n47425_ = ~new_n47298_ & ~new_n47301_;
  assign new_n47426_ = ~new_n47424_ & ~new_n47425_;
  assign new_n47427_ = new_n288_ & ~new_n47426_;
  assign new_n47428_ = ~new_n47348_ & new_n47427_;
  assign new_n47429_ = ~new_n47422_ & ~new_n47428_;
  assign new_n47430_ = ~\b[43]  & ~new_n47429_;
  assign new_n47431_ = ~new_n46736_ & ~new_n47349_;
  assign new_n47432_ = ~new_n46746_ & new_n47296_;
  assign new_n47433_ = ~new_n47292_ & new_n47432_;
  assign new_n47434_ = ~new_n47293_ & ~new_n47296_;
  assign new_n47435_ = ~new_n47433_ & ~new_n47434_;
  assign new_n47436_ = new_n288_ & ~new_n47435_;
  assign new_n47437_ = ~new_n47348_ & new_n47436_;
  assign new_n47438_ = ~new_n47431_ & ~new_n47437_;
  assign new_n47439_ = ~\b[42]  & ~new_n47438_;
  assign new_n47440_ = ~new_n46745_ & ~new_n47349_;
  assign new_n47441_ = ~new_n46755_ & new_n47291_;
  assign new_n47442_ = ~new_n47287_ & new_n47441_;
  assign new_n47443_ = ~new_n47288_ & ~new_n47291_;
  assign new_n47444_ = ~new_n47442_ & ~new_n47443_;
  assign new_n47445_ = new_n288_ & ~new_n47444_;
  assign new_n47446_ = ~new_n47348_ & new_n47445_;
  assign new_n47447_ = ~new_n47440_ & ~new_n47446_;
  assign new_n47448_ = ~\b[41]  & ~new_n47447_;
  assign new_n47449_ = ~new_n46754_ & ~new_n47349_;
  assign new_n47450_ = ~new_n46764_ & new_n47286_;
  assign new_n47451_ = ~new_n47282_ & new_n47450_;
  assign new_n47452_ = ~new_n47283_ & ~new_n47286_;
  assign new_n47453_ = ~new_n47451_ & ~new_n47452_;
  assign new_n47454_ = new_n288_ & ~new_n47453_;
  assign new_n47455_ = ~new_n47348_ & new_n47454_;
  assign new_n47456_ = ~new_n47449_ & ~new_n47455_;
  assign new_n47457_ = ~\b[40]  & ~new_n47456_;
  assign new_n47458_ = ~new_n46763_ & ~new_n47349_;
  assign new_n47459_ = ~new_n46773_ & new_n47281_;
  assign new_n47460_ = ~new_n47277_ & new_n47459_;
  assign new_n47461_ = ~new_n47278_ & ~new_n47281_;
  assign new_n47462_ = ~new_n47460_ & ~new_n47461_;
  assign new_n47463_ = new_n288_ & ~new_n47462_;
  assign new_n47464_ = ~new_n47348_ & new_n47463_;
  assign new_n47465_ = ~new_n47458_ & ~new_n47464_;
  assign new_n47466_ = ~\b[39]  & ~new_n47465_;
  assign new_n47467_ = ~new_n46772_ & ~new_n47349_;
  assign new_n47468_ = ~new_n46782_ & new_n47276_;
  assign new_n47469_ = ~new_n47272_ & new_n47468_;
  assign new_n47470_ = ~new_n47273_ & ~new_n47276_;
  assign new_n47471_ = ~new_n47469_ & ~new_n47470_;
  assign new_n47472_ = new_n288_ & ~new_n47471_;
  assign new_n47473_ = ~new_n47348_ & new_n47472_;
  assign new_n47474_ = ~new_n47467_ & ~new_n47473_;
  assign new_n47475_ = ~\b[38]  & ~new_n47474_;
  assign new_n47476_ = ~new_n46781_ & ~new_n47349_;
  assign new_n47477_ = ~new_n46791_ & new_n47271_;
  assign new_n47478_ = ~new_n47267_ & new_n47477_;
  assign new_n47479_ = ~new_n47268_ & ~new_n47271_;
  assign new_n47480_ = ~new_n47478_ & ~new_n47479_;
  assign new_n47481_ = new_n288_ & ~new_n47480_;
  assign new_n47482_ = ~new_n47348_ & new_n47481_;
  assign new_n47483_ = ~new_n47476_ & ~new_n47482_;
  assign new_n47484_ = ~\b[37]  & ~new_n47483_;
  assign new_n47485_ = ~new_n46790_ & ~new_n47349_;
  assign new_n47486_ = ~new_n46800_ & new_n47266_;
  assign new_n47487_ = ~new_n47262_ & new_n47486_;
  assign new_n47488_ = ~new_n47263_ & ~new_n47266_;
  assign new_n47489_ = ~new_n47487_ & ~new_n47488_;
  assign new_n47490_ = new_n288_ & ~new_n47489_;
  assign new_n47491_ = ~new_n47348_ & new_n47490_;
  assign new_n47492_ = ~new_n47485_ & ~new_n47491_;
  assign new_n47493_ = ~\b[36]  & ~new_n47492_;
  assign new_n47494_ = ~new_n46799_ & ~new_n47349_;
  assign new_n47495_ = ~new_n46809_ & new_n47261_;
  assign new_n47496_ = ~new_n47257_ & new_n47495_;
  assign new_n47497_ = ~new_n47258_ & ~new_n47261_;
  assign new_n47498_ = ~new_n47496_ & ~new_n47497_;
  assign new_n47499_ = new_n288_ & ~new_n47498_;
  assign new_n47500_ = ~new_n47348_ & new_n47499_;
  assign new_n47501_ = ~new_n47494_ & ~new_n47500_;
  assign new_n47502_ = ~\b[35]  & ~new_n47501_;
  assign new_n47503_ = ~new_n46808_ & ~new_n47349_;
  assign new_n47504_ = ~new_n46818_ & new_n47256_;
  assign new_n47505_ = ~new_n47252_ & new_n47504_;
  assign new_n47506_ = ~new_n47253_ & ~new_n47256_;
  assign new_n47507_ = ~new_n47505_ & ~new_n47506_;
  assign new_n47508_ = new_n288_ & ~new_n47507_;
  assign new_n47509_ = ~new_n47348_ & new_n47508_;
  assign new_n47510_ = ~new_n47503_ & ~new_n47509_;
  assign new_n47511_ = ~\b[34]  & ~new_n47510_;
  assign new_n47512_ = ~new_n46817_ & ~new_n47349_;
  assign new_n47513_ = ~new_n46827_ & new_n47251_;
  assign new_n47514_ = ~new_n47247_ & new_n47513_;
  assign new_n47515_ = ~new_n47248_ & ~new_n47251_;
  assign new_n47516_ = ~new_n47514_ & ~new_n47515_;
  assign new_n47517_ = new_n288_ & ~new_n47516_;
  assign new_n47518_ = ~new_n47348_ & new_n47517_;
  assign new_n47519_ = ~new_n47512_ & ~new_n47518_;
  assign new_n47520_ = ~\b[33]  & ~new_n47519_;
  assign new_n47521_ = ~new_n46826_ & ~new_n47349_;
  assign new_n47522_ = ~new_n46836_ & new_n47246_;
  assign new_n47523_ = ~new_n47242_ & new_n47522_;
  assign new_n47524_ = ~new_n47243_ & ~new_n47246_;
  assign new_n47525_ = ~new_n47523_ & ~new_n47524_;
  assign new_n47526_ = new_n288_ & ~new_n47525_;
  assign new_n47527_ = ~new_n47348_ & new_n47526_;
  assign new_n47528_ = ~new_n47521_ & ~new_n47527_;
  assign new_n47529_ = ~\b[32]  & ~new_n47528_;
  assign new_n47530_ = ~new_n46835_ & ~new_n47349_;
  assign new_n47531_ = ~new_n46845_ & new_n47241_;
  assign new_n47532_ = ~new_n47237_ & new_n47531_;
  assign new_n47533_ = ~new_n47238_ & ~new_n47241_;
  assign new_n47534_ = ~new_n47532_ & ~new_n47533_;
  assign new_n47535_ = new_n288_ & ~new_n47534_;
  assign new_n47536_ = ~new_n47348_ & new_n47535_;
  assign new_n47537_ = ~new_n47530_ & ~new_n47536_;
  assign new_n47538_ = ~\b[31]  & ~new_n47537_;
  assign new_n47539_ = ~new_n46844_ & ~new_n47349_;
  assign new_n47540_ = ~new_n46854_ & new_n47236_;
  assign new_n47541_ = ~new_n47232_ & new_n47540_;
  assign new_n47542_ = ~new_n47233_ & ~new_n47236_;
  assign new_n47543_ = ~new_n47541_ & ~new_n47542_;
  assign new_n47544_ = new_n288_ & ~new_n47543_;
  assign new_n47545_ = ~new_n47348_ & new_n47544_;
  assign new_n47546_ = ~new_n47539_ & ~new_n47545_;
  assign new_n47547_ = ~\b[30]  & ~new_n47546_;
  assign new_n47548_ = ~new_n46853_ & ~new_n47349_;
  assign new_n47549_ = ~new_n46863_ & new_n47231_;
  assign new_n47550_ = ~new_n47227_ & new_n47549_;
  assign new_n47551_ = ~new_n47228_ & ~new_n47231_;
  assign new_n47552_ = ~new_n47550_ & ~new_n47551_;
  assign new_n47553_ = new_n288_ & ~new_n47552_;
  assign new_n47554_ = ~new_n47348_ & new_n47553_;
  assign new_n47555_ = ~new_n47548_ & ~new_n47554_;
  assign new_n47556_ = ~\b[29]  & ~new_n47555_;
  assign new_n47557_ = ~new_n46862_ & ~new_n47349_;
  assign new_n47558_ = ~new_n46872_ & new_n47226_;
  assign new_n47559_ = ~new_n47222_ & new_n47558_;
  assign new_n47560_ = ~new_n47223_ & ~new_n47226_;
  assign new_n47561_ = ~new_n47559_ & ~new_n47560_;
  assign new_n47562_ = new_n288_ & ~new_n47561_;
  assign new_n47563_ = ~new_n47348_ & new_n47562_;
  assign new_n47564_ = ~new_n47557_ & ~new_n47563_;
  assign new_n47565_ = ~\b[28]  & ~new_n47564_;
  assign new_n47566_ = ~new_n46871_ & ~new_n47349_;
  assign new_n47567_ = ~new_n46881_ & new_n47221_;
  assign new_n47568_ = ~new_n47217_ & new_n47567_;
  assign new_n47569_ = ~new_n47218_ & ~new_n47221_;
  assign new_n47570_ = ~new_n47568_ & ~new_n47569_;
  assign new_n47571_ = new_n288_ & ~new_n47570_;
  assign new_n47572_ = ~new_n47348_ & new_n47571_;
  assign new_n47573_ = ~new_n47566_ & ~new_n47572_;
  assign new_n47574_ = ~\b[27]  & ~new_n47573_;
  assign new_n47575_ = ~new_n46880_ & ~new_n47349_;
  assign new_n47576_ = ~new_n46890_ & new_n47216_;
  assign new_n47577_ = ~new_n47212_ & new_n47576_;
  assign new_n47578_ = ~new_n47213_ & ~new_n47216_;
  assign new_n47579_ = ~new_n47577_ & ~new_n47578_;
  assign new_n47580_ = new_n288_ & ~new_n47579_;
  assign new_n47581_ = ~new_n47348_ & new_n47580_;
  assign new_n47582_ = ~new_n47575_ & ~new_n47581_;
  assign new_n47583_ = ~\b[26]  & ~new_n47582_;
  assign new_n47584_ = ~new_n46889_ & ~new_n47349_;
  assign new_n47585_ = ~new_n46899_ & new_n47211_;
  assign new_n47586_ = ~new_n47207_ & new_n47585_;
  assign new_n47587_ = ~new_n47208_ & ~new_n47211_;
  assign new_n47588_ = ~new_n47586_ & ~new_n47587_;
  assign new_n47589_ = new_n288_ & ~new_n47588_;
  assign new_n47590_ = ~new_n47348_ & new_n47589_;
  assign new_n47591_ = ~new_n47584_ & ~new_n47590_;
  assign new_n47592_ = ~\b[25]  & ~new_n47591_;
  assign new_n47593_ = ~new_n46898_ & ~new_n47349_;
  assign new_n47594_ = ~new_n46908_ & new_n47206_;
  assign new_n47595_ = ~new_n47202_ & new_n47594_;
  assign new_n47596_ = ~new_n47203_ & ~new_n47206_;
  assign new_n47597_ = ~new_n47595_ & ~new_n47596_;
  assign new_n47598_ = new_n288_ & ~new_n47597_;
  assign new_n47599_ = ~new_n47348_ & new_n47598_;
  assign new_n47600_ = ~new_n47593_ & ~new_n47599_;
  assign new_n47601_ = ~\b[24]  & ~new_n47600_;
  assign new_n47602_ = ~new_n46907_ & ~new_n47349_;
  assign new_n47603_ = ~new_n46917_ & new_n47201_;
  assign new_n47604_ = ~new_n47197_ & new_n47603_;
  assign new_n47605_ = ~new_n47198_ & ~new_n47201_;
  assign new_n47606_ = ~new_n47604_ & ~new_n47605_;
  assign new_n47607_ = new_n288_ & ~new_n47606_;
  assign new_n47608_ = ~new_n47348_ & new_n47607_;
  assign new_n47609_ = ~new_n47602_ & ~new_n47608_;
  assign new_n47610_ = ~\b[23]  & ~new_n47609_;
  assign new_n47611_ = ~new_n46916_ & ~new_n47349_;
  assign new_n47612_ = ~new_n46926_ & new_n47196_;
  assign new_n47613_ = ~new_n47192_ & new_n47612_;
  assign new_n47614_ = ~new_n47193_ & ~new_n47196_;
  assign new_n47615_ = ~new_n47613_ & ~new_n47614_;
  assign new_n47616_ = new_n288_ & ~new_n47615_;
  assign new_n47617_ = ~new_n47348_ & new_n47616_;
  assign new_n47618_ = ~new_n47611_ & ~new_n47617_;
  assign new_n47619_ = ~\b[22]  & ~new_n47618_;
  assign new_n47620_ = ~new_n46925_ & ~new_n47349_;
  assign new_n47621_ = ~new_n46935_ & new_n47191_;
  assign new_n47622_ = ~new_n47187_ & new_n47621_;
  assign new_n47623_ = ~new_n47188_ & ~new_n47191_;
  assign new_n47624_ = ~new_n47622_ & ~new_n47623_;
  assign new_n47625_ = new_n288_ & ~new_n47624_;
  assign new_n47626_ = ~new_n47348_ & new_n47625_;
  assign new_n47627_ = ~new_n47620_ & ~new_n47626_;
  assign new_n47628_ = ~\b[21]  & ~new_n47627_;
  assign new_n47629_ = ~new_n46934_ & ~new_n47349_;
  assign new_n47630_ = ~new_n46944_ & new_n47186_;
  assign new_n47631_ = ~new_n47182_ & new_n47630_;
  assign new_n47632_ = ~new_n47183_ & ~new_n47186_;
  assign new_n47633_ = ~new_n47631_ & ~new_n47632_;
  assign new_n47634_ = new_n288_ & ~new_n47633_;
  assign new_n47635_ = ~new_n47348_ & new_n47634_;
  assign new_n47636_ = ~new_n47629_ & ~new_n47635_;
  assign new_n47637_ = ~\b[20]  & ~new_n47636_;
  assign new_n47638_ = ~new_n46943_ & ~new_n47349_;
  assign new_n47639_ = ~new_n46953_ & new_n47181_;
  assign new_n47640_ = ~new_n47177_ & new_n47639_;
  assign new_n47641_ = ~new_n47178_ & ~new_n47181_;
  assign new_n47642_ = ~new_n47640_ & ~new_n47641_;
  assign new_n47643_ = new_n288_ & ~new_n47642_;
  assign new_n47644_ = ~new_n47348_ & new_n47643_;
  assign new_n47645_ = ~new_n47638_ & ~new_n47644_;
  assign new_n47646_ = ~\b[19]  & ~new_n47645_;
  assign new_n47647_ = ~new_n46952_ & ~new_n47349_;
  assign new_n47648_ = ~new_n46962_ & new_n47176_;
  assign new_n47649_ = ~new_n47172_ & new_n47648_;
  assign new_n47650_ = ~new_n47173_ & ~new_n47176_;
  assign new_n47651_ = ~new_n47649_ & ~new_n47650_;
  assign new_n47652_ = new_n288_ & ~new_n47651_;
  assign new_n47653_ = ~new_n47348_ & new_n47652_;
  assign new_n47654_ = ~new_n47647_ & ~new_n47653_;
  assign new_n47655_ = ~\b[18]  & ~new_n47654_;
  assign new_n47656_ = ~new_n46961_ & ~new_n47349_;
  assign new_n47657_ = ~new_n46971_ & new_n47171_;
  assign new_n47658_ = ~new_n47167_ & new_n47657_;
  assign new_n47659_ = ~new_n47168_ & ~new_n47171_;
  assign new_n47660_ = ~new_n47658_ & ~new_n47659_;
  assign new_n47661_ = new_n288_ & ~new_n47660_;
  assign new_n47662_ = ~new_n47348_ & new_n47661_;
  assign new_n47663_ = ~new_n47656_ & ~new_n47662_;
  assign new_n47664_ = ~\b[17]  & ~new_n47663_;
  assign new_n47665_ = ~new_n46970_ & ~new_n47349_;
  assign new_n47666_ = ~new_n46980_ & new_n47166_;
  assign new_n47667_ = ~new_n47162_ & new_n47666_;
  assign new_n47668_ = ~new_n47163_ & ~new_n47166_;
  assign new_n47669_ = ~new_n47667_ & ~new_n47668_;
  assign new_n47670_ = new_n288_ & ~new_n47669_;
  assign new_n47671_ = ~new_n47348_ & new_n47670_;
  assign new_n47672_ = ~new_n47665_ & ~new_n47671_;
  assign new_n47673_ = ~\b[16]  & ~new_n47672_;
  assign new_n47674_ = ~new_n46979_ & ~new_n47349_;
  assign new_n47675_ = ~new_n46989_ & new_n47161_;
  assign new_n47676_ = ~new_n47157_ & new_n47675_;
  assign new_n47677_ = ~new_n47158_ & ~new_n47161_;
  assign new_n47678_ = ~new_n47676_ & ~new_n47677_;
  assign new_n47679_ = new_n288_ & ~new_n47678_;
  assign new_n47680_ = ~new_n47348_ & new_n47679_;
  assign new_n47681_ = ~new_n47674_ & ~new_n47680_;
  assign new_n47682_ = ~\b[15]  & ~new_n47681_;
  assign new_n47683_ = ~new_n46988_ & ~new_n47349_;
  assign new_n47684_ = ~new_n46998_ & new_n47156_;
  assign new_n47685_ = ~new_n47152_ & new_n47684_;
  assign new_n47686_ = ~new_n47153_ & ~new_n47156_;
  assign new_n47687_ = ~new_n47685_ & ~new_n47686_;
  assign new_n47688_ = new_n288_ & ~new_n47687_;
  assign new_n47689_ = ~new_n47348_ & new_n47688_;
  assign new_n47690_ = ~new_n47683_ & ~new_n47689_;
  assign new_n47691_ = ~\b[14]  & ~new_n47690_;
  assign new_n47692_ = ~new_n46997_ & ~new_n47349_;
  assign new_n47693_ = ~new_n47007_ & new_n47151_;
  assign new_n47694_ = ~new_n47147_ & new_n47693_;
  assign new_n47695_ = ~new_n47148_ & ~new_n47151_;
  assign new_n47696_ = ~new_n47694_ & ~new_n47695_;
  assign new_n47697_ = new_n288_ & ~new_n47696_;
  assign new_n47698_ = ~new_n47348_ & new_n47697_;
  assign new_n47699_ = ~new_n47692_ & ~new_n47698_;
  assign new_n47700_ = ~\b[13]  & ~new_n47699_;
  assign new_n47701_ = ~new_n47006_ & ~new_n47349_;
  assign new_n47702_ = ~new_n47016_ & new_n47146_;
  assign new_n47703_ = ~new_n47142_ & new_n47702_;
  assign new_n47704_ = ~new_n47143_ & ~new_n47146_;
  assign new_n47705_ = ~new_n47703_ & ~new_n47704_;
  assign new_n47706_ = new_n288_ & ~new_n47705_;
  assign new_n47707_ = ~new_n47348_ & new_n47706_;
  assign new_n47708_ = ~new_n47701_ & ~new_n47707_;
  assign new_n47709_ = ~\b[12]  & ~new_n47708_;
  assign new_n47710_ = ~new_n47015_ & ~new_n47349_;
  assign new_n47711_ = ~new_n47025_ & new_n47141_;
  assign new_n47712_ = ~new_n47137_ & new_n47711_;
  assign new_n47713_ = ~new_n47138_ & ~new_n47141_;
  assign new_n47714_ = ~new_n47712_ & ~new_n47713_;
  assign new_n47715_ = new_n288_ & ~new_n47714_;
  assign new_n47716_ = ~new_n47348_ & new_n47715_;
  assign new_n47717_ = ~new_n47710_ & ~new_n47716_;
  assign new_n47718_ = ~\b[11]  & ~new_n47717_;
  assign new_n47719_ = ~new_n47024_ & ~new_n47349_;
  assign new_n47720_ = ~new_n47034_ & new_n47136_;
  assign new_n47721_ = ~new_n47132_ & new_n47720_;
  assign new_n47722_ = ~new_n47133_ & ~new_n47136_;
  assign new_n47723_ = ~new_n47721_ & ~new_n47722_;
  assign new_n47724_ = new_n288_ & ~new_n47723_;
  assign new_n47725_ = ~new_n47348_ & new_n47724_;
  assign new_n47726_ = ~new_n47719_ & ~new_n47725_;
  assign new_n47727_ = ~\b[10]  & ~new_n47726_;
  assign new_n47728_ = ~new_n47033_ & ~new_n47349_;
  assign new_n47729_ = ~new_n47043_ & new_n47131_;
  assign new_n47730_ = ~new_n47127_ & new_n47729_;
  assign new_n47731_ = ~new_n47128_ & ~new_n47131_;
  assign new_n47732_ = ~new_n47730_ & ~new_n47731_;
  assign new_n47733_ = new_n288_ & ~new_n47732_;
  assign new_n47734_ = ~new_n47348_ & new_n47733_;
  assign new_n47735_ = ~new_n47728_ & ~new_n47734_;
  assign new_n47736_ = ~\b[9]  & ~new_n47735_;
  assign new_n47737_ = ~new_n47042_ & ~new_n47349_;
  assign new_n47738_ = ~new_n47052_ & new_n47126_;
  assign new_n47739_ = ~new_n47122_ & new_n47738_;
  assign new_n47740_ = ~new_n47123_ & ~new_n47126_;
  assign new_n47741_ = ~new_n47739_ & ~new_n47740_;
  assign new_n47742_ = new_n288_ & ~new_n47741_;
  assign new_n47743_ = ~new_n47348_ & new_n47742_;
  assign new_n47744_ = ~new_n47737_ & ~new_n47743_;
  assign new_n47745_ = ~\b[8]  & ~new_n47744_;
  assign new_n47746_ = ~new_n47051_ & ~new_n47349_;
  assign new_n47747_ = ~new_n47061_ & new_n47121_;
  assign new_n47748_ = ~new_n47117_ & new_n47747_;
  assign new_n47749_ = ~new_n47118_ & ~new_n47121_;
  assign new_n47750_ = ~new_n47748_ & ~new_n47749_;
  assign new_n47751_ = new_n288_ & ~new_n47750_;
  assign new_n47752_ = ~new_n47348_ & new_n47751_;
  assign new_n47753_ = ~new_n47746_ & ~new_n47752_;
  assign new_n47754_ = ~\b[7]  & ~new_n47753_;
  assign new_n47755_ = ~new_n47060_ & ~new_n47349_;
  assign new_n47756_ = ~new_n47070_ & new_n47116_;
  assign new_n47757_ = ~new_n47112_ & new_n47756_;
  assign new_n47758_ = ~new_n47113_ & ~new_n47116_;
  assign new_n47759_ = ~new_n47757_ & ~new_n47758_;
  assign new_n47760_ = new_n288_ & ~new_n47759_;
  assign new_n47761_ = ~new_n47348_ & new_n47760_;
  assign new_n47762_ = ~new_n47755_ & ~new_n47761_;
  assign new_n47763_ = ~\b[6]  & ~new_n47762_;
  assign new_n47764_ = ~new_n47069_ & ~new_n47349_;
  assign new_n47765_ = ~new_n47079_ & new_n47111_;
  assign new_n47766_ = ~new_n47107_ & new_n47765_;
  assign new_n47767_ = ~new_n47108_ & ~new_n47111_;
  assign new_n47768_ = ~new_n47766_ & ~new_n47767_;
  assign new_n47769_ = new_n288_ & ~new_n47768_;
  assign new_n47770_ = ~new_n47348_ & new_n47769_;
  assign new_n47771_ = ~new_n47764_ & ~new_n47770_;
  assign new_n47772_ = ~\b[5]  & ~new_n47771_;
  assign new_n47773_ = ~new_n47078_ & ~new_n47349_;
  assign new_n47774_ = ~new_n47087_ & new_n47106_;
  assign new_n47775_ = ~new_n47102_ & new_n47774_;
  assign new_n47776_ = ~new_n47103_ & ~new_n47106_;
  assign new_n47777_ = ~new_n47775_ & ~new_n47776_;
  assign new_n47778_ = new_n288_ & ~new_n47777_;
  assign new_n47779_ = ~new_n47348_ & new_n47778_;
  assign new_n47780_ = ~new_n47773_ & ~new_n47779_;
  assign new_n47781_ = ~\b[4]  & ~new_n47780_;
  assign new_n47782_ = ~new_n47086_ & ~new_n47349_;
  assign new_n47783_ = ~new_n47097_ & new_n47101_;
  assign new_n47784_ = ~new_n47096_ & new_n47783_;
  assign new_n47785_ = ~new_n47098_ & ~new_n47101_;
  assign new_n47786_ = ~new_n47784_ & ~new_n47785_;
  assign new_n47787_ = new_n288_ & ~new_n47786_;
  assign new_n47788_ = ~new_n47348_ & new_n47787_;
  assign new_n47789_ = ~new_n47782_ & ~new_n47788_;
  assign new_n47790_ = ~\b[3]  & ~new_n47789_;
  assign new_n47791_ = ~new_n47091_ & ~new_n47349_;
  assign new_n47792_ = new_n19050_ & ~new_n47094_;
  assign new_n47793_ = ~new_n47092_ & new_n47792_;
  assign new_n47794_ = new_n288_ & ~new_n47793_;
  assign new_n47795_ = ~new_n47096_ & new_n47794_;
  assign new_n47796_ = ~new_n47348_ & new_n47795_;
  assign new_n47797_ = ~new_n47791_ & ~new_n47796_;
  assign new_n47798_ = ~\b[2]  & ~new_n47797_;
  assign new_n47799_ = new_n19756_ & ~new_n47348_;
  assign new_n47800_ = \a[12]  & ~new_n47799_;
  assign new_n47801_ = new_n19760_ & ~new_n47348_;
  assign new_n47802_ = ~new_n47800_ & ~new_n47801_;
  assign new_n47803_ = \b[1]  & ~new_n47802_;
  assign new_n47804_ = ~\b[1]  & ~new_n47801_;
  assign new_n47805_ = ~new_n47800_ & new_n47804_;
  assign new_n47806_ = ~new_n47803_ & ~new_n47805_;
  assign new_n47807_ = ~new_n19767_ & ~new_n47806_;
  assign new_n47808_ = ~\b[1]  & ~new_n47802_;
  assign new_n47809_ = ~new_n47807_ & ~new_n47808_;
  assign new_n47810_ = \b[2]  & ~new_n47796_;
  assign new_n47811_ = ~new_n47791_ & new_n47810_;
  assign new_n47812_ = ~new_n47798_ & ~new_n47811_;
  assign new_n47813_ = ~new_n47809_ & new_n47812_;
  assign new_n47814_ = ~new_n47798_ & ~new_n47813_;
  assign new_n47815_ = \b[3]  & ~new_n47788_;
  assign new_n47816_ = ~new_n47782_ & new_n47815_;
  assign new_n47817_ = ~new_n47790_ & ~new_n47816_;
  assign new_n47818_ = ~new_n47814_ & new_n47817_;
  assign new_n47819_ = ~new_n47790_ & ~new_n47818_;
  assign new_n47820_ = \b[4]  & ~new_n47779_;
  assign new_n47821_ = ~new_n47773_ & new_n47820_;
  assign new_n47822_ = ~new_n47781_ & ~new_n47821_;
  assign new_n47823_ = ~new_n47819_ & new_n47822_;
  assign new_n47824_ = ~new_n47781_ & ~new_n47823_;
  assign new_n47825_ = \b[5]  & ~new_n47770_;
  assign new_n47826_ = ~new_n47764_ & new_n47825_;
  assign new_n47827_ = ~new_n47772_ & ~new_n47826_;
  assign new_n47828_ = ~new_n47824_ & new_n47827_;
  assign new_n47829_ = ~new_n47772_ & ~new_n47828_;
  assign new_n47830_ = \b[6]  & ~new_n47761_;
  assign new_n47831_ = ~new_n47755_ & new_n47830_;
  assign new_n47832_ = ~new_n47763_ & ~new_n47831_;
  assign new_n47833_ = ~new_n47829_ & new_n47832_;
  assign new_n47834_ = ~new_n47763_ & ~new_n47833_;
  assign new_n47835_ = \b[7]  & ~new_n47752_;
  assign new_n47836_ = ~new_n47746_ & new_n47835_;
  assign new_n47837_ = ~new_n47754_ & ~new_n47836_;
  assign new_n47838_ = ~new_n47834_ & new_n47837_;
  assign new_n47839_ = ~new_n47754_ & ~new_n47838_;
  assign new_n47840_ = \b[8]  & ~new_n47743_;
  assign new_n47841_ = ~new_n47737_ & new_n47840_;
  assign new_n47842_ = ~new_n47745_ & ~new_n47841_;
  assign new_n47843_ = ~new_n47839_ & new_n47842_;
  assign new_n47844_ = ~new_n47745_ & ~new_n47843_;
  assign new_n47845_ = \b[9]  & ~new_n47734_;
  assign new_n47846_ = ~new_n47728_ & new_n47845_;
  assign new_n47847_ = ~new_n47736_ & ~new_n47846_;
  assign new_n47848_ = ~new_n47844_ & new_n47847_;
  assign new_n47849_ = ~new_n47736_ & ~new_n47848_;
  assign new_n47850_ = \b[10]  & ~new_n47725_;
  assign new_n47851_ = ~new_n47719_ & new_n47850_;
  assign new_n47852_ = ~new_n47727_ & ~new_n47851_;
  assign new_n47853_ = ~new_n47849_ & new_n47852_;
  assign new_n47854_ = ~new_n47727_ & ~new_n47853_;
  assign new_n47855_ = \b[11]  & ~new_n47716_;
  assign new_n47856_ = ~new_n47710_ & new_n47855_;
  assign new_n47857_ = ~new_n47718_ & ~new_n47856_;
  assign new_n47858_ = ~new_n47854_ & new_n47857_;
  assign new_n47859_ = ~new_n47718_ & ~new_n47858_;
  assign new_n47860_ = \b[12]  & ~new_n47707_;
  assign new_n47861_ = ~new_n47701_ & new_n47860_;
  assign new_n47862_ = ~new_n47709_ & ~new_n47861_;
  assign new_n47863_ = ~new_n47859_ & new_n47862_;
  assign new_n47864_ = ~new_n47709_ & ~new_n47863_;
  assign new_n47865_ = \b[13]  & ~new_n47698_;
  assign new_n47866_ = ~new_n47692_ & new_n47865_;
  assign new_n47867_ = ~new_n47700_ & ~new_n47866_;
  assign new_n47868_ = ~new_n47864_ & new_n47867_;
  assign new_n47869_ = ~new_n47700_ & ~new_n47868_;
  assign new_n47870_ = \b[14]  & ~new_n47689_;
  assign new_n47871_ = ~new_n47683_ & new_n47870_;
  assign new_n47872_ = ~new_n47691_ & ~new_n47871_;
  assign new_n47873_ = ~new_n47869_ & new_n47872_;
  assign new_n47874_ = ~new_n47691_ & ~new_n47873_;
  assign new_n47875_ = \b[15]  & ~new_n47680_;
  assign new_n47876_ = ~new_n47674_ & new_n47875_;
  assign new_n47877_ = ~new_n47682_ & ~new_n47876_;
  assign new_n47878_ = ~new_n47874_ & new_n47877_;
  assign new_n47879_ = ~new_n47682_ & ~new_n47878_;
  assign new_n47880_ = \b[16]  & ~new_n47671_;
  assign new_n47881_ = ~new_n47665_ & new_n47880_;
  assign new_n47882_ = ~new_n47673_ & ~new_n47881_;
  assign new_n47883_ = ~new_n47879_ & new_n47882_;
  assign new_n47884_ = ~new_n47673_ & ~new_n47883_;
  assign new_n47885_ = \b[17]  & ~new_n47662_;
  assign new_n47886_ = ~new_n47656_ & new_n47885_;
  assign new_n47887_ = ~new_n47664_ & ~new_n47886_;
  assign new_n47888_ = ~new_n47884_ & new_n47887_;
  assign new_n47889_ = ~new_n47664_ & ~new_n47888_;
  assign new_n47890_ = \b[18]  & ~new_n47653_;
  assign new_n47891_ = ~new_n47647_ & new_n47890_;
  assign new_n47892_ = ~new_n47655_ & ~new_n47891_;
  assign new_n47893_ = ~new_n47889_ & new_n47892_;
  assign new_n47894_ = ~new_n47655_ & ~new_n47893_;
  assign new_n47895_ = \b[19]  & ~new_n47644_;
  assign new_n47896_ = ~new_n47638_ & new_n47895_;
  assign new_n47897_ = ~new_n47646_ & ~new_n47896_;
  assign new_n47898_ = ~new_n47894_ & new_n47897_;
  assign new_n47899_ = ~new_n47646_ & ~new_n47898_;
  assign new_n47900_ = \b[20]  & ~new_n47635_;
  assign new_n47901_ = ~new_n47629_ & new_n47900_;
  assign new_n47902_ = ~new_n47637_ & ~new_n47901_;
  assign new_n47903_ = ~new_n47899_ & new_n47902_;
  assign new_n47904_ = ~new_n47637_ & ~new_n47903_;
  assign new_n47905_ = \b[21]  & ~new_n47626_;
  assign new_n47906_ = ~new_n47620_ & new_n47905_;
  assign new_n47907_ = ~new_n47628_ & ~new_n47906_;
  assign new_n47908_ = ~new_n47904_ & new_n47907_;
  assign new_n47909_ = ~new_n47628_ & ~new_n47908_;
  assign new_n47910_ = \b[22]  & ~new_n47617_;
  assign new_n47911_ = ~new_n47611_ & new_n47910_;
  assign new_n47912_ = ~new_n47619_ & ~new_n47911_;
  assign new_n47913_ = ~new_n47909_ & new_n47912_;
  assign new_n47914_ = ~new_n47619_ & ~new_n47913_;
  assign new_n47915_ = \b[23]  & ~new_n47608_;
  assign new_n47916_ = ~new_n47602_ & new_n47915_;
  assign new_n47917_ = ~new_n47610_ & ~new_n47916_;
  assign new_n47918_ = ~new_n47914_ & new_n47917_;
  assign new_n47919_ = ~new_n47610_ & ~new_n47918_;
  assign new_n47920_ = \b[24]  & ~new_n47599_;
  assign new_n47921_ = ~new_n47593_ & new_n47920_;
  assign new_n47922_ = ~new_n47601_ & ~new_n47921_;
  assign new_n47923_ = ~new_n47919_ & new_n47922_;
  assign new_n47924_ = ~new_n47601_ & ~new_n47923_;
  assign new_n47925_ = \b[25]  & ~new_n47590_;
  assign new_n47926_ = ~new_n47584_ & new_n47925_;
  assign new_n47927_ = ~new_n47592_ & ~new_n47926_;
  assign new_n47928_ = ~new_n47924_ & new_n47927_;
  assign new_n47929_ = ~new_n47592_ & ~new_n47928_;
  assign new_n47930_ = \b[26]  & ~new_n47581_;
  assign new_n47931_ = ~new_n47575_ & new_n47930_;
  assign new_n47932_ = ~new_n47583_ & ~new_n47931_;
  assign new_n47933_ = ~new_n47929_ & new_n47932_;
  assign new_n47934_ = ~new_n47583_ & ~new_n47933_;
  assign new_n47935_ = \b[27]  & ~new_n47572_;
  assign new_n47936_ = ~new_n47566_ & new_n47935_;
  assign new_n47937_ = ~new_n47574_ & ~new_n47936_;
  assign new_n47938_ = ~new_n47934_ & new_n47937_;
  assign new_n47939_ = ~new_n47574_ & ~new_n47938_;
  assign new_n47940_ = \b[28]  & ~new_n47563_;
  assign new_n47941_ = ~new_n47557_ & new_n47940_;
  assign new_n47942_ = ~new_n47565_ & ~new_n47941_;
  assign new_n47943_ = ~new_n47939_ & new_n47942_;
  assign new_n47944_ = ~new_n47565_ & ~new_n47943_;
  assign new_n47945_ = \b[29]  & ~new_n47554_;
  assign new_n47946_ = ~new_n47548_ & new_n47945_;
  assign new_n47947_ = ~new_n47556_ & ~new_n47946_;
  assign new_n47948_ = ~new_n47944_ & new_n47947_;
  assign new_n47949_ = ~new_n47556_ & ~new_n47948_;
  assign new_n47950_ = \b[30]  & ~new_n47545_;
  assign new_n47951_ = ~new_n47539_ & new_n47950_;
  assign new_n47952_ = ~new_n47547_ & ~new_n47951_;
  assign new_n47953_ = ~new_n47949_ & new_n47952_;
  assign new_n47954_ = ~new_n47547_ & ~new_n47953_;
  assign new_n47955_ = \b[31]  & ~new_n47536_;
  assign new_n47956_ = ~new_n47530_ & new_n47955_;
  assign new_n47957_ = ~new_n47538_ & ~new_n47956_;
  assign new_n47958_ = ~new_n47954_ & new_n47957_;
  assign new_n47959_ = ~new_n47538_ & ~new_n47958_;
  assign new_n47960_ = \b[32]  & ~new_n47527_;
  assign new_n47961_ = ~new_n47521_ & new_n47960_;
  assign new_n47962_ = ~new_n47529_ & ~new_n47961_;
  assign new_n47963_ = ~new_n47959_ & new_n47962_;
  assign new_n47964_ = ~new_n47529_ & ~new_n47963_;
  assign new_n47965_ = \b[33]  & ~new_n47518_;
  assign new_n47966_ = ~new_n47512_ & new_n47965_;
  assign new_n47967_ = ~new_n47520_ & ~new_n47966_;
  assign new_n47968_ = ~new_n47964_ & new_n47967_;
  assign new_n47969_ = ~new_n47520_ & ~new_n47968_;
  assign new_n47970_ = \b[34]  & ~new_n47509_;
  assign new_n47971_ = ~new_n47503_ & new_n47970_;
  assign new_n47972_ = ~new_n47511_ & ~new_n47971_;
  assign new_n47973_ = ~new_n47969_ & new_n47972_;
  assign new_n47974_ = ~new_n47511_ & ~new_n47973_;
  assign new_n47975_ = \b[35]  & ~new_n47500_;
  assign new_n47976_ = ~new_n47494_ & new_n47975_;
  assign new_n47977_ = ~new_n47502_ & ~new_n47976_;
  assign new_n47978_ = ~new_n47974_ & new_n47977_;
  assign new_n47979_ = ~new_n47502_ & ~new_n47978_;
  assign new_n47980_ = \b[36]  & ~new_n47491_;
  assign new_n47981_ = ~new_n47485_ & new_n47980_;
  assign new_n47982_ = ~new_n47493_ & ~new_n47981_;
  assign new_n47983_ = ~new_n47979_ & new_n47982_;
  assign new_n47984_ = ~new_n47493_ & ~new_n47983_;
  assign new_n47985_ = \b[37]  & ~new_n47482_;
  assign new_n47986_ = ~new_n47476_ & new_n47985_;
  assign new_n47987_ = ~new_n47484_ & ~new_n47986_;
  assign new_n47988_ = ~new_n47984_ & new_n47987_;
  assign new_n47989_ = ~new_n47484_ & ~new_n47988_;
  assign new_n47990_ = \b[38]  & ~new_n47473_;
  assign new_n47991_ = ~new_n47467_ & new_n47990_;
  assign new_n47992_ = ~new_n47475_ & ~new_n47991_;
  assign new_n47993_ = ~new_n47989_ & new_n47992_;
  assign new_n47994_ = ~new_n47475_ & ~new_n47993_;
  assign new_n47995_ = \b[39]  & ~new_n47464_;
  assign new_n47996_ = ~new_n47458_ & new_n47995_;
  assign new_n47997_ = ~new_n47466_ & ~new_n47996_;
  assign new_n47998_ = ~new_n47994_ & new_n47997_;
  assign new_n47999_ = ~new_n47466_ & ~new_n47998_;
  assign new_n48000_ = \b[40]  & ~new_n47455_;
  assign new_n48001_ = ~new_n47449_ & new_n48000_;
  assign new_n48002_ = ~new_n47457_ & ~new_n48001_;
  assign new_n48003_ = ~new_n47999_ & new_n48002_;
  assign new_n48004_ = ~new_n47457_ & ~new_n48003_;
  assign new_n48005_ = \b[41]  & ~new_n47446_;
  assign new_n48006_ = ~new_n47440_ & new_n48005_;
  assign new_n48007_ = ~new_n47448_ & ~new_n48006_;
  assign new_n48008_ = ~new_n48004_ & new_n48007_;
  assign new_n48009_ = ~new_n47448_ & ~new_n48008_;
  assign new_n48010_ = \b[42]  & ~new_n47437_;
  assign new_n48011_ = ~new_n47431_ & new_n48010_;
  assign new_n48012_ = ~new_n47439_ & ~new_n48011_;
  assign new_n48013_ = ~new_n48009_ & new_n48012_;
  assign new_n48014_ = ~new_n47439_ & ~new_n48013_;
  assign new_n48015_ = \b[43]  & ~new_n47428_;
  assign new_n48016_ = ~new_n47422_ & new_n48015_;
  assign new_n48017_ = ~new_n47430_ & ~new_n48016_;
  assign new_n48018_ = ~new_n48014_ & new_n48017_;
  assign new_n48019_ = ~new_n47430_ & ~new_n48018_;
  assign new_n48020_ = \b[44]  & ~new_n47419_;
  assign new_n48021_ = ~new_n47413_ & new_n48020_;
  assign new_n48022_ = ~new_n47421_ & ~new_n48021_;
  assign new_n48023_ = ~new_n48019_ & new_n48022_;
  assign new_n48024_ = ~new_n47421_ & ~new_n48023_;
  assign new_n48025_ = \b[45]  & ~new_n47410_;
  assign new_n48026_ = ~new_n47404_ & new_n48025_;
  assign new_n48027_ = ~new_n47412_ & ~new_n48026_;
  assign new_n48028_ = ~new_n48024_ & new_n48027_;
  assign new_n48029_ = ~new_n47412_ & ~new_n48028_;
  assign new_n48030_ = \b[46]  & ~new_n47401_;
  assign new_n48031_ = ~new_n47395_ & new_n48030_;
  assign new_n48032_ = ~new_n47403_ & ~new_n48031_;
  assign new_n48033_ = ~new_n48029_ & new_n48032_;
  assign new_n48034_ = ~new_n47403_ & ~new_n48033_;
  assign new_n48035_ = \b[47]  & ~new_n47392_;
  assign new_n48036_ = ~new_n47386_ & new_n48035_;
  assign new_n48037_ = ~new_n47394_ & ~new_n48036_;
  assign new_n48038_ = ~new_n48034_ & new_n48037_;
  assign new_n48039_ = ~new_n47394_ & ~new_n48038_;
  assign new_n48040_ = \b[48]  & ~new_n47383_;
  assign new_n48041_ = ~new_n47377_ & new_n48040_;
  assign new_n48042_ = ~new_n47385_ & ~new_n48041_;
  assign new_n48043_ = ~new_n48039_ & new_n48042_;
  assign new_n48044_ = ~new_n47385_ & ~new_n48043_;
  assign new_n48045_ = \b[49]  & ~new_n47374_;
  assign new_n48046_ = ~new_n47368_ & new_n48045_;
  assign new_n48047_ = ~new_n47376_ & ~new_n48046_;
  assign new_n48048_ = ~new_n48044_ & new_n48047_;
  assign new_n48049_ = ~new_n47376_ & ~new_n48048_;
  assign new_n48050_ = \b[50]  & ~new_n47365_;
  assign new_n48051_ = ~new_n47359_ & new_n48050_;
  assign new_n48052_ = ~new_n47367_ & ~new_n48051_;
  assign new_n48053_ = ~new_n48049_ & new_n48052_;
  assign new_n48054_ = ~new_n47367_ & ~new_n48053_;
  assign new_n48055_ = \b[51]  & ~new_n47356_;
  assign new_n48056_ = ~new_n47350_ & new_n48055_;
  assign new_n48057_ = ~new_n47358_ & ~new_n48056_;
  assign new_n48058_ = ~new_n48054_ & new_n48057_;
  assign new_n48059_ = ~new_n47358_ & ~new_n48058_;
  assign new_n48060_ = ~new_n46654_ & ~new_n47349_;
  assign new_n48061_ = ~new_n46656_ & new_n47346_;
  assign new_n48062_ = ~new_n47342_ & new_n48061_;
  assign new_n48063_ = ~new_n47343_ & ~new_n47346_;
  assign new_n48064_ = ~new_n48062_ & ~new_n48063_;
  assign new_n48065_ = new_n47349_ & ~new_n48064_;
  assign new_n48066_ = ~new_n48060_ & ~new_n48065_;
  assign new_n48067_ = ~\b[52]  & ~new_n48066_;
  assign new_n48068_ = \b[52]  & ~new_n48060_;
  assign new_n48069_ = ~new_n48065_ & new_n48068_;
  assign new_n48070_ = new_n595_ & ~new_n48069_;
  assign new_n48071_ = ~new_n48067_ & new_n48070_;
  assign new_n48072_ = ~new_n48059_ & new_n48071_;
  assign new_n48073_ = new_n288_ & ~new_n48066_;
  assign new_n48074_ = ~new_n48072_ & ~new_n48073_;
  assign new_n48075_ = ~new_n47367_ & new_n48057_;
  assign new_n48076_ = ~new_n48053_ & new_n48075_;
  assign new_n48077_ = ~new_n48054_ & ~new_n48057_;
  assign new_n48078_ = ~new_n48076_ & ~new_n48077_;
  assign new_n48079_ = ~new_n48074_ & ~new_n48078_;
  assign new_n48080_ = ~new_n47357_ & ~new_n48073_;
  assign new_n48081_ = ~new_n48072_ & new_n48080_;
  assign new_n48082_ = ~new_n48079_ & ~new_n48081_;
  assign new_n48083_ = ~\b[52]  & ~new_n48082_;
  assign new_n48084_ = ~new_n47376_ & new_n48052_;
  assign new_n48085_ = ~new_n48048_ & new_n48084_;
  assign new_n48086_ = ~new_n48049_ & ~new_n48052_;
  assign new_n48087_ = ~new_n48085_ & ~new_n48086_;
  assign new_n48088_ = ~new_n48074_ & ~new_n48087_;
  assign new_n48089_ = ~new_n47366_ & ~new_n48073_;
  assign new_n48090_ = ~new_n48072_ & new_n48089_;
  assign new_n48091_ = ~new_n48088_ & ~new_n48090_;
  assign new_n48092_ = ~\b[51]  & ~new_n48091_;
  assign new_n48093_ = ~new_n47385_ & new_n48047_;
  assign new_n48094_ = ~new_n48043_ & new_n48093_;
  assign new_n48095_ = ~new_n48044_ & ~new_n48047_;
  assign new_n48096_ = ~new_n48094_ & ~new_n48095_;
  assign new_n48097_ = ~new_n48074_ & ~new_n48096_;
  assign new_n48098_ = ~new_n47375_ & ~new_n48073_;
  assign new_n48099_ = ~new_n48072_ & new_n48098_;
  assign new_n48100_ = ~new_n48097_ & ~new_n48099_;
  assign new_n48101_ = ~\b[50]  & ~new_n48100_;
  assign new_n48102_ = ~new_n47394_ & new_n48042_;
  assign new_n48103_ = ~new_n48038_ & new_n48102_;
  assign new_n48104_ = ~new_n48039_ & ~new_n48042_;
  assign new_n48105_ = ~new_n48103_ & ~new_n48104_;
  assign new_n48106_ = ~new_n48074_ & ~new_n48105_;
  assign new_n48107_ = ~new_n47384_ & ~new_n48073_;
  assign new_n48108_ = ~new_n48072_ & new_n48107_;
  assign new_n48109_ = ~new_n48106_ & ~new_n48108_;
  assign new_n48110_ = ~\b[49]  & ~new_n48109_;
  assign new_n48111_ = ~new_n47403_ & new_n48037_;
  assign new_n48112_ = ~new_n48033_ & new_n48111_;
  assign new_n48113_ = ~new_n48034_ & ~new_n48037_;
  assign new_n48114_ = ~new_n48112_ & ~new_n48113_;
  assign new_n48115_ = ~new_n48074_ & ~new_n48114_;
  assign new_n48116_ = ~new_n47393_ & ~new_n48073_;
  assign new_n48117_ = ~new_n48072_ & new_n48116_;
  assign new_n48118_ = ~new_n48115_ & ~new_n48117_;
  assign new_n48119_ = ~\b[48]  & ~new_n48118_;
  assign new_n48120_ = ~new_n47412_ & new_n48032_;
  assign new_n48121_ = ~new_n48028_ & new_n48120_;
  assign new_n48122_ = ~new_n48029_ & ~new_n48032_;
  assign new_n48123_ = ~new_n48121_ & ~new_n48122_;
  assign new_n48124_ = ~new_n48074_ & ~new_n48123_;
  assign new_n48125_ = ~new_n47402_ & ~new_n48073_;
  assign new_n48126_ = ~new_n48072_ & new_n48125_;
  assign new_n48127_ = ~new_n48124_ & ~new_n48126_;
  assign new_n48128_ = ~\b[47]  & ~new_n48127_;
  assign new_n48129_ = ~new_n47421_ & new_n48027_;
  assign new_n48130_ = ~new_n48023_ & new_n48129_;
  assign new_n48131_ = ~new_n48024_ & ~new_n48027_;
  assign new_n48132_ = ~new_n48130_ & ~new_n48131_;
  assign new_n48133_ = ~new_n48074_ & ~new_n48132_;
  assign new_n48134_ = ~new_n47411_ & ~new_n48073_;
  assign new_n48135_ = ~new_n48072_ & new_n48134_;
  assign new_n48136_ = ~new_n48133_ & ~new_n48135_;
  assign new_n48137_ = ~\b[46]  & ~new_n48136_;
  assign new_n48138_ = ~new_n47430_ & new_n48022_;
  assign new_n48139_ = ~new_n48018_ & new_n48138_;
  assign new_n48140_ = ~new_n48019_ & ~new_n48022_;
  assign new_n48141_ = ~new_n48139_ & ~new_n48140_;
  assign new_n48142_ = ~new_n48074_ & ~new_n48141_;
  assign new_n48143_ = ~new_n47420_ & ~new_n48073_;
  assign new_n48144_ = ~new_n48072_ & new_n48143_;
  assign new_n48145_ = ~new_n48142_ & ~new_n48144_;
  assign new_n48146_ = ~\b[45]  & ~new_n48145_;
  assign new_n48147_ = ~new_n47439_ & new_n48017_;
  assign new_n48148_ = ~new_n48013_ & new_n48147_;
  assign new_n48149_ = ~new_n48014_ & ~new_n48017_;
  assign new_n48150_ = ~new_n48148_ & ~new_n48149_;
  assign new_n48151_ = ~new_n48074_ & ~new_n48150_;
  assign new_n48152_ = ~new_n47429_ & ~new_n48073_;
  assign new_n48153_ = ~new_n48072_ & new_n48152_;
  assign new_n48154_ = ~new_n48151_ & ~new_n48153_;
  assign new_n48155_ = ~\b[44]  & ~new_n48154_;
  assign new_n48156_ = ~new_n47448_ & new_n48012_;
  assign new_n48157_ = ~new_n48008_ & new_n48156_;
  assign new_n48158_ = ~new_n48009_ & ~new_n48012_;
  assign new_n48159_ = ~new_n48157_ & ~new_n48158_;
  assign new_n48160_ = ~new_n48074_ & ~new_n48159_;
  assign new_n48161_ = ~new_n47438_ & ~new_n48073_;
  assign new_n48162_ = ~new_n48072_ & new_n48161_;
  assign new_n48163_ = ~new_n48160_ & ~new_n48162_;
  assign new_n48164_ = ~\b[43]  & ~new_n48163_;
  assign new_n48165_ = ~new_n47457_ & new_n48007_;
  assign new_n48166_ = ~new_n48003_ & new_n48165_;
  assign new_n48167_ = ~new_n48004_ & ~new_n48007_;
  assign new_n48168_ = ~new_n48166_ & ~new_n48167_;
  assign new_n48169_ = ~new_n48074_ & ~new_n48168_;
  assign new_n48170_ = ~new_n47447_ & ~new_n48073_;
  assign new_n48171_ = ~new_n48072_ & new_n48170_;
  assign new_n48172_ = ~new_n48169_ & ~new_n48171_;
  assign new_n48173_ = ~\b[42]  & ~new_n48172_;
  assign new_n48174_ = ~new_n47466_ & new_n48002_;
  assign new_n48175_ = ~new_n47998_ & new_n48174_;
  assign new_n48176_ = ~new_n47999_ & ~new_n48002_;
  assign new_n48177_ = ~new_n48175_ & ~new_n48176_;
  assign new_n48178_ = ~new_n48074_ & ~new_n48177_;
  assign new_n48179_ = ~new_n47456_ & ~new_n48073_;
  assign new_n48180_ = ~new_n48072_ & new_n48179_;
  assign new_n48181_ = ~new_n48178_ & ~new_n48180_;
  assign new_n48182_ = ~\b[41]  & ~new_n48181_;
  assign new_n48183_ = ~new_n47475_ & new_n47997_;
  assign new_n48184_ = ~new_n47993_ & new_n48183_;
  assign new_n48185_ = ~new_n47994_ & ~new_n47997_;
  assign new_n48186_ = ~new_n48184_ & ~new_n48185_;
  assign new_n48187_ = ~new_n48074_ & ~new_n48186_;
  assign new_n48188_ = ~new_n47465_ & ~new_n48073_;
  assign new_n48189_ = ~new_n48072_ & new_n48188_;
  assign new_n48190_ = ~new_n48187_ & ~new_n48189_;
  assign new_n48191_ = ~\b[40]  & ~new_n48190_;
  assign new_n48192_ = ~new_n47484_ & new_n47992_;
  assign new_n48193_ = ~new_n47988_ & new_n48192_;
  assign new_n48194_ = ~new_n47989_ & ~new_n47992_;
  assign new_n48195_ = ~new_n48193_ & ~new_n48194_;
  assign new_n48196_ = ~new_n48074_ & ~new_n48195_;
  assign new_n48197_ = ~new_n47474_ & ~new_n48073_;
  assign new_n48198_ = ~new_n48072_ & new_n48197_;
  assign new_n48199_ = ~new_n48196_ & ~new_n48198_;
  assign new_n48200_ = ~\b[39]  & ~new_n48199_;
  assign new_n48201_ = ~new_n47493_ & new_n47987_;
  assign new_n48202_ = ~new_n47983_ & new_n48201_;
  assign new_n48203_ = ~new_n47984_ & ~new_n47987_;
  assign new_n48204_ = ~new_n48202_ & ~new_n48203_;
  assign new_n48205_ = ~new_n48074_ & ~new_n48204_;
  assign new_n48206_ = ~new_n47483_ & ~new_n48073_;
  assign new_n48207_ = ~new_n48072_ & new_n48206_;
  assign new_n48208_ = ~new_n48205_ & ~new_n48207_;
  assign new_n48209_ = ~\b[38]  & ~new_n48208_;
  assign new_n48210_ = ~new_n47502_ & new_n47982_;
  assign new_n48211_ = ~new_n47978_ & new_n48210_;
  assign new_n48212_ = ~new_n47979_ & ~new_n47982_;
  assign new_n48213_ = ~new_n48211_ & ~new_n48212_;
  assign new_n48214_ = ~new_n48074_ & ~new_n48213_;
  assign new_n48215_ = ~new_n47492_ & ~new_n48073_;
  assign new_n48216_ = ~new_n48072_ & new_n48215_;
  assign new_n48217_ = ~new_n48214_ & ~new_n48216_;
  assign new_n48218_ = ~\b[37]  & ~new_n48217_;
  assign new_n48219_ = ~new_n47511_ & new_n47977_;
  assign new_n48220_ = ~new_n47973_ & new_n48219_;
  assign new_n48221_ = ~new_n47974_ & ~new_n47977_;
  assign new_n48222_ = ~new_n48220_ & ~new_n48221_;
  assign new_n48223_ = ~new_n48074_ & ~new_n48222_;
  assign new_n48224_ = ~new_n47501_ & ~new_n48073_;
  assign new_n48225_ = ~new_n48072_ & new_n48224_;
  assign new_n48226_ = ~new_n48223_ & ~new_n48225_;
  assign new_n48227_ = ~\b[36]  & ~new_n48226_;
  assign new_n48228_ = ~new_n47520_ & new_n47972_;
  assign new_n48229_ = ~new_n47968_ & new_n48228_;
  assign new_n48230_ = ~new_n47969_ & ~new_n47972_;
  assign new_n48231_ = ~new_n48229_ & ~new_n48230_;
  assign new_n48232_ = ~new_n48074_ & ~new_n48231_;
  assign new_n48233_ = ~new_n47510_ & ~new_n48073_;
  assign new_n48234_ = ~new_n48072_ & new_n48233_;
  assign new_n48235_ = ~new_n48232_ & ~new_n48234_;
  assign new_n48236_ = ~\b[35]  & ~new_n48235_;
  assign new_n48237_ = ~new_n47529_ & new_n47967_;
  assign new_n48238_ = ~new_n47963_ & new_n48237_;
  assign new_n48239_ = ~new_n47964_ & ~new_n47967_;
  assign new_n48240_ = ~new_n48238_ & ~new_n48239_;
  assign new_n48241_ = ~new_n48074_ & ~new_n48240_;
  assign new_n48242_ = ~new_n47519_ & ~new_n48073_;
  assign new_n48243_ = ~new_n48072_ & new_n48242_;
  assign new_n48244_ = ~new_n48241_ & ~new_n48243_;
  assign new_n48245_ = ~\b[34]  & ~new_n48244_;
  assign new_n48246_ = ~new_n47538_ & new_n47962_;
  assign new_n48247_ = ~new_n47958_ & new_n48246_;
  assign new_n48248_ = ~new_n47959_ & ~new_n47962_;
  assign new_n48249_ = ~new_n48247_ & ~new_n48248_;
  assign new_n48250_ = ~new_n48074_ & ~new_n48249_;
  assign new_n48251_ = ~new_n47528_ & ~new_n48073_;
  assign new_n48252_ = ~new_n48072_ & new_n48251_;
  assign new_n48253_ = ~new_n48250_ & ~new_n48252_;
  assign new_n48254_ = ~\b[33]  & ~new_n48253_;
  assign new_n48255_ = ~new_n47547_ & new_n47957_;
  assign new_n48256_ = ~new_n47953_ & new_n48255_;
  assign new_n48257_ = ~new_n47954_ & ~new_n47957_;
  assign new_n48258_ = ~new_n48256_ & ~new_n48257_;
  assign new_n48259_ = ~new_n48074_ & ~new_n48258_;
  assign new_n48260_ = ~new_n47537_ & ~new_n48073_;
  assign new_n48261_ = ~new_n48072_ & new_n48260_;
  assign new_n48262_ = ~new_n48259_ & ~new_n48261_;
  assign new_n48263_ = ~\b[32]  & ~new_n48262_;
  assign new_n48264_ = ~new_n47556_ & new_n47952_;
  assign new_n48265_ = ~new_n47948_ & new_n48264_;
  assign new_n48266_ = ~new_n47949_ & ~new_n47952_;
  assign new_n48267_ = ~new_n48265_ & ~new_n48266_;
  assign new_n48268_ = ~new_n48074_ & ~new_n48267_;
  assign new_n48269_ = ~new_n47546_ & ~new_n48073_;
  assign new_n48270_ = ~new_n48072_ & new_n48269_;
  assign new_n48271_ = ~new_n48268_ & ~new_n48270_;
  assign new_n48272_ = ~\b[31]  & ~new_n48271_;
  assign new_n48273_ = ~new_n47565_ & new_n47947_;
  assign new_n48274_ = ~new_n47943_ & new_n48273_;
  assign new_n48275_ = ~new_n47944_ & ~new_n47947_;
  assign new_n48276_ = ~new_n48274_ & ~new_n48275_;
  assign new_n48277_ = ~new_n48074_ & ~new_n48276_;
  assign new_n48278_ = ~new_n47555_ & ~new_n48073_;
  assign new_n48279_ = ~new_n48072_ & new_n48278_;
  assign new_n48280_ = ~new_n48277_ & ~new_n48279_;
  assign new_n48281_ = ~\b[30]  & ~new_n48280_;
  assign new_n48282_ = ~new_n47574_ & new_n47942_;
  assign new_n48283_ = ~new_n47938_ & new_n48282_;
  assign new_n48284_ = ~new_n47939_ & ~new_n47942_;
  assign new_n48285_ = ~new_n48283_ & ~new_n48284_;
  assign new_n48286_ = ~new_n48074_ & ~new_n48285_;
  assign new_n48287_ = ~new_n47564_ & ~new_n48073_;
  assign new_n48288_ = ~new_n48072_ & new_n48287_;
  assign new_n48289_ = ~new_n48286_ & ~new_n48288_;
  assign new_n48290_ = ~\b[29]  & ~new_n48289_;
  assign new_n48291_ = ~new_n47583_ & new_n47937_;
  assign new_n48292_ = ~new_n47933_ & new_n48291_;
  assign new_n48293_ = ~new_n47934_ & ~new_n47937_;
  assign new_n48294_ = ~new_n48292_ & ~new_n48293_;
  assign new_n48295_ = ~new_n48074_ & ~new_n48294_;
  assign new_n48296_ = ~new_n47573_ & ~new_n48073_;
  assign new_n48297_ = ~new_n48072_ & new_n48296_;
  assign new_n48298_ = ~new_n48295_ & ~new_n48297_;
  assign new_n48299_ = ~\b[28]  & ~new_n48298_;
  assign new_n48300_ = ~new_n47592_ & new_n47932_;
  assign new_n48301_ = ~new_n47928_ & new_n48300_;
  assign new_n48302_ = ~new_n47929_ & ~new_n47932_;
  assign new_n48303_ = ~new_n48301_ & ~new_n48302_;
  assign new_n48304_ = ~new_n48074_ & ~new_n48303_;
  assign new_n48305_ = ~new_n47582_ & ~new_n48073_;
  assign new_n48306_ = ~new_n48072_ & new_n48305_;
  assign new_n48307_ = ~new_n48304_ & ~new_n48306_;
  assign new_n48308_ = ~\b[27]  & ~new_n48307_;
  assign new_n48309_ = ~new_n47601_ & new_n47927_;
  assign new_n48310_ = ~new_n47923_ & new_n48309_;
  assign new_n48311_ = ~new_n47924_ & ~new_n47927_;
  assign new_n48312_ = ~new_n48310_ & ~new_n48311_;
  assign new_n48313_ = ~new_n48074_ & ~new_n48312_;
  assign new_n48314_ = ~new_n47591_ & ~new_n48073_;
  assign new_n48315_ = ~new_n48072_ & new_n48314_;
  assign new_n48316_ = ~new_n48313_ & ~new_n48315_;
  assign new_n48317_ = ~\b[26]  & ~new_n48316_;
  assign new_n48318_ = ~new_n47610_ & new_n47922_;
  assign new_n48319_ = ~new_n47918_ & new_n48318_;
  assign new_n48320_ = ~new_n47919_ & ~new_n47922_;
  assign new_n48321_ = ~new_n48319_ & ~new_n48320_;
  assign new_n48322_ = ~new_n48074_ & ~new_n48321_;
  assign new_n48323_ = ~new_n47600_ & ~new_n48073_;
  assign new_n48324_ = ~new_n48072_ & new_n48323_;
  assign new_n48325_ = ~new_n48322_ & ~new_n48324_;
  assign new_n48326_ = ~\b[25]  & ~new_n48325_;
  assign new_n48327_ = ~new_n47619_ & new_n47917_;
  assign new_n48328_ = ~new_n47913_ & new_n48327_;
  assign new_n48329_ = ~new_n47914_ & ~new_n47917_;
  assign new_n48330_ = ~new_n48328_ & ~new_n48329_;
  assign new_n48331_ = ~new_n48074_ & ~new_n48330_;
  assign new_n48332_ = ~new_n47609_ & ~new_n48073_;
  assign new_n48333_ = ~new_n48072_ & new_n48332_;
  assign new_n48334_ = ~new_n48331_ & ~new_n48333_;
  assign new_n48335_ = ~\b[24]  & ~new_n48334_;
  assign new_n48336_ = ~new_n47628_ & new_n47912_;
  assign new_n48337_ = ~new_n47908_ & new_n48336_;
  assign new_n48338_ = ~new_n47909_ & ~new_n47912_;
  assign new_n48339_ = ~new_n48337_ & ~new_n48338_;
  assign new_n48340_ = ~new_n48074_ & ~new_n48339_;
  assign new_n48341_ = ~new_n47618_ & ~new_n48073_;
  assign new_n48342_ = ~new_n48072_ & new_n48341_;
  assign new_n48343_ = ~new_n48340_ & ~new_n48342_;
  assign new_n48344_ = ~\b[23]  & ~new_n48343_;
  assign new_n48345_ = ~new_n47637_ & new_n47907_;
  assign new_n48346_ = ~new_n47903_ & new_n48345_;
  assign new_n48347_ = ~new_n47904_ & ~new_n47907_;
  assign new_n48348_ = ~new_n48346_ & ~new_n48347_;
  assign new_n48349_ = ~new_n48074_ & ~new_n48348_;
  assign new_n48350_ = ~new_n47627_ & ~new_n48073_;
  assign new_n48351_ = ~new_n48072_ & new_n48350_;
  assign new_n48352_ = ~new_n48349_ & ~new_n48351_;
  assign new_n48353_ = ~\b[22]  & ~new_n48352_;
  assign new_n48354_ = ~new_n47646_ & new_n47902_;
  assign new_n48355_ = ~new_n47898_ & new_n48354_;
  assign new_n48356_ = ~new_n47899_ & ~new_n47902_;
  assign new_n48357_ = ~new_n48355_ & ~new_n48356_;
  assign new_n48358_ = ~new_n48074_ & ~new_n48357_;
  assign new_n48359_ = ~new_n47636_ & ~new_n48073_;
  assign new_n48360_ = ~new_n48072_ & new_n48359_;
  assign new_n48361_ = ~new_n48358_ & ~new_n48360_;
  assign new_n48362_ = ~\b[21]  & ~new_n48361_;
  assign new_n48363_ = ~new_n47655_ & new_n47897_;
  assign new_n48364_ = ~new_n47893_ & new_n48363_;
  assign new_n48365_ = ~new_n47894_ & ~new_n47897_;
  assign new_n48366_ = ~new_n48364_ & ~new_n48365_;
  assign new_n48367_ = ~new_n48074_ & ~new_n48366_;
  assign new_n48368_ = ~new_n47645_ & ~new_n48073_;
  assign new_n48369_ = ~new_n48072_ & new_n48368_;
  assign new_n48370_ = ~new_n48367_ & ~new_n48369_;
  assign new_n48371_ = ~\b[20]  & ~new_n48370_;
  assign new_n48372_ = ~new_n47664_ & new_n47892_;
  assign new_n48373_ = ~new_n47888_ & new_n48372_;
  assign new_n48374_ = ~new_n47889_ & ~new_n47892_;
  assign new_n48375_ = ~new_n48373_ & ~new_n48374_;
  assign new_n48376_ = ~new_n48074_ & ~new_n48375_;
  assign new_n48377_ = ~new_n47654_ & ~new_n48073_;
  assign new_n48378_ = ~new_n48072_ & new_n48377_;
  assign new_n48379_ = ~new_n48376_ & ~new_n48378_;
  assign new_n48380_ = ~\b[19]  & ~new_n48379_;
  assign new_n48381_ = ~new_n47673_ & new_n47887_;
  assign new_n48382_ = ~new_n47883_ & new_n48381_;
  assign new_n48383_ = ~new_n47884_ & ~new_n47887_;
  assign new_n48384_ = ~new_n48382_ & ~new_n48383_;
  assign new_n48385_ = ~new_n48074_ & ~new_n48384_;
  assign new_n48386_ = ~new_n47663_ & ~new_n48073_;
  assign new_n48387_ = ~new_n48072_ & new_n48386_;
  assign new_n48388_ = ~new_n48385_ & ~new_n48387_;
  assign new_n48389_ = ~\b[18]  & ~new_n48388_;
  assign new_n48390_ = ~new_n47682_ & new_n47882_;
  assign new_n48391_ = ~new_n47878_ & new_n48390_;
  assign new_n48392_ = ~new_n47879_ & ~new_n47882_;
  assign new_n48393_ = ~new_n48391_ & ~new_n48392_;
  assign new_n48394_ = ~new_n48074_ & ~new_n48393_;
  assign new_n48395_ = ~new_n47672_ & ~new_n48073_;
  assign new_n48396_ = ~new_n48072_ & new_n48395_;
  assign new_n48397_ = ~new_n48394_ & ~new_n48396_;
  assign new_n48398_ = ~\b[17]  & ~new_n48397_;
  assign new_n48399_ = ~new_n47691_ & new_n47877_;
  assign new_n48400_ = ~new_n47873_ & new_n48399_;
  assign new_n48401_ = ~new_n47874_ & ~new_n47877_;
  assign new_n48402_ = ~new_n48400_ & ~new_n48401_;
  assign new_n48403_ = ~new_n48074_ & ~new_n48402_;
  assign new_n48404_ = ~new_n47681_ & ~new_n48073_;
  assign new_n48405_ = ~new_n48072_ & new_n48404_;
  assign new_n48406_ = ~new_n48403_ & ~new_n48405_;
  assign new_n48407_ = ~\b[16]  & ~new_n48406_;
  assign new_n48408_ = ~new_n47700_ & new_n47872_;
  assign new_n48409_ = ~new_n47868_ & new_n48408_;
  assign new_n48410_ = ~new_n47869_ & ~new_n47872_;
  assign new_n48411_ = ~new_n48409_ & ~new_n48410_;
  assign new_n48412_ = ~new_n48074_ & ~new_n48411_;
  assign new_n48413_ = ~new_n47690_ & ~new_n48073_;
  assign new_n48414_ = ~new_n48072_ & new_n48413_;
  assign new_n48415_ = ~new_n48412_ & ~new_n48414_;
  assign new_n48416_ = ~\b[15]  & ~new_n48415_;
  assign new_n48417_ = ~new_n47709_ & new_n47867_;
  assign new_n48418_ = ~new_n47863_ & new_n48417_;
  assign new_n48419_ = ~new_n47864_ & ~new_n47867_;
  assign new_n48420_ = ~new_n48418_ & ~new_n48419_;
  assign new_n48421_ = ~new_n48074_ & ~new_n48420_;
  assign new_n48422_ = ~new_n47699_ & ~new_n48073_;
  assign new_n48423_ = ~new_n48072_ & new_n48422_;
  assign new_n48424_ = ~new_n48421_ & ~new_n48423_;
  assign new_n48425_ = ~\b[14]  & ~new_n48424_;
  assign new_n48426_ = ~new_n47718_ & new_n47862_;
  assign new_n48427_ = ~new_n47858_ & new_n48426_;
  assign new_n48428_ = ~new_n47859_ & ~new_n47862_;
  assign new_n48429_ = ~new_n48427_ & ~new_n48428_;
  assign new_n48430_ = ~new_n48074_ & ~new_n48429_;
  assign new_n48431_ = ~new_n47708_ & ~new_n48073_;
  assign new_n48432_ = ~new_n48072_ & new_n48431_;
  assign new_n48433_ = ~new_n48430_ & ~new_n48432_;
  assign new_n48434_ = ~\b[13]  & ~new_n48433_;
  assign new_n48435_ = ~new_n47727_ & new_n47857_;
  assign new_n48436_ = ~new_n47853_ & new_n48435_;
  assign new_n48437_ = ~new_n47854_ & ~new_n47857_;
  assign new_n48438_ = ~new_n48436_ & ~new_n48437_;
  assign new_n48439_ = ~new_n48074_ & ~new_n48438_;
  assign new_n48440_ = ~new_n47717_ & ~new_n48073_;
  assign new_n48441_ = ~new_n48072_ & new_n48440_;
  assign new_n48442_ = ~new_n48439_ & ~new_n48441_;
  assign new_n48443_ = ~\b[12]  & ~new_n48442_;
  assign new_n48444_ = ~new_n47736_ & new_n47852_;
  assign new_n48445_ = ~new_n47848_ & new_n48444_;
  assign new_n48446_ = ~new_n47849_ & ~new_n47852_;
  assign new_n48447_ = ~new_n48445_ & ~new_n48446_;
  assign new_n48448_ = ~new_n48074_ & ~new_n48447_;
  assign new_n48449_ = ~new_n47726_ & ~new_n48073_;
  assign new_n48450_ = ~new_n48072_ & new_n48449_;
  assign new_n48451_ = ~new_n48448_ & ~new_n48450_;
  assign new_n48452_ = ~\b[11]  & ~new_n48451_;
  assign new_n48453_ = ~new_n47745_ & new_n47847_;
  assign new_n48454_ = ~new_n47843_ & new_n48453_;
  assign new_n48455_ = ~new_n47844_ & ~new_n47847_;
  assign new_n48456_ = ~new_n48454_ & ~new_n48455_;
  assign new_n48457_ = ~new_n48074_ & ~new_n48456_;
  assign new_n48458_ = ~new_n47735_ & ~new_n48073_;
  assign new_n48459_ = ~new_n48072_ & new_n48458_;
  assign new_n48460_ = ~new_n48457_ & ~new_n48459_;
  assign new_n48461_ = ~\b[10]  & ~new_n48460_;
  assign new_n48462_ = ~new_n47754_ & new_n47842_;
  assign new_n48463_ = ~new_n47838_ & new_n48462_;
  assign new_n48464_ = ~new_n47839_ & ~new_n47842_;
  assign new_n48465_ = ~new_n48463_ & ~new_n48464_;
  assign new_n48466_ = ~new_n48074_ & ~new_n48465_;
  assign new_n48467_ = ~new_n47744_ & ~new_n48073_;
  assign new_n48468_ = ~new_n48072_ & new_n48467_;
  assign new_n48469_ = ~new_n48466_ & ~new_n48468_;
  assign new_n48470_ = ~\b[9]  & ~new_n48469_;
  assign new_n48471_ = ~new_n47763_ & new_n47837_;
  assign new_n48472_ = ~new_n47833_ & new_n48471_;
  assign new_n48473_ = ~new_n47834_ & ~new_n47837_;
  assign new_n48474_ = ~new_n48472_ & ~new_n48473_;
  assign new_n48475_ = ~new_n48074_ & ~new_n48474_;
  assign new_n48476_ = ~new_n47753_ & ~new_n48073_;
  assign new_n48477_ = ~new_n48072_ & new_n48476_;
  assign new_n48478_ = ~new_n48475_ & ~new_n48477_;
  assign new_n48479_ = ~\b[8]  & ~new_n48478_;
  assign new_n48480_ = ~new_n47772_ & new_n47832_;
  assign new_n48481_ = ~new_n47828_ & new_n48480_;
  assign new_n48482_ = ~new_n47829_ & ~new_n47832_;
  assign new_n48483_ = ~new_n48481_ & ~new_n48482_;
  assign new_n48484_ = ~new_n48074_ & ~new_n48483_;
  assign new_n48485_ = ~new_n47762_ & ~new_n48073_;
  assign new_n48486_ = ~new_n48072_ & new_n48485_;
  assign new_n48487_ = ~new_n48484_ & ~new_n48486_;
  assign new_n48488_ = ~\b[7]  & ~new_n48487_;
  assign new_n48489_ = ~new_n47781_ & new_n47827_;
  assign new_n48490_ = ~new_n47823_ & new_n48489_;
  assign new_n48491_ = ~new_n47824_ & ~new_n47827_;
  assign new_n48492_ = ~new_n48490_ & ~new_n48491_;
  assign new_n48493_ = ~new_n48074_ & ~new_n48492_;
  assign new_n48494_ = ~new_n47771_ & ~new_n48073_;
  assign new_n48495_ = ~new_n48072_ & new_n48494_;
  assign new_n48496_ = ~new_n48493_ & ~new_n48495_;
  assign new_n48497_ = ~\b[6]  & ~new_n48496_;
  assign new_n48498_ = ~new_n47790_ & new_n47822_;
  assign new_n48499_ = ~new_n47818_ & new_n48498_;
  assign new_n48500_ = ~new_n47819_ & ~new_n47822_;
  assign new_n48501_ = ~new_n48499_ & ~new_n48500_;
  assign new_n48502_ = ~new_n48074_ & ~new_n48501_;
  assign new_n48503_ = ~new_n47780_ & ~new_n48073_;
  assign new_n48504_ = ~new_n48072_ & new_n48503_;
  assign new_n48505_ = ~new_n48502_ & ~new_n48504_;
  assign new_n48506_ = ~\b[5]  & ~new_n48505_;
  assign new_n48507_ = ~new_n47798_ & new_n47817_;
  assign new_n48508_ = ~new_n47813_ & new_n48507_;
  assign new_n48509_ = ~new_n47814_ & ~new_n47817_;
  assign new_n48510_ = ~new_n48508_ & ~new_n48509_;
  assign new_n48511_ = ~new_n48074_ & ~new_n48510_;
  assign new_n48512_ = ~new_n47789_ & ~new_n48073_;
  assign new_n48513_ = ~new_n48072_ & new_n48512_;
  assign new_n48514_ = ~new_n48511_ & ~new_n48513_;
  assign new_n48515_ = ~\b[4]  & ~new_n48514_;
  assign new_n48516_ = ~new_n47808_ & new_n47812_;
  assign new_n48517_ = ~new_n47807_ & new_n48516_;
  assign new_n48518_ = ~new_n47809_ & ~new_n47812_;
  assign new_n48519_ = ~new_n48517_ & ~new_n48518_;
  assign new_n48520_ = ~new_n48074_ & ~new_n48519_;
  assign new_n48521_ = ~new_n47797_ & ~new_n48073_;
  assign new_n48522_ = ~new_n48072_ & new_n48521_;
  assign new_n48523_ = ~new_n48520_ & ~new_n48522_;
  assign new_n48524_ = ~\b[3]  & ~new_n48523_;
  assign new_n48525_ = new_n19767_ & ~new_n47805_;
  assign new_n48526_ = ~new_n47803_ & new_n48525_;
  assign new_n48527_ = ~new_n47807_ & ~new_n48526_;
  assign new_n48528_ = ~new_n48074_ & new_n48527_;
  assign new_n48529_ = ~new_n47802_ & ~new_n48073_;
  assign new_n48530_ = ~new_n48072_ & new_n48529_;
  assign new_n48531_ = ~new_n48528_ & ~new_n48530_;
  assign new_n48532_ = ~\b[2]  & ~new_n48531_;
  assign new_n48533_ = \b[0]  & ~new_n48074_;
  assign new_n48534_ = \a[11]  & ~new_n48533_;
  assign new_n48535_ = new_n19767_ & ~new_n48074_;
  assign new_n48536_ = ~new_n48534_ & ~new_n48535_;
  assign new_n48537_ = \b[1]  & ~new_n48536_;
  assign new_n48538_ = ~\b[1]  & ~new_n48535_;
  assign new_n48539_ = ~new_n48534_ & new_n48538_;
  assign new_n48540_ = ~new_n48537_ & ~new_n48539_;
  assign new_n48541_ = ~new_n20502_ & ~new_n48540_;
  assign new_n48542_ = ~\b[1]  & ~new_n48536_;
  assign new_n48543_ = ~new_n48541_ & ~new_n48542_;
  assign new_n48544_ = \b[2]  & ~new_n48530_;
  assign new_n48545_ = ~new_n48528_ & new_n48544_;
  assign new_n48546_ = ~new_n48532_ & ~new_n48545_;
  assign new_n48547_ = ~new_n48543_ & new_n48546_;
  assign new_n48548_ = ~new_n48532_ & ~new_n48547_;
  assign new_n48549_ = \b[3]  & ~new_n48522_;
  assign new_n48550_ = ~new_n48520_ & new_n48549_;
  assign new_n48551_ = ~new_n48524_ & ~new_n48550_;
  assign new_n48552_ = ~new_n48548_ & new_n48551_;
  assign new_n48553_ = ~new_n48524_ & ~new_n48552_;
  assign new_n48554_ = \b[4]  & ~new_n48513_;
  assign new_n48555_ = ~new_n48511_ & new_n48554_;
  assign new_n48556_ = ~new_n48515_ & ~new_n48555_;
  assign new_n48557_ = ~new_n48553_ & new_n48556_;
  assign new_n48558_ = ~new_n48515_ & ~new_n48557_;
  assign new_n48559_ = \b[5]  & ~new_n48504_;
  assign new_n48560_ = ~new_n48502_ & new_n48559_;
  assign new_n48561_ = ~new_n48506_ & ~new_n48560_;
  assign new_n48562_ = ~new_n48558_ & new_n48561_;
  assign new_n48563_ = ~new_n48506_ & ~new_n48562_;
  assign new_n48564_ = \b[6]  & ~new_n48495_;
  assign new_n48565_ = ~new_n48493_ & new_n48564_;
  assign new_n48566_ = ~new_n48497_ & ~new_n48565_;
  assign new_n48567_ = ~new_n48563_ & new_n48566_;
  assign new_n48568_ = ~new_n48497_ & ~new_n48567_;
  assign new_n48569_ = \b[7]  & ~new_n48486_;
  assign new_n48570_ = ~new_n48484_ & new_n48569_;
  assign new_n48571_ = ~new_n48488_ & ~new_n48570_;
  assign new_n48572_ = ~new_n48568_ & new_n48571_;
  assign new_n48573_ = ~new_n48488_ & ~new_n48572_;
  assign new_n48574_ = \b[8]  & ~new_n48477_;
  assign new_n48575_ = ~new_n48475_ & new_n48574_;
  assign new_n48576_ = ~new_n48479_ & ~new_n48575_;
  assign new_n48577_ = ~new_n48573_ & new_n48576_;
  assign new_n48578_ = ~new_n48479_ & ~new_n48577_;
  assign new_n48579_ = \b[9]  & ~new_n48468_;
  assign new_n48580_ = ~new_n48466_ & new_n48579_;
  assign new_n48581_ = ~new_n48470_ & ~new_n48580_;
  assign new_n48582_ = ~new_n48578_ & new_n48581_;
  assign new_n48583_ = ~new_n48470_ & ~new_n48582_;
  assign new_n48584_ = \b[10]  & ~new_n48459_;
  assign new_n48585_ = ~new_n48457_ & new_n48584_;
  assign new_n48586_ = ~new_n48461_ & ~new_n48585_;
  assign new_n48587_ = ~new_n48583_ & new_n48586_;
  assign new_n48588_ = ~new_n48461_ & ~new_n48587_;
  assign new_n48589_ = \b[11]  & ~new_n48450_;
  assign new_n48590_ = ~new_n48448_ & new_n48589_;
  assign new_n48591_ = ~new_n48452_ & ~new_n48590_;
  assign new_n48592_ = ~new_n48588_ & new_n48591_;
  assign new_n48593_ = ~new_n48452_ & ~new_n48592_;
  assign new_n48594_ = \b[12]  & ~new_n48441_;
  assign new_n48595_ = ~new_n48439_ & new_n48594_;
  assign new_n48596_ = ~new_n48443_ & ~new_n48595_;
  assign new_n48597_ = ~new_n48593_ & new_n48596_;
  assign new_n48598_ = ~new_n48443_ & ~new_n48597_;
  assign new_n48599_ = \b[13]  & ~new_n48432_;
  assign new_n48600_ = ~new_n48430_ & new_n48599_;
  assign new_n48601_ = ~new_n48434_ & ~new_n48600_;
  assign new_n48602_ = ~new_n48598_ & new_n48601_;
  assign new_n48603_ = ~new_n48434_ & ~new_n48602_;
  assign new_n48604_ = \b[14]  & ~new_n48423_;
  assign new_n48605_ = ~new_n48421_ & new_n48604_;
  assign new_n48606_ = ~new_n48425_ & ~new_n48605_;
  assign new_n48607_ = ~new_n48603_ & new_n48606_;
  assign new_n48608_ = ~new_n48425_ & ~new_n48607_;
  assign new_n48609_ = \b[15]  & ~new_n48414_;
  assign new_n48610_ = ~new_n48412_ & new_n48609_;
  assign new_n48611_ = ~new_n48416_ & ~new_n48610_;
  assign new_n48612_ = ~new_n48608_ & new_n48611_;
  assign new_n48613_ = ~new_n48416_ & ~new_n48612_;
  assign new_n48614_ = \b[16]  & ~new_n48405_;
  assign new_n48615_ = ~new_n48403_ & new_n48614_;
  assign new_n48616_ = ~new_n48407_ & ~new_n48615_;
  assign new_n48617_ = ~new_n48613_ & new_n48616_;
  assign new_n48618_ = ~new_n48407_ & ~new_n48617_;
  assign new_n48619_ = \b[17]  & ~new_n48396_;
  assign new_n48620_ = ~new_n48394_ & new_n48619_;
  assign new_n48621_ = ~new_n48398_ & ~new_n48620_;
  assign new_n48622_ = ~new_n48618_ & new_n48621_;
  assign new_n48623_ = ~new_n48398_ & ~new_n48622_;
  assign new_n48624_ = \b[18]  & ~new_n48387_;
  assign new_n48625_ = ~new_n48385_ & new_n48624_;
  assign new_n48626_ = ~new_n48389_ & ~new_n48625_;
  assign new_n48627_ = ~new_n48623_ & new_n48626_;
  assign new_n48628_ = ~new_n48389_ & ~new_n48627_;
  assign new_n48629_ = \b[19]  & ~new_n48378_;
  assign new_n48630_ = ~new_n48376_ & new_n48629_;
  assign new_n48631_ = ~new_n48380_ & ~new_n48630_;
  assign new_n48632_ = ~new_n48628_ & new_n48631_;
  assign new_n48633_ = ~new_n48380_ & ~new_n48632_;
  assign new_n48634_ = \b[20]  & ~new_n48369_;
  assign new_n48635_ = ~new_n48367_ & new_n48634_;
  assign new_n48636_ = ~new_n48371_ & ~new_n48635_;
  assign new_n48637_ = ~new_n48633_ & new_n48636_;
  assign new_n48638_ = ~new_n48371_ & ~new_n48637_;
  assign new_n48639_ = \b[21]  & ~new_n48360_;
  assign new_n48640_ = ~new_n48358_ & new_n48639_;
  assign new_n48641_ = ~new_n48362_ & ~new_n48640_;
  assign new_n48642_ = ~new_n48638_ & new_n48641_;
  assign new_n48643_ = ~new_n48362_ & ~new_n48642_;
  assign new_n48644_ = \b[22]  & ~new_n48351_;
  assign new_n48645_ = ~new_n48349_ & new_n48644_;
  assign new_n48646_ = ~new_n48353_ & ~new_n48645_;
  assign new_n48647_ = ~new_n48643_ & new_n48646_;
  assign new_n48648_ = ~new_n48353_ & ~new_n48647_;
  assign new_n48649_ = \b[23]  & ~new_n48342_;
  assign new_n48650_ = ~new_n48340_ & new_n48649_;
  assign new_n48651_ = ~new_n48344_ & ~new_n48650_;
  assign new_n48652_ = ~new_n48648_ & new_n48651_;
  assign new_n48653_ = ~new_n48344_ & ~new_n48652_;
  assign new_n48654_ = \b[24]  & ~new_n48333_;
  assign new_n48655_ = ~new_n48331_ & new_n48654_;
  assign new_n48656_ = ~new_n48335_ & ~new_n48655_;
  assign new_n48657_ = ~new_n48653_ & new_n48656_;
  assign new_n48658_ = ~new_n48335_ & ~new_n48657_;
  assign new_n48659_ = \b[25]  & ~new_n48324_;
  assign new_n48660_ = ~new_n48322_ & new_n48659_;
  assign new_n48661_ = ~new_n48326_ & ~new_n48660_;
  assign new_n48662_ = ~new_n48658_ & new_n48661_;
  assign new_n48663_ = ~new_n48326_ & ~new_n48662_;
  assign new_n48664_ = \b[26]  & ~new_n48315_;
  assign new_n48665_ = ~new_n48313_ & new_n48664_;
  assign new_n48666_ = ~new_n48317_ & ~new_n48665_;
  assign new_n48667_ = ~new_n48663_ & new_n48666_;
  assign new_n48668_ = ~new_n48317_ & ~new_n48667_;
  assign new_n48669_ = \b[27]  & ~new_n48306_;
  assign new_n48670_ = ~new_n48304_ & new_n48669_;
  assign new_n48671_ = ~new_n48308_ & ~new_n48670_;
  assign new_n48672_ = ~new_n48668_ & new_n48671_;
  assign new_n48673_ = ~new_n48308_ & ~new_n48672_;
  assign new_n48674_ = \b[28]  & ~new_n48297_;
  assign new_n48675_ = ~new_n48295_ & new_n48674_;
  assign new_n48676_ = ~new_n48299_ & ~new_n48675_;
  assign new_n48677_ = ~new_n48673_ & new_n48676_;
  assign new_n48678_ = ~new_n48299_ & ~new_n48677_;
  assign new_n48679_ = \b[29]  & ~new_n48288_;
  assign new_n48680_ = ~new_n48286_ & new_n48679_;
  assign new_n48681_ = ~new_n48290_ & ~new_n48680_;
  assign new_n48682_ = ~new_n48678_ & new_n48681_;
  assign new_n48683_ = ~new_n48290_ & ~new_n48682_;
  assign new_n48684_ = \b[30]  & ~new_n48279_;
  assign new_n48685_ = ~new_n48277_ & new_n48684_;
  assign new_n48686_ = ~new_n48281_ & ~new_n48685_;
  assign new_n48687_ = ~new_n48683_ & new_n48686_;
  assign new_n48688_ = ~new_n48281_ & ~new_n48687_;
  assign new_n48689_ = \b[31]  & ~new_n48270_;
  assign new_n48690_ = ~new_n48268_ & new_n48689_;
  assign new_n48691_ = ~new_n48272_ & ~new_n48690_;
  assign new_n48692_ = ~new_n48688_ & new_n48691_;
  assign new_n48693_ = ~new_n48272_ & ~new_n48692_;
  assign new_n48694_ = \b[32]  & ~new_n48261_;
  assign new_n48695_ = ~new_n48259_ & new_n48694_;
  assign new_n48696_ = ~new_n48263_ & ~new_n48695_;
  assign new_n48697_ = ~new_n48693_ & new_n48696_;
  assign new_n48698_ = ~new_n48263_ & ~new_n48697_;
  assign new_n48699_ = \b[33]  & ~new_n48252_;
  assign new_n48700_ = ~new_n48250_ & new_n48699_;
  assign new_n48701_ = ~new_n48254_ & ~new_n48700_;
  assign new_n48702_ = ~new_n48698_ & new_n48701_;
  assign new_n48703_ = ~new_n48254_ & ~new_n48702_;
  assign new_n48704_ = \b[34]  & ~new_n48243_;
  assign new_n48705_ = ~new_n48241_ & new_n48704_;
  assign new_n48706_ = ~new_n48245_ & ~new_n48705_;
  assign new_n48707_ = ~new_n48703_ & new_n48706_;
  assign new_n48708_ = ~new_n48245_ & ~new_n48707_;
  assign new_n48709_ = \b[35]  & ~new_n48234_;
  assign new_n48710_ = ~new_n48232_ & new_n48709_;
  assign new_n48711_ = ~new_n48236_ & ~new_n48710_;
  assign new_n48712_ = ~new_n48708_ & new_n48711_;
  assign new_n48713_ = ~new_n48236_ & ~new_n48712_;
  assign new_n48714_ = \b[36]  & ~new_n48225_;
  assign new_n48715_ = ~new_n48223_ & new_n48714_;
  assign new_n48716_ = ~new_n48227_ & ~new_n48715_;
  assign new_n48717_ = ~new_n48713_ & new_n48716_;
  assign new_n48718_ = ~new_n48227_ & ~new_n48717_;
  assign new_n48719_ = \b[37]  & ~new_n48216_;
  assign new_n48720_ = ~new_n48214_ & new_n48719_;
  assign new_n48721_ = ~new_n48218_ & ~new_n48720_;
  assign new_n48722_ = ~new_n48718_ & new_n48721_;
  assign new_n48723_ = ~new_n48218_ & ~new_n48722_;
  assign new_n48724_ = \b[38]  & ~new_n48207_;
  assign new_n48725_ = ~new_n48205_ & new_n48724_;
  assign new_n48726_ = ~new_n48209_ & ~new_n48725_;
  assign new_n48727_ = ~new_n48723_ & new_n48726_;
  assign new_n48728_ = ~new_n48209_ & ~new_n48727_;
  assign new_n48729_ = \b[39]  & ~new_n48198_;
  assign new_n48730_ = ~new_n48196_ & new_n48729_;
  assign new_n48731_ = ~new_n48200_ & ~new_n48730_;
  assign new_n48732_ = ~new_n48728_ & new_n48731_;
  assign new_n48733_ = ~new_n48200_ & ~new_n48732_;
  assign new_n48734_ = \b[40]  & ~new_n48189_;
  assign new_n48735_ = ~new_n48187_ & new_n48734_;
  assign new_n48736_ = ~new_n48191_ & ~new_n48735_;
  assign new_n48737_ = ~new_n48733_ & new_n48736_;
  assign new_n48738_ = ~new_n48191_ & ~new_n48737_;
  assign new_n48739_ = \b[41]  & ~new_n48180_;
  assign new_n48740_ = ~new_n48178_ & new_n48739_;
  assign new_n48741_ = ~new_n48182_ & ~new_n48740_;
  assign new_n48742_ = ~new_n48738_ & new_n48741_;
  assign new_n48743_ = ~new_n48182_ & ~new_n48742_;
  assign new_n48744_ = \b[42]  & ~new_n48171_;
  assign new_n48745_ = ~new_n48169_ & new_n48744_;
  assign new_n48746_ = ~new_n48173_ & ~new_n48745_;
  assign new_n48747_ = ~new_n48743_ & new_n48746_;
  assign new_n48748_ = ~new_n48173_ & ~new_n48747_;
  assign new_n48749_ = \b[43]  & ~new_n48162_;
  assign new_n48750_ = ~new_n48160_ & new_n48749_;
  assign new_n48751_ = ~new_n48164_ & ~new_n48750_;
  assign new_n48752_ = ~new_n48748_ & new_n48751_;
  assign new_n48753_ = ~new_n48164_ & ~new_n48752_;
  assign new_n48754_ = \b[44]  & ~new_n48153_;
  assign new_n48755_ = ~new_n48151_ & new_n48754_;
  assign new_n48756_ = ~new_n48155_ & ~new_n48755_;
  assign new_n48757_ = ~new_n48753_ & new_n48756_;
  assign new_n48758_ = ~new_n48155_ & ~new_n48757_;
  assign new_n48759_ = \b[45]  & ~new_n48144_;
  assign new_n48760_ = ~new_n48142_ & new_n48759_;
  assign new_n48761_ = ~new_n48146_ & ~new_n48760_;
  assign new_n48762_ = ~new_n48758_ & new_n48761_;
  assign new_n48763_ = ~new_n48146_ & ~new_n48762_;
  assign new_n48764_ = \b[46]  & ~new_n48135_;
  assign new_n48765_ = ~new_n48133_ & new_n48764_;
  assign new_n48766_ = ~new_n48137_ & ~new_n48765_;
  assign new_n48767_ = ~new_n48763_ & new_n48766_;
  assign new_n48768_ = ~new_n48137_ & ~new_n48767_;
  assign new_n48769_ = \b[47]  & ~new_n48126_;
  assign new_n48770_ = ~new_n48124_ & new_n48769_;
  assign new_n48771_ = ~new_n48128_ & ~new_n48770_;
  assign new_n48772_ = ~new_n48768_ & new_n48771_;
  assign new_n48773_ = ~new_n48128_ & ~new_n48772_;
  assign new_n48774_ = \b[48]  & ~new_n48117_;
  assign new_n48775_ = ~new_n48115_ & new_n48774_;
  assign new_n48776_ = ~new_n48119_ & ~new_n48775_;
  assign new_n48777_ = ~new_n48773_ & new_n48776_;
  assign new_n48778_ = ~new_n48119_ & ~new_n48777_;
  assign new_n48779_ = \b[49]  & ~new_n48108_;
  assign new_n48780_ = ~new_n48106_ & new_n48779_;
  assign new_n48781_ = ~new_n48110_ & ~new_n48780_;
  assign new_n48782_ = ~new_n48778_ & new_n48781_;
  assign new_n48783_ = ~new_n48110_ & ~new_n48782_;
  assign new_n48784_ = \b[50]  & ~new_n48099_;
  assign new_n48785_ = ~new_n48097_ & new_n48784_;
  assign new_n48786_ = ~new_n48101_ & ~new_n48785_;
  assign new_n48787_ = ~new_n48783_ & new_n48786_;
  assign new_n48788_ = ~new_n48101_ & ~new_n48787_;
  assign new_n48789_ = \b[51]  & ~new_n48090_;
  assign new_n48790_ = ~new_n48088_ & new_n48789_;
  assign new_n48791_ = ~new_n48092_ & ~new_n48790_;
  assign new_n48792_ = ~new_n48788_ & new_n48791_;
  assign new_n48793_ = ~new_n48092_ & ~new_n48792_;
  assign new_n48794_ = \b[52]  & ~new_n48081_;
  assign new_n48795_ = ~new_n48079_ & new_n48794_;
  assign new_n48796_ = ~new_n48083_ & ~new_n48795_;
  assign new_n48797_ = ~new_n48793_ & new_n48796_;
  assign new_n48798_ = ~new_n48083_ & ~new_n48797_;
  assign new_n48799_ = ~new_n47358_ & ~new_n48069_;
  assign new_n48800_ = ~new_n48067_ & new_n48799_;
  assign new_n48801_ = ~new_n48058_ & new_n48800_;
  assign new_n48802_ = ~new_n48067_ & ~new_n48069_;
  assign new_n48803_ = ~new_n48059_ & ~new_n48802_;
  assign new_n48804_ = ~new_n48801_ & ~new_n48803_;
  assign new_n48805_ = ~new_n48074_ & ~new_n48804_;
  assign new_n48806_ = ~new_n48066_ & ~new_n48073_;
  assign new_n48807_ = ~new_n48072_ & new_n48806_;
  assign new_n48808_ = ~new_n48805_ & ~new_n48807_;
  assign new_n48809_ = ~\b[53]  & ~new_n48808_;
  assign new_n48810_ = \b[53]  & ~new_n48807_;
  assign new_n48811_ = ~new_n48805_ & new_n48810_;
  assign new_n48812_ = new_n20775_ & ~new_n48811_;
  assign new_n48813_ = ~new_n48809_ & new_n48812_;
  assign new_n48814_ = ~new_n48798_ & new_n48813_;
  assign new_n48815_ = new_n595_ & ~new_n48808_;
  assign new_n48816_ = ~new_n48814_ & ~new_n48815_;
  assign new_n48817_ = ~new_n48092_ & new_n48796_;
  assign new_n48818_ = ~new_n48792_ & new_n48817_;
  assign new_n48819_ = ~new_n48793_ & ~new_n48796_;
  assign new_n48820_ = ~new_n48818_ & ~new_n48819_;
  assign new_n48821_ = ~new_n48816_ & ~new_n48820_;
  assign new_n48822_ = ~new_n48082_ & ~new_n48815_;
  assign new_n48823_ = ~new_n48814_ & new_n48822_;
  assign new_n48824_ = ~new_n48821_ & ~new_n48823_;
  assign new_n48825_ = ~new_n48083_ & ~new_n48811_;
  assign new_n48826_ = ~new_n48809_ & new_n48825_;
  assign new_n48827_ = ~new_n48797_ & new_n48826_;
  assign new_n48828_ = ~new_n48809_ & ~new_n48811_;
  assign new_n48829_ = ~new_n48798_ & ~new_n48828_;
  assign new_n48830_ = ~new_n48827_ & ~new_n48829_;
  assign new_n48831_ = ~new_n48816_ & ~new_n48830_;
  assign new_n48832_ = ~new_n48808_ & ~new_n48815_;
  assign new_n48833_ = ~new_n48814_ & new_n48832_;
  assign new_n48834_ = ~new_n48831_ & ~new_n48833_;
  assign new_n48835_ = ~\b[54]  & ~new_n48834_;
  assign new_n48836_ = ~\b[53]  & ~new_n48824_;
  assign new_n48837_ = ~new_n48101_ & new_n48791_;
  assign new_n48838_ = ~new_n48787_ & new_n48837_;
  assign new_n48839_ = ~new_n48788_ & ~new_n48791_;
  assign new_n48840_ = ~new_n48838_ & ~new_n48839_;
  assign new_n48841_ = ~new_n48816_ & ~new_n48840_;
  assign new_n48842_ = ~new_n48091_ & ~new_n48815_;
  assign new_n48843_ = ~new_n48814_ & new_n48842_;
  assign new_n48844_ = ~new_n48841_ & ~new_n48843_;
  assign new_n48845_ = ~\b[52]  & ~new_n48844_;
  assign new_n48846_ = ~new_n48110_ & new_n48786_;
  assign new_n48847_ = ~new_n48782_ & new_n48846_;
  assign new_n48848_ = ~new_n48783_ & ~new_n48786_;
  assign new_n48849_ = ~new_n48847_ & ~new_n48848_;
  assign new_n48850_ = ~new_n48816_ & ~new_n48849_;
  assign new_n48851_ = ~new_n48100_ & ~new_n48815_;
  assign new_n48852_ = ~new_n48814_ & new_n48851_;
  assign new_n48853_ = ~new_n48850_ & ~new_n48852_;
  assign new_n48854_ = ~\b[51]  & ~new_n48853_;
  assign new_n48855_ = ~new_n48119_ & new_n48781_;
  assign new_n48856_ = ~new_n48777_ & new_n48855_;
  assign new_n48857_ = ~new_n48778_ & ~new_n48781_;
  assign new_n48858_ = ~new_n48856_ & ~new_n48857_;
  assign new_n48859_ = ~new_n48816_ & ~new_n48858_;
  assign new_n48860_ = ~new_n48109_ & ~new_n48815_;
  assign new_n48861_ = ~new_n48814_ & new_n48860_;
  assign new_n48862_ = ~new_n48859_ & ~new_n48861_;
  assign new_n48863_ = ~\b[50]  & ~new_n48862_;
  assign new_n48864_ = ~new_n48128_ & new_n48776_;
  assign new_n48865_ = ~new_n48772_ & new_n48864_;
  assign new_n48866_ = ~new_n48773_ & ~new_n48776_;
  assign new_n48867_ = ~new_n48865_ & ~new_n48866_;
  assign new_n48868_ = ~new_n48816_ & ~new_n48867_;
  assign new_n48869_ = ~new_n48118_ & ~new_n48815_;
  assign new_n48870_ = ~new_n48814_ & new_n48869_;
  assign new_n48871_ = ~new_n48868_ & ~new_n48870_;
  assign new_n48872_ = ~\b[49]  & ~new_n48871_;
  assign new_n48873_ = ~new_n48137_ & new_n48771_;
  assign new_n48874_ = ~new_n48767_ & new_n48873_;
  assign new_n48875_ = ~new_n48768_ & ~new_n48771_;
  assign new_n48876_ = ~new_n48874_ & ~new_n48875_;
  assign new_n48877_ = ~new_n48816_ & ~new_n48876_;
  assign new_n48878_ = ~new_n48127_ & ~new_n48815_;
  assign new_n48879_ = ~new_n48814_ & new_n48878_;
  assign new_n48880_ = ~new_n48877_ & ~new_n48879_;
  assign new_n48881_ = ~\b[48]  & ~new_n48880_;
  assign new_n48882_ = ~new_n48146_ & new_n48766_;
  assign new_n48883_ = ~new_n48762_ & new_n48882_;
  assign new_n48884_ = ~new_n48763_ & ~new_n48766_;
  assign new_n48885_ = ~new_n48883_ & ~new_n48884_;
  assign new_n48886_ = ~new_n48816_ & ~new_n48885_;
  assign new_n48887_ = ~new_n48136_ & ~new_n48815_;
  assign new_n48888_ = ~new_n48814_ & new_n48887_;
  assign new_n48889_ = ~new_n48886_ & ~new_n48888_;
  assign new_n48890_ = ~\b[47]  & ~new_n48889_;
  assign new_n48891_ = ~new_n48155_ & new_n48761_;
  assign new_n48892_ = ~new_n48757_ & new_n48891_;
  assign new_n48893_ = ~new_n48758_ & ~new_n48761_;
  assign new_n48894_ = ~new_n48892_ & ~new_n48893_;
  assign new_n48895_ = ~new_n48816_ & ~new_n48894_;
  assign new_n48896_ = ~new_n48145_ & ~new_n48815_;
  assign new_n48897_ = ~new_n48814_ & new_n48896_;
  assign new_n48898_ = ~new_n48895_ & ~new_n48897_;
  assign new_n48899_ = ~\b[46]  & ~new_n48898_;
  assign new_n48900_ = ~new_n48164_ & new_n48756_;
  assign new_n48901_ = ~new_n48752_ & new_n48900_;
  assign new_n48902_ = ~new_n48753_ & ~new_n48756_;
  assign new_n48903_ = ~new_n48901_ & ~new_n48902_;
  assign new_n48904_ = ~new_n48816_ & ~new_n48903_;
  assign new_n48905_ = ~new_n48154_ & ~new_n48815_;
  assign new_n48906_ = ~new_n48814_ & new_n48905_;
  assign new_n48907_ = ~new_n48904_ & ~new_n48906_;
  assign new_n48908_ = ~\b[45]  & ~new_n48907_;
  assign new_n48909_ = ~new_n48173_ & new_n48751_;
  assign new_n48910_ = ~new_n48747_ & new_n48909_;
  assign new_n48911_ = ~new_n48748_ & ~new_n48751_;
  assign new_n48912_ = ~new_n48910_ & ~new_n48911_;
  assign new_n48913_ = ~new_n48816_ & ~new_n48912_;
  assign new_n48914_ = ~new_n48163_ & ~new_n48815_;
  assign new_n48915_ = ~new_n48814_ & new_n48914_;
  assign new_n48916_ = ~new_n48913_ & ~new_n48915_;
  assign new_n48917_ = ~\b[44]  & ~new_n48916_;
  assign new_n48918_ = ~new_n48182_ & new_n48746_;
  assign new_n48919_ = ~new_n48742_ & new_n48918_;
  assign new_n48920_ = ~new_n48743_ & ~new_n48746_;
  assign new_n48921_ = ~new_n48919_ & ~new_n48920_;
  assign new_n48922_ = ~new_n48816_ & ~new_n48921_;
  assign new_n48923_ = ~new_n48172_ & ~new_n48815_;
  assign new_n48924_ = ~new_n48814_ & new_n48923_;
  assign new_n48925_ = ~new_n48922_ & ~new_n48924_;
  assign new_n48926_ = ~\b[43]  & ~new_n48925_;
  assign new_n48927_ = ~new_n48191_ & new_n48741_;
  assign new_n48928_ = ~new_n48737_ & new_n48927_;
  assign new_n48929_ = ~new_n48738_ & ~new_n48741_;
  assign new_n48930_ = ~new_n48928_ & ~new_n48929_;
  assign new_n48931_ = ~new_n48816_ & ~new_n48930_;
  assign new_n48932_ = ~new_n48181_ & ~new_n48815_;
  assign new_n48933_ = ~new_n48814_ & new_n48932_;
  assign new_n48934_ = ~new_n48931_ & ~new_n48933_;
  assign new_n48935_ = ~\b[42]  & ~new_n48934_;
  assign new_n48936_ = ~new_n48200_ & new_n48736_;
  assign new_n48937_ = ~new_n48732_ & new_n48936_;
  assign new_n48938_ = ~new_n48733_ & ~new_n48736_;
  assign new_n48939_ = ~new_n48937_ & ~new_n48938_;
  assign new_n48940_ = ~new_n48816_ & ~new_n48939_;
  assign new_n48941_ = ~new_n48190_ & ~new_n48815_;
  assign new_n48942_ = ~new_n48814_ & new_n48941_;
  assign new_n48943_ = ~new_n48940_ & ~new_n48942_;
  assign new_n48944_ = ~\b[41]  & ~new_n48943_;
  assign new_n48945_ = ~new_n48209_ & new_n48731_;
  assign new_n48946_ = ~new_n48727_ & new_n48945_;
  assign new_n48947_ = ~new_n48728_ & ~new_n48731_;
  assign new_n48948_ = ~new_n48946_ & ~new_n48947_;
  assign new_n48949_ = ~new_n48816_ & ~new_n48948_;
  assign new_n48950_ = ~new_n48199_ & ~new_n48815_;
  assign new_n48951_ = ~new_n48814_ & new_n48950_;
  assign new_n48952_ = ~new_n48949_ & ~new_n48951_;
  assign new_n48953_ = ~\b[40]  & ~new_n48952_;
  assign new_n48954_ = ~new_n48218_ & new_n48726_;
  assign new_n48955_ = ~new_n48722_ & new_n48954_;
  assign new_n48956_ = ~new_n48723_ & ~new_n48726_;
  assign new_n48957_ = ~new_n48955_ & ~new_n48956_;
  assign new_n48958_ = ~new_n48816_ & ~new_n48957_;
  assign new_n48959_ = ~new_n48208_ & ~new_n48815_;
  assign new_n48960_ = ~new_n48814_ & new_n48959_;
  assign new_n48961_ = ~new_n48958_ & ~new_n48960_;
  assign new_n48962_ = ~\b[39]  & ~new_n48961_;
  assign new_n48963_ = ~new_n48227_ & new_n48721_;
  assign new_n48964_ = ~new_n48717_ & new_n48963_;
  assign new_n48965_ = ~new_n48718_ & ~new_n48721_;
  assign new_n48966_ = ~new_n48964_ & ~new_n48965_;
  assign new_n48967_ = ~new_n48816_ & ~new_n48966_;
  assign new_n48968_ = ~new_n48217_ & ~new_n48815_;
  assign new_n48969_ = ~new_n48814_ & new_n48968_;
  assign new_n48970_ = ~new_n48967_ & ~new_n48969_;
  assign new_n48971_ = ~\b[38]  & ~new_n48970_;
  assign new_n48972_ = ~new_n48236_ & new_n48716_;
  assign new_n48973_ = ~new_n48712_ & new_n48972_;
  assign new_n48974_ = ~new_n48713_ & ~new_n48716_;
  assign new_n48975_ = ~new_n48973_ & ~new_n48974_;
  assign new_n48976_ = ~new_n48816_ & ~new_n48975_;
  assign new_n48977_ = ~new_n48226_ & ~new_n48815_;
  assign new_n48978_ = ~new_n48814_ & new_n48977_;
  assign new_n48979_ = ~new_n48976_ & ~new_n48978_;
  assign new_n48980_ = ~\b[37]  & ~new_n48979_;
  assign new_n48981_ = ~new_n48245_ & new_n48711_;
  assign new_n48982_ = ~new_n48707_ & new_n48981_;
  assign new_n48983_ = ~new_n48708_ & ~new_n48711_;
  assign new_n48984_ = ~new_n48982_ & ~new_n48983_;
  assign new_n48985_ = ~new_n48816_ & ~new_n48984_;
  assign new_n48986_ = ~new_n48235_ & ~new_n48815_;
  assign new_n48987_ = ~new_n48814_ & new_n48986_;
  assign new_n48988_ = ~new_n48985_ & ~new_n48987_;
  assign new_n48989_ = ~\b[36]  & ~new_n48988_;
  assign new_n48990_ = ~new_n48254_ & new_n48706_;
  assign new_n48991_ = ~new_n48702_ & new_n48990_;
  assign new_n48992_ = ~new_n48703_ & ~new_n48706_;
  assign new_n48993_ = ~new_n48991_ & ~new_n48992_;
  assign new_n48994_ = ~new_n48816_ & ~new_n48993_;
  assign new_n48995_ = ~new_n48244_ & ~new_n48815_;
  assign new_n48996_ = ~new_n48814_ & new_n48995_;
  assign new_n48997_ = ~new_n48994_ & ~new_n48996_;
  assign new_n48998_ = ~\b[35]  & ~new_n48997_;
  assign new_n48999_ = ~new_n48263_ & new_n48701_;
  assign new_n49000_ = ~new_n48697_ & new_n48999_;
  assign new_n49001_ = ~new_n48698_ & ~new_n48701_;
  assign new_n49002_ = ~new_n49000_ & ~new_n49001_;
  assign new_n49003_ = ~new_n48816_ & ~new_n49002_;
  assign new_n49004_ = ~new_n48253_ & ~new_n48815_;
  assign new_n49005_ = ~new_n48814_ & new_n49004_;
  assign new_n49006_ = ~new_n49003_ & ~new_n49005_;
  assign new_n49007_ = ~\b[34]  & ~new_n49006_;
  assign new_n49008_ = ~new_n48272_ & new_n48696_;
  assign new_n49009_ = ~new_n48692_ & new_n49008_;
  assign new_n49010_ = ~new_n48693_ & ~new_n48696_;
  assign new_n49011_ = ~new_n49009_ & ~new_n49010_;
  assign new_n49012_ = ~new_n48816_ & ~new_n49011_;
  assign new_n49013_ = ~new_n48262_ & ~new_n48815_;
  assign new_n49014_ = ~new_n48814_ & new_n49013_;
  assign new_n49015_ = ~new_n49012_ & ~new_n49014_;
  assign new_n49016_ = ~\b[33]  & ~new_n49015_;
  assign new_n49017_ = ~new_n48281_ & new_n48691_;
  assign new_n49018_ = ~new_n48687_ & new_n49017_;
  assign new_n49019_ = ~new_n48688_ & ~new_n48691_;
  assign new_n49020_ = ~new_n49018_ & ~new_n49019_;
  assign new_n49021_ = ~new_n48816_ & ~new_n49020_;
  assign new_n49022_ = ~new_n48271_ & ~new_n48815_;
  assign new_n49023_ = ~new_n48814_ & new_n49022_;
  assign new_n49024_ = ~new_n49021_ & ~new_n49023_;
  assign new_n49025_ = ~\b[32]  & ~new_n49024_;
  assign new_n49026_ = ~new_n48290_ & new_n48686_;
  assign new_n49027_ = ~new_n48682_ & new_n49026_;
  assign new_n49028_ = ~new_n48683_ & ~new_n48686_;
  assign new_n49029_ = ~new_n49027_ & ~new_n49028_;
  assign new_n49030_ = ~new_n48816_ & ~new_n49029_;
  assign new_n49031_ = ~new_n48280_ & ~new_n48815_;
  assign new_n49032_ = ~new_n48814_ & new_n49031_;
  assign new_n49033_ = ~new_n49030_ & ~new_n49032_;
  assign new_n49034_ = ~\b[31]  & ~new_n49033_;
  assign new_n49035_ = ~new_n48299_ & new_n48681_;
  assign new_n49036_ = ~new_n48677_ & new_n49035_;
  assign new_n49037_ = ~new_n48678_ & ~new_n48681_;
  assign new_n49038_ = ~new_n49036_ & ~new_n49037_;
  assign new_n49039_ = ~new_n48816_ & ~new_n49038_;
  assign new_n49040_ = ~new_n48289_ & ~new_n48815_;
  assign new_n49041_ = ~new_n48814_ & new_n49040_;
  assign new_n49042_ = ~new_n49039_ & ~new_n49041_;
  assign new_n49043_ = ~\b[30]  & ~new_n49042_;
  assign new_n49044_ = ~new_n48308_ & new_n48676_;
  assign new_n49045_ = ~new_n48672_ & new_n49044_;
  assign new_n49046_ = ~new_n48673_ & ~new_n48676_;
  assign new_n49047_ = ~new_n49045_ & ~new_n49046_;
  assign new_n49048_ = ~new_n48816_ & ~new_n49047_;
  assign new_n49049_ = ~new_n48298_ & ~new_n48815_;
  assign new_n49050_ = ~new_n48814_ & new_n49049_;
  assign new_n49051_ = ~new_n49048_ & ~new_n49050_;
  assign new_n49052_ = ~\b[29]  & ~new_n49051_;
  assign new_n49053_ = ~new_n48317_ & new_n48671_;
  assign new_n49054_ = ~new_n48667_ & new_n49053_;
  assign new_n49055_ = ~new_n48668_ & ~new_n48671_;
  assign new_n49056_ = ~new_n49054_ & ~new_n49055_;
  assign new_n49057_ = ~new_n48816_ & ~new_n49056_;
  assign new_n49058_ = ~new_n48307_ & ~new_n48815_;
  assign new_n49059_ = ~new_n48814_ & new_n49058_;
  assign new_n49060_ = ~new_n49057_ & ~new_n49059_;
  assign new_n49061_ = ~\b[28]  & ~new_n49060_;
  assign new_n49062_ = ~new_n48326_ & new_n48666_;
  assign new_n49063_ = ~new_n48662_ & new_n49062_;
  assign new_n49064_ = ~new_n48663_ & ~new_n48666_;
  assign new_n49065_ = ~new_n49063_ & ~new_n49064_;
  assign new_n49066_ = ~new_n48816_ & ~new_n49065_;
  assign new_n49067_ = ~new_n48316_ & ~new_n48815_;
  assign new_n49068_ = ~new_n48814_ & new_n49067_;
  assign new_n49069_ = ~new_n49066_ & ~new_n49068_;
  assign new_n49070_ = ~\b[27]  & ~new_n49069_;
  assign new_n49071_ = ~new_n48335_ & new_n48661_;
  assign new_n49072_ = ~new_n48657_ & new_n49071_;
  assign new_n49073_ = ~new_n48658_ & ~new_n48661_;
  assign new_n49074_ = ~new_n49072_ & ~new_n49073_;
  assign new_n49075_ = ~new_n48816_ & ~new_n49074_;
  assign new_n49076_ = ~new_n48325_ & ~new_n48815_;
  assign new_n49077_ = ~new_n48814_ & new_n49076_;
  assign new_n49078_ = ~new_n49075_ & ~new_n49077_;
  assign new_n49079_ = ~\b[26]  & ~new_n49078_;
  assign new_n49080_ = ~new_n48344_ & new_n48656_;
  assign new_n49081_ = ~new_n48652_ & new_n49080_;
  assign new_n49082_ = ~new_n48653_ & ~new_n48656_;
  assign new_n49083_ = ~new_n49081_ & ~new_n49082_;
  assign new_n49084_ = ~new_n48816_ & ~new_n49083_;
  assign new_n49085_ = ~new_n48334_ & ~new_n48815_;
  assign new_n49086_ = ~new_n48814_ & new_n49085_;
  assign new_n49087_ = ~new_n49084_ & ~new_n49086_;
  assign new_n49088_ = ~\b[25]  & ~new_n49087_;
  assign new_n49089_ = ~new_n48353_ & new_n48651_;
  assign new_n49090_ = ~new_n48647_ & new_n49089_;
  assign new_n49091_ = ~new_n48648_ & ~new_n48651_;
  assign new_n49092_ = ~new_n49090_ & ~new_n49091_;
  assign new_n49093_ = ~new_n48816_ & ~new_n49092_;
  assign new_n49094_ = ~new_n48343_ & ~new_n48815_;
  assign new_n49095_ = ~new_n48814_ & new_n49094_;
  assign new_n49096_ = ~new_n49093_ & ~new_n49095_;
  assign new_n49097_ = ~\b[24]  & ~new_n49096_;
  assign new_n49098_ = ~new_n48362_ & new_n48646_;
  assign new_n49099_ = ~new_n48642_ & new_n49098_;
  assign new_n49100_ = ~new_n48643_ & ~new_n48646_;
  assign new_n49101_ = ~new_n49099_ & ~new_n49100_;
  assign new_n49102_ = ~new_n48816_ & ~new_n49101_;
  assign new_n49103_ = ~new_n48352_ & ~new_n48815_;
  assign new_n49104_ = ~new_n48814_ & new_n49103_;
  assign new_n49105_ = ~new_n49102_ & ~new_n49104_;
  assign new_n49106_ = ~\b[23]  & ~new_n49105_;
  assign new_n49107_ = ~new_n48371_ & new_n48641_;
  assign new_n49108_ = ~new_n48637_ & new_n49107_;
  assign new_n49109_ = ~new_n48638_ & ~new_n48641_;
  assign new_n49110_ = ~new_n49108_ & ~new_n49109_;
  assign new_n49111_ = ~new_n48816_ & ~new_n49110_;
  assign new_n49112_ = ~new_n48361_ & ~new_n48815_;
  assign new_n49113_ = ~new_n48814_ & new_n49112_;
  assign new_n49114_ = ~new_n49111_ & ~new_n49113_;
  assign new_n49115_ = ~\b[22]  & ~new_n49114_;
  assign new_n49116_ = ~new_n48380_ & new_n48636_;
  assign new_n49117_ = ~new_n48632_ & new_n49116_;
  assign new_n49118_ = ~new_n48633_ & ~new_n48636_;
  assign new_n49119_ = ~new_n49117_ & ~new_n49118_;
  assign new_n49120_ = ~new_n48816_ & ~new_n49119_;
  assign new_n49121_ = ~new_n48370_ & ~new_n48815_;
  assign new_n49122_ = ~new_n48814_ & new_n49121_;
  assign new_n49123_ = ~new_n49120_ & ~new_n49122_;
  assign new_n49124_ = ~\b[21]  & ~new_n49123_;
  assign new_n49125_ = ~new_n48389_ & new_n48631_;
  assign new_n49126_ = ~new_n48627_ & new_n49125_;
  assign new_n49127_ = ~new_n48628_ & ~new_n48631_;
  assign new_n49128_ = ~new_n49126_ & ~new_n49127_;
  assign new_n49129_ = ~new_n48816_ & ~new_n49128_;
  assign new_n49130_ = ~new_n48379_ & ~new_n48815_;
  assign new_n49131_ = ~new_n48814_ & new_n49130_;
  assign new_n49132_ = ~new_n49129_ & ~new_n49131_;
  assign new_n49133_ = ~\b[20]  & ~new_n49132_;
  assign new_n49134_ = ~new_n48398_ & new_n48626_;
  assign new_n49135_ = ~new_n48622_ & new_n49134_;
  assign new_n49136_ = ~new_n48623_ & ~new_n48626_;
  assign new_n49137_ = ~new_n49135_ & ~new_n49136_;
  assign new_n49138_ = ~new_n48816_ & ~new_n49137_;
  assign new_n49139_ = ~new_n48388_ & ~new_n48815_;
  assign new_n49140_ = ~new_n48814_ & new_n49139_;
  assign new_n49141_ = ~new_n49138_ & ~new_n49140_;
  assign new_n49142_ = ~\b[19]  & ~new_n49141_;
  assign new_n49143_ = ~new_n48407_ & new_n48621_;
  assign new_n49144_ = ~new_n48617_ & new_n49143_;
  assign new_n49145_ = ~new_n48618_ & ~new_n48621_;
  assign new_n49146_ = ~new_n49144_ & ~new_n49145_;
  assign new_n49147_ = ~new_n48816_ & ~new_n49146_;
  assign new_n49148_ = ~new_n48397_ & ~new_n48815_;
  assign new_n49149_ = ~new_n48814_ & new_n49148_;
  assign new_n49150_ = ~new_n49147_ & ~new_n49149_;
  assign new_n49151_ = ~\b[18]  & ~new_n49150_;
  assign new_n49152_ = ~new_n48416_ & new_n48616_;
  assign new_n49153_ = ~new_n48612_ & new_n49152_;
  assign new_n49154_ = ~new_n48613_ & ~new_n48616_;
  assign new_n49155_ = ~new_n49153_ & ~new_n49154_;
  assign new_n49156_ = ~new_n48816_ & ~new_n49155_;
  assign new_n49157_ = ~new_n48406_ & ~new_n48815_;
  assign new_n49158_ = ~new_n48814_ & new_n49157_;
  assign new_n49159_ = ~new_n49156_ & ~new_n49158_;
  assign new_n49160_ = ~\b[17]  & ~new_n49159_;
  assign new_n49161_ = ~new_n48425_ & new_n48611_;
  assign new_n49162_ = ~new_n48607_ & new_n49161_;
  assign new_n49163_ = ~new_n48608_ & ~new_n48611_;
  assign new_n49164_ = ~new_n49162_ & ~new_n49163_;
  assign new_n49165_ = ~new_n48816_ & ~new_n49164_;
  assign new_n49166_ = ~new_n48415_ & ~new_n48815_;
  assign new_n49167_ = ~new_n48814_ & new_n49166_;
  assign new_n49168_ = ~new_n49165_ & ~new_n49167_;
  assign new_n49169_ = ~\b[16]  & ~new_n49168_;
  assign new_n49170_ = ~new_n48434_ & new_n48606_;
  assign new_n49171_ = ~new_n48602_ & new_n49170_;
  assign new_n49172_ = ~new_n48603_ & ~new_n48606_;
  assign new_n49173_ = ~new_n49171_ & ~new_n49172_;
  assign new_n49174_ = ~new_n48816_ & ~new_n49173_;
  assign new_n49175_ = ~new_n48424_ & ~new_n48815_;
  assign new_n49176_ = ~new_n48814_ & new_n49175_;
  assign new_n49177_ = ~new_n49174_ & ~new_n49176_;
  assign new_n49178_ = ~\b[15]  & ~new_n49177_;
  assign new_n49179_ = ~new_n48443_ & new_n48601_;
  assign new_n49180_ = ~new_n48597_ & new_n49179_;
  assign new_n49181_ = ~new_n48598_ & ~new_n48601_;
  assign new_n49182_ = ~new_n49180_ & ~new_n49181_;
  assign new_n49183_ = ~new_n48816_ & ~new_n49182_;
  assign new_n49184_ = ~new_n48433_ & ~new_n48815_;
  assign new_n49185_ = ~new_n48814_ & new_n49184_;
  assign new_n49186_ = ~new_n49183_ & ~new_n49185_;
  assign new_n49187_ = ~\b[14]  & ~new_n49186_;
  assign new_n49188_ = ~new_n48452_ & new_n48596_;
  assign new_n49189_ = ~new_n48592_ & new_n49188_;
  assign new_n49190_ = ~new_n48593_ & ~new_n48596_;
  assign new_n49191_ = ~new_n49189_ & ~new_n49190_;
  assign new_n49192_ = ~new_n48816_ & ~new_n49191_;
  assign new_n49193_ = ~new_n48442_ & ~new_n48815_;
  assign new_n49194_ = ~new_n48814_ & new_n49193_;
  assign new_n49195_ = ~new_n49192_ & ~new_n49194_;
  assign new_n49196_ = ~\b[13]  & ~new_n49195_;
  assign new_n49197_ = ~new_n48461_ & new_n48591_;
  assign new_n49198_ = ~new_n48587_ & new_n49197_;
  assign new_n49199_ = ~new_n48588_ & ~new_n48591_;
  assign new_n49200_ = ~new_n49198_ & ~new_n49199_;
  assign new_n49201_ = ~new_n48816_ & ~new_n49200_;
  assign new_n49202_ = ~new_n48451_ & ~new_n48815_;
  assign new_n49203_ = ~new_n48814_ & new_n49202_;
  assign new_n49204_ = ~new_n49201_ & ~new_n49203_;
  assign new_n49205_ = ~\b[12]  & ~new_n49204_;
  assign new_n49206_ = ~new_n48470_ & new_n48586_;
  assign new_n49207_ = ~new_n48582_ & new_n49206_;
  assign new_n49208_ = ~new_n48583_ & ~new_n48586_;
  assign new_n49209_ = ~new_n49207_ & ~new_n49208_;
  assign new_n49210_ = ~new_n48816_ & ~new_n49209_;
  assign new_n49211_ = ~new_n48460_ & ~new_n48815_;
  assign new_n49212_ = ~new_n48814_ & new_n49211_;
  assign new_n49213_ = ~new_n49210_ & ~new_n49212_;
  assign new_n49214_ = ~\b[11]  & ~new_n49213_;
  assign new_n49215_ = ~new_n48479_ & new_n48581_;
  assign new_n49216_ = ~new_n48577_ & new_n49215_;
  assign new_n49217_ = ~new_n48578_ & ~new_n48581_;
  assign new_n49218_ = ~new_n49216_ & ~new_n49217_;
  assign new_n49219_ = ~new_n48816_ & ~new_n49218_;
  assign new_n49220_ = ~new_n48469_ & ~new_n48815_;
  assign new_n49221_ = ~new_n48814_ & new_n49220_;
  assign new_n49222_ = ~new_n49219_ & ~new_n49221_;
  assign new_n49223_ = ~\b[10]  & ~new_n49222_;
  assign new_n49224_ = ~new_n48488_ & new_n48576_;
  assign new_n49225_ = ~new_n48572_ & new_n49224_;
  assign new_n49226_ = ~new_n48573_ & ~new_n48576_;
  assign new_n49227_ = ~new_n49225_ & ~new_n49226_;
  assign new_n49228_ = ~new_n48816_ & ~new_n49227_;
  assign new_n49229_ = ~new_n48478_ & ~new_n48815_;
  assign new_n49230_ = ~new_n48814_ & new_n49229_;
  assign new_n49231_ = ~new_n49228_ & ~new_n49230_;
  assign new_n49232_ = ~\b[9]  & ~new_n49231_;
  assign new_n49233_ = ~new_n48497_ & new_n48571_;
  assign new_n49234_ = ~new_n48567_ & new_n49233_;
  assign new_n49235_ = ~new_n48568_ & ~new_n48571_;
  assign new_n49236_ = ~new_n49234_ & ~new_n49235_;
  assign new_n49237_ = ~new_n48816_ & ~new_n49236_;
  assign new_n49238_ = ~new_n48487_ & ~new_n48815_;
  assign new_n49239_ = ~new_n48814_ & new_n49238_;
  assign new_n49240_ = ~new_n49237_ & ~new_n49239_;
  assign new_n49241_ = ~\b[8]  & ~new_n49240_;
  assign new_n49242_ = ~new_n48506_ & new_n48566_;
  assign new_n49243_ = ~new_n48562_ & new_n49242_;
  assign new_n49244_ = ~new_n48563_ & ~new_n48566_;
  assign new_n49245_ = ~new_n49243_ & ~new_n49244_;
  assign new_n49246_ = ~new_n48816_ & ~new_n49245_;
  assign new_n49247_ = ~new_n48496_ & ~new_n48815_;
  assign new_n49248_ = ~new_n48814_ & new_n49247_;
  assign new_n49249_ = ~new_n49246_ & ~new_n49248_;
  assign new_n49250_ = ~\b[7]  & ~new_n49249_;
  assign new_n49251_ = ~new_n48515_ & new_n48561_;
  assign new_n49252_ = ~new_n48557_ & new_n49251_;
  assign new_n49253_ = ~new_n48558_ & ~new_n48561_;
  assign new_n49254_ = ~new_n49252_ & ~new_n49253_;
  assign new_n49255_ = ~new_n48816_ & ~new_n49254_;
  assign new_n49256_ = ~new_n48505_ & ~new_n48815_;
  assign new_n49257_ = ~new_n48814_ & new_n49256_;
  assign new_n49258_ = ~new_n49255_ & ~new_n49257_;
  assign new_n49259_ = ~\b[6]  & ~new_n49258_;
  assign new_n49260_ = ~new_n48524_ & new_n48556_;
  assign new_n49261_ = ~new_n48552_ & new_n49260_;
  assign new_n49262_ = ~new_n48553_ & ~new_n48556_;
  assign new_n49263_ = ~new_n49261_ & ~new_n49262_;
  assign new_n49264_ = ~new_n48816_ & ~new_n49263_;
  assign new_n49265_ = ~new_n48514_ & ~new_n48815_;
  assign new_n49266_ = ~new_n48814_ & new_n49265_;
  assign new_n49267_ = ~new_n49264_ & ~new_n49266_;
  assign new_n49268_ = ~\b[5]  & ~new_n49267_;
  assign new_n49269_ = ~new_n48532_ & new_n48551_;
  assign new_n49270_ = ~new_n48547_ & new_n49269_;
  assign new_n49271_ = ~new_n48548_ & ~new_n48551_;
  assign new_n49272_ = ~new_n49270_ & ~new_n49271_;
  assign new_n49273_ = ~new_n48816_ & ~new_n49272_;
  assign new_n49274_ = ~new_n48523_ & ~new_n48815_;
  assign new_n49275_ = ~new_n48814_ & new_n49274_;
  assign new_n49276_ = ~new_n49273_ & ~new_n49275_;
  assign new_n49277_ = ~\b[4]  & ~new_n49276_;
  assign new_n49278_ = ~new_n48542_ & new_n48546_;
  assign new_n49279_ = ~new_n48541_ & new_n49278_;
  assign new_n49280_ = ~new_n48543_ & ~new_n48546_;
  assign new_n49281_ = ~new_n49279_ & ~new_n49280_;
  assign new_n49282_ = ~new_n48816_ & ~new_n49281_;
  assign new_n49283_ = ~new_n48531_ & ~new_n48815_;
  assign new_n49284_ = ~new_n48814_ & new_n49283_;
  assign new_n49285_ = ~new_n49282_ & ~new_n49284_;
  assign new_n49286_ = ~\b[3]  & ~new_n49285_;
  assign new_n49287_ = new_n20502_ & ~new_n48539_;
  assign new_n49288_ = ~new_n48537_ & new_n49287_;
  assign new_n49289_ = ~new_n48541_ & ~new_n49288_;
  assign new_n49290_ = ~new_n48816_ & new_n49289_;
  assign new_n49291_ = ~new_n48536_ & ~new_n48815_;
  assign new_n49292_ = ~new_n48814_ & new_n49291_;
  assign new_n49293_ = ~new_n49290_ & ~new_n49292_;
  assign new_n49294_ = ~\b[2]  & ~new_n49293_;
  assign new_n49295_ = \b[0]  & ~new_n48816_;
  assign new_n49296_ = \a[10]  & ~new_n49295_;
  assign new_n49297_ = new_n20502_ & ~new_n48816_;
  assign new_n49298_ = ~new_n49296_ & ~new_n49297_;
  assign new_n49299_ = \b[1]  & ~new_n49298_;
  assign new_n49300_ = ~\b[1]  & ~new_n49297_;
  assign new_n49301_ = ~new_n49296_ & new_n49300_;
  assign new_n49302_ = ~new_n49299_ & ~new_n49301_;
  assign new_n49303_ = ~new_n21267_ & ~new_n49302_;
  assign new_n49304_ = ~\b[1]  & ~new_n49298_;
  assign new_n49305_ = ~new_n49303_ & ~new_n49304_;
  assign new_n49306_ = \b[2]  & ~new_n49292_;
  assign new_n49307_ = ~new_n49290_ & new_n49306_;
  assign new_n49308_ = ~new_n49294_ & ~new_n49307_;
  assign new_n49309_ = ~new_n49305_ & new_n49308_;
  assign new_n49310_ = ~new_n49294_ & ~new_n49309_;
  assign new_n49311_ = \b[3]  & ~new_n49284_;
  assign new_n49312_ = ~new_n49282_ & new_n49311_;
  assign new_n49313_ = ~new_n49286_ & ~new_n49312_;
  assign new_n49314_ = ~new_n49310_ & new_n49313_;
  assign new_n49315_ = ~new_n49286_ & ~new_n49314_;
  assign new_n49316_ = \b[4]  & ~new_n49275_;
  assign new_n49317_ = ~new_n49273_ & new_n49316_;
  assign new_n49318_ = ~new_n49277_ & ~new_n49317_;
  assign new_n49319_ = ~new_n49315_ & new_n49318_;
  assign new_n49320_ = ~new_n49277_ & ~new_n49319_;
  assign new_n49321_ = \b[5]  & ~new_n49266_;
  assign new_n49322_ = ~new_n49264_ & new_n49321_;
  assign new_n49323_ = ~new_n49268_ & ~new_n49322_;
  assign new_n49324_ = ~new_n49320_ & new_n49323_;
  assign new_n49325_ = ~new_n49268_ & ~new_n49324_;
  assign new_n49326_ = \b[6]  & ~new_n49257_;
  assign new_n49327_ = ~new_n49255_ & new_n49326_;
  assign new_n49328_ = ~new_n49259_ & ~new_n49327_;
  assign new_n49329_ = ~new_n49325_ & new_n49328_;
  assign new_n49330_ = ~new_n49259_ & ~new_n49329_;
  assign new_n49331_ = \b[7]  & ~new_n49248_;
  assign new_n49332_ = ~new_n49246_ & new_n49331_;
  assign new_n49333_ = ~new_n49250_ & ~new_n49332_;
  assign new_n49334_ = ~new_n49330_ & new_n49333_;
  assign new_n49335_ = ~new_n49250_ & ~new_n49334_;
  assign new_n49336_ = \b[8]  & ~new_n49239_;
  assign new_n49337_ = ~new_n49237_ & new_n49336_;
  assign new_n49338_ = ~new_n49241_ & ~new_n49337_;
  assign new_n49339_ = ~new_n49335_ & new_n49338_;
  assign new_n49340_ = ~new_n49241_ & ~new_n49339_;
  assign new_n49341_ = \b[9]  & ~new_n49230_;
  assign new_n49342_ = ~new_n49228_ & new_n49341_;
  assign new_n49343_ = ~new_n49232_ & ~new_n49342_;
  assign new_n49344_ = ~new_n49340_ & new_n49343_;
  assign new_n49345_ = ~new_n49232_ & ~new_n49344_;
  assign new_n49346_ = \b[10]  & ~new_n49221_;
  assign new_n49347_ = ~new_n49219_ & new_n49346_;
  assign new_n49348_ = ~new_n49223_ & ~new_n49347_;
  assign new_n49349_ = ~new_n49345_ & new_n49348_;
  assign new_n49350_ = ~new_n49223_ & ~new_n49349_;
  assign new_n49351_ = \b[11]  & ~new_n49212_;
  assign new_n49352_ = ~new_n49210_ & new_n49351_;
  assign new_n49353_ = ~new_n49214_ & ~new_n49352_;
  assign new_n49354_ = ~new_n49350_ & new_n49353_;
  assign new_n49355_ = ~new_n49214_ & ~new_n49354_;
  assign new_n49356_ = \b[12]  & ~new_n49203_;
  assign new_n49357_ = ~new_n49201_ & new_n49356_;
  assign new_n49358_ = ~new_n49205_ & ~new_n49357_;
  assign new_n49359_ = ~new_n49355_ & new_n49358_;
  assign new_n49360_ = ~new_n49205_ & ~new_n49359_;
  assign new_n49361_ = \b[13]  & ~new_n49194_;
  assign new_n49362_ = ~new_n49192_ & new_n49361_;
  assign new_n49363_ = ~new_n49196_ & ~new_n49362_;
  assign new_n49364_ = ~new_n49360_ & new_n49363_;
  assign new_n49365_ = ~new_n49196_ & ~new_n49364_;
  assign new_n49366_ = \b[14]  & ~new_n49185_;
  assign new_n49367_ = ~new_n49183_ & new_n49366_;
  assign new_n49368_ = ~new_n49187_ & ~new_n49367_;
  assign new_n49369_ = ~new_n49365_ & new_n49368_;
  assign new_n49370_ = ~new_n49187_ & ~new_n49369_;
  assign new_n49371_ = \b[15]  & ~new_n49176_;
  assign new_n49372_ = ~new_n49174_ & new_n49371_;
  assign new_n49373_ = ~new_n49178_ & ~new_n49372_;
  assign new_n49374_ = ~new_n49370_ & new_n49373_;
  assign new_n49375_ = ~new_n49178_ & ~new_n49374_;
  assign new_n49376_ = \b[16]  & ~new_n49167_;
  assign new_n49377_ = ~new_n49165_ & new_n49376_;
  assign new_n49378_ = ~new_n49169_ & ~new_n49377_;
  assign new_n49379_ = ~new_n49375_ & new_n49378_;
  assign new_n49380_ = ~new_n49169_ & ~new_n49379_;
  assign new_n49381_ = \b[17]  & ~new_n49158_;
  assign new_n49382_ = ~new_n49156_ & new_n49381_;
  assign new_n49383_ = ~new_n49160_ & ~new_n49382_;
  assign new_n49384_ = ~new_n49380_ & new_n49383_;
  assign new_n49385_ = ~new_n49160_ & ~new_n49384_;
  assign new_n49386_ = \b[18]  & ~new_n49149_;
  assign new_n49387_ = ~new_n49147_ & new_n49386_;
  assign new_n49388_ = ~new_n49151_ & ~new_n49387_;
  assign new_n49389_ = ~new_n49385_ & new_n49388_;
  assign new_n49390_ = ~new_n49151_ & ~new_n49389_;
  assign new_n49391_ = \b[19]  & ~new_n49140_;
  assign new_n49392_ = ~new_n49138_ & new_n49391_;
  assign new_n49393_ = ~new_n49142_ & ~new_n49392_;
  assign new_n49394_ = ~new_n49390_ & new_n49393_;
  assign new_n49395_ = ~new_n49142_ & ~new_n49394_;
  assign new_n49396_ = \b[20]  & ~new_n49131_;
  assign new_n49397_ = ~new_n49129_ & new_n49396_;
  assign new_n49398_ = ~new_n49133_ & ~new_n49397_;
  assign new_n49399_ = ~new_n49395_ & new_n49398_;
  assign new_n49400_ = ~new_n49133_ & ~new_n49399_;
  assign new_n49401_ = \b[21]  & ~new_n49122_;
  assign new_n49402_ = ~new_n49120_ & new_n49401_;
  assign new_n49403_ = ~new_n49124_ & ~new_n49402_;
  assign new_n49404_ = ~new_n49400_ & new_n49403_;
  assign new_n49405_ = ~new_n49124_ & ~new_n49404_;
  assign new_n49406_ = \b[22]  & ~new_n49113_;
  assign new_n49407_ = ~new_n49111_ & new_n49406_;
  assign new_n49408_ = ~new_n49115_ & ~new_n49407_;
  assign new_n49409_ = ~new_n49405_ & new_n49408_;
  assign new_n49410_ = ~new_n49115_ & ~new_n49409_;
  assign new_n49411_ = \b[23]  & ~new_n49104_;
  assign new_n49412_ = ~new_n49102_ & new_n49411_;
  assign new_n49413_ = ~new_n49106_ & ~new_n49412_;
  assign new_n49414_ = ~new_n49410_ & new_n49413_;
  assign new_n49415_ = ~new_n49106_ & ~new_n49414_;
  assign new_n49416_ = \b[24]  & ~new_n49095_;
  assign new_n49417_ = ~new_n49093_ & new_n49416_;
  assign new_n49418_ = ~new_n49097_ & ~new_n49417_;
  assign new_n49419_ = ~new_n49415_ & new_n49418_;
  assign new_n49420_ = ~new_n49097_ & ~new_n49419_;
  assign new_n49421_ = \b[25]  & ~new_n49086_;
  assign new_n49422_ = ~new_n49084_ & new_n49421_;
  assign new_n49423_ = ~new_n49088_ & ~new_n49422_;
  assign new_n49424_ = ~new_n49420_ & new_n49423_;
  assign new_n49425_ = ~new_n49088_ & ~new_n49424_;
  assign new_n49426_ = \b[26]  & ~new_n49077_;
  assign new_n49427_ = ~new_n49075_ & new_n49426_;
  assign new_n49428_ = ~new_n49079_ & ~new_n49427_;
  assign new_n49429_ = ~new_n49425_ & new_n49428_;
  assign new_n49430_ = ~new_n49079_ & ~new_n49429_;
  assign new_n49431_ = \b[27]  & ~new_n49068_;
  assign new_n49432_ = ~new_n49066_ & new_n49431_;
  assign new_n49433_ = ~new_n49070_ & ~new_n49432_;
  assign new_n49434_ = ~new_n49430_ & new_n49433_;
  assign new_n49435_ = ~new_n49070_ & ~new_n49434_;
  assign new_n49436_ = \b[28]  & ~new_n49059_;
  assign new_n49437_ = ~new_n49057_ & new_n49436_;
  assign new_n49438_ = ~new_n49061_ & ~new_n49437_;
  assign new_n49439_ = ~new_n49435_ & new_n49438_;
  assign new_n49440_ = ~new_n49061_ & ~new_n49439_;
  assign new_n49441_ = \b[29]  & ~new_n49050_;
  assign new_n49442_ = ~new_n49048_ & new_n49441_;
  assign new_n49443_ = ~new_n49052_ & ~new_n49442_;
  assign new_n49444_ = ~new_n49440_ & new_n49443_;
  assign new_n49445_ = ~new_n49052_ & ~new_n49444_;
  assign new_n49446_ = \b[30]  & ~new_n49041_;
  assign new_n49447_ = ~new_n49039_ & new_n49446_;
  assign new_n49448_ = ~new_n49043_ & ~new_n49447_;
  assign new_n49449_ = ~new_n49445_ & new_n49448_;
  assign new_n49450_ = ~new_n49043_ & ~new_n49449_;
  assign new_n49451_ = \b[31]  & ~new_n49032_;
  assign new_n49452_ = ~new_n49030_ & new_n49451_;
  assign new_n49453_ = ~new_n49034_ & ~new_n49452_;
  assign new_n49454_ = ~new_n49450_ & new_n49453_;
  assign new_n49455_ = ~new_n49034_ & ~new_n49454_;
  assign new_n49456_ = \b[32]  & ~new_n49023_;
  assign new_n49457_ = ~new_n49021_ & new_n49456_;
  assign new_n49458_ = ~new_n49025_ & ~new_n49457_;
  assign new_n49459_ = ~new_n49455_ & new_n49458_;
  assign new_n49460_ = ~new_n49025_ & ~new_n49459_;
  assign new_n49461_ = \b[33]  & ~new_n49014_;
  assign new_n49462_ = ~new_n49012_ & new_n49461_;
  assign new_n49463_ = ~new_n49016_ & ~new_n49462_;
  assign new_n49464_ = ~new_n49460_ & new_n49463_;
  assign new_n49465_ = ~new_n49016_ & ~new_n49464_;
  assign new_n49466_ = \b[34]  & ~new_n49005_;
  assign new_n49467_ = ~new_n49003_ & new_n49466_;
  assign new_n49468_ = ~new_n49007_ & ~new_n49467_;
  assign new_n49469_ = ~new_n49465_ & new_n49468_;
  assign new_n49470_ = ~new_n49007_ & ~new_n49469_;
  assign new_n49471_ = \b[35]  & ~new_n48996_;
  assign new_n49472_ = ~new_n48994_ & new_n49471_;
  assign new_n49473_ = ~new_n48998_ & ~new_n49472_;
  assign new_n49474_ = ~new_n49470_ & new_n49473_;
  assign new_n49475_ = ~new_n48998_ & ~new_n49474_;
  assign new_n49476_ = \b[36]  & ~new_n48987_;
  assign new_n49477_ = ~new_n48985_ & new_n49476_;
  assign new_n49478_ = ~new_n48989_ & ~new_n49477_;
  assign new_n49479_ = ~new_n49475_ & new_n49478_;
  assign new_n49480_ = ~new_n48989_ & ~new_n49479_;
  assign new_n49481_ = \b[37]  & ~new_n48978_;
  assign new_n49482_ = ~new_n48976_ & new_n49481_;
  assign new_n49483_ = ~new_n48980_ & ~new_n49482_;
  assign new_n49484_ = ~new_n49480_ & new_n49483_;
  assign new_n49485_ = ~new_n48980_ & ~new_n49484_;
  assign new_n49486_ = \b[38]  & ~new_n48969_;
  assign new_n49487_ = ~new_n48967_ & new_n49486_;
  assign new_n49488_ = ~new_n48971_ & ~new_n49487_;
  assign new_n49489_ = ~new_n49485_ & new_n49488_;
  assign new_n49490_ = ~new_n48971_ & ~new_n49489_;
  assign new_n49491_ = \b[39]  & ~new_n48960_;
  assign new_n49492_ = ~new_n48958_ & new_n49491_;
  assign new_n49493_ = ~new_n48962_ & ~new_n49492_;
  assign new_n49494_ = ~new_n49490_ & new_n49493_;
  assign new_n49495_ = ~new_n48962_ & ~new_n49494_;
  assign new_n49496_ = \b[40]  & ~new_n48951_;
  assign new_n49497_ = ~new_n48949_ & new_n49496_;
  assign new_n49498_ = ~new_n48953_ & ~new_n49497_;
  assign new_n49499_ = ~new_n49495_ & new_n49498_;
  assign new_n49500_ = ~new_n48953_ & ~new_n49499_;
  assign new_n49501_ = \b[41]  & ~new_n48942_;
  assign new_n49502_ = ~new_n48940_ & new_n49501_;
  assign new_n49503_ = ~new_n48944_ & ~new_n49502_;
  assign new_n49504_ = ~new_n49500_ & new_n49503_;
  assign new_n49505_ = ~new_n48944_ & ~new_n49504_;
  assign new_n49506_ = \b[42]  & ~new_n48933_;
  assign new_n49507_ = ~new_n48931_ & new_n49506_;
  assign new_n49508_ = ~new_n48935_ & ~new_n49507_;
  assign new_n49509_ = ~new_n49505_ & new_n49508_;
  assign new_n49510_ = ~new_n48935_ & ~new_n49509_;
  assign new_n49511_ = \b[43]  & ~new_n48924_;
  assign new_n49512_ = ~new_n48922_ & new_n49511_;
  assign new_n49513_ = ~new_n48926_ & ~new_n49512_;
  assign new_n49514_ = ~new_n49510_ & new_n49513_;
  assign new_n49515_ = ~new_n48926_ & ~new_n49514_;
  assign new_n49516_ = \b[44]  & ~new_n48915_;
  assign new_n49517_ = ~new_n48913_ & new_n49516_;
  assign new_n49518_ = ~new_n48917_ & ~new_n49517_;
  assign new_n49519_ = ~new_n49515_ & new_n49518_;
  assign new_n49520_ = ~new_n48917_ & ~new_n49519_;
  assign new_n49521_ = \b[45]  & ~new_n48906_;
  assign new_n49522_ = ~new_n48904_ & new_n49521_;
  assign new_n49523_ = ~new_n48908_ & ~new_n49522_;
  assign new_n49524_ = ~new_n49520_ & new_n49523_;
  assign new_n49525_ = ~new_n48908_ & ~new_n49524_;
  assign new_n49526_ = \b[46]  & ~new_n48897_;
  assign new_n49527_ = ~new_n48895_ & new_n49526_;
  assign new_n49528_ = ~new_n48899_ & ~new_n49527_;
  assign new_n49529_ = ~new_n49525_ & new_n49528_;
  assign new_n49530_ = ~new_n48899_ & ~new_n49529_;
  assign new_n49531_ = \b[47]  & ~new_n48888_;
  assign new_n49532_ = ~new_n48886_ & new_n49531_;
  assign new_n49533_ = ~new_n48890_ & ~new_n49532_;
  assign new_n49534_ = ~new_n49530_ & new_n49533_;
  assign new_n49535_ = ~new_n48890_ & ~new_n49534_;
  assign new_n49536_ = \b[48]  & ~new_n48879_;
  assign new_n49537_ = ~new_n48877_ & new_n49536_;
  assign new_n49538_ = ~new_n48881_ & ~new_n49537_;
  assign new_n49539_ = ~new_n49535_ & new_n49538_;
  assign new_n49540_ = ~new_n48881_ & ~new_n49539_;
  assign new_n49541_ = \b[49]  & ~new_n48870_;
  assign new_n49542_ = ~new_n48868_ & new_n49541_;
  assign new_n49543_ = ~new_n48872_ & ~new_n49542_;
  assign new_n49544_ = ~new_n49540_ & new_n49543_;
  assign new_n49545_ = ~new_n48872_ & ~new_n49544_;
  assign new_n49546_ = \b[50]  & ~new_n48861_;
  assign new_n49547_ = ~new_n48859_ & new_n49546_;
  assign new_n49548_ = ~new_n48863_ & ~new_n49547_;
  assign new_n49549_ = ~new_n49545_ & new_n49548_;
  assign new_n49550_ = ~new_n48863_ & ~new_n49549_;
  assign new_n49551_ = \b[51]  & ~new_n48852_;
  assign new_n49552_ = ~new_n48850_ & new_n49551_;
  assign new_n49553_ = ~new_n48854_ & ~new_n49552_;
  assign new_n49554_ = ~new_n49550_ & new_n49553_;
  assign new_n49555_ = ~new_n48854_ & ~new_n49554_;
  assign new_n49556_ = \b[52]  & ~new_n48843_;
  assign new_n49557_ = ~new_n48841_ & new_n49556_;
  assign new_n49558_ = ~new_n48845_ & ~new_n49557_;
  assign new_n49559_ = ~new_n49555_ & new_n49558_;
  assign new_n49560_ = ~new_n48845_ & ~new_n49559_;
  assign new_n49561_ = \b[53]  & ~new_n48823_;
  assign new_n49562_ = ~new_n48821_ & new_n49561_;
  assign new_n49563_ = ~new_n48836_ & ~new_n49562_;
  assign new_n49564_ = ~new_n49560_ & new_n49563_;
  assign new_n49565_ = ~new_n48836_ & ~new_n49564_;
  assign new_n49566_ = \b[54]  & ~new_n48833_;
  assign new_n49567_ = ~new_n48831_ & new_n49566_;
  assign new_n49568_ = ~new_n48835_ & ~new_n49567_;
  assign new_n49569_ = ~new_n49565_ & new_n49568_;
  assign new_n49570_ = ~new_n48835_ & ~new_n49569_;
  assign new_n49571_ = new_n21537_ & ~new_n49570_;
  assign new_n49572_ = ~new_n48824_ & ~new_n49571_;
  assign new_n49573_ = ~new_n48845_ & new_n49563_;
  assign new_n49574_ = ~new_n49559_ & new_n49573_;
  assign new_n49575_ = ~new_n49560_ & ~new_n49563_;
  assign new_n49576_ = ~new_n49574_ & ~new_n49575_;
  assign new_n49577_ = new_n21537_ & ~new_n49576_;
  assign new_n49578_ = ~new_n49570_ & new_n49577_;
  assign new_n49579_ = ~new_n49572_ & ~new_n49578_;
  assign new_n49580_ = ~\b[54]  & ~new_n49579_;
  assign new_n49581_ = ~new_n48844_ & ~new_n49571_;
  assign new_n49582_ = ~new_n48854_ & new_n49558_;
  assign new_n49583_ = ~new_n49554_ & new_n49582_;
  assign new_n49584_ = ~new_n49555_ & ~new_n49558_;
  assign new_n49585_ = ~new_n49583_ & ~new_n49584_;
  assign new_n49586_ = new_n21537_ & ~new_n49585_;
  assign new_n49587_ = ~new_n49570_ & new_n49586_;
  assign new_n49588_ = ~new_n49581_ & ~new_n49587_;
  assign new_n49589_ = ~\b[53]  & ~new_n49588_;
  assign new_n49590_ = ~new_n48853_ & ~new_n49571_;
  assign new_n49591_ = ~new_n48863_ & new_n49553_;
  assign new_n49592_ = ~new_n49549_ & new_n49591_;
  assign new_n49593_ = ~new_n49550_ & ~new_n49553_;
  assign new_n49594_ = ~new_n49592_ & ~new_n49593_;
  assign new_n49595_ = new_n21537_ & ~new_n49594_;
  assign new_n49596_ = ~new_n49570_ & new_n49595_;
  assign new_n49597_ = ~new_n49590_ & ~new_n49596_;
  assign new_n49598_ = ~\b[52]  & ~new_n49597_;
  assign new_n49599_ = ~new_n48862_ & ~new_n49571_;
  assign new_n49600_ = ~new_n48872_ & new_n49548_;
  assign new_n49601_ = ~new_n49544_ & new_n49600_;
  assign new_n49602_ = ~new_n49545_ & ~new_n49548_;
  assign new_n49603_ = ~new_n49601_ & ~new_n49602_;
  assign new_n49604_ = new_n21537_ & ~new_n49603_;
  assign new_n49605_ = ~new_n49570_ & new_n49604_;
  assign new_n49606_ = ~new_n49599_ & ~new_n49605_;
  assign new_n49607_ = ~\b[51]  & ~new_n49606_;
  assign new_n49608_ = ~new_n48871_ & ~new_n49571_;
  assign new_n49609_ = ~new_n48881_ & new_n49543_;
  assign new_n49610_ = ~new_n49539_ & new_n49609_;
  assign new_n49611_ = ~new_n49540_ & ~new_n49543_;
  assign new_n49612_ = ~new_n49610_ & ~new_n49611_;
  assign new_n49613_ = new_n21537_ & ~new_n49612_;
  assign new_n49614_ = ~new_n49570_ & new_n49613_;
  assign new_n49615_ = ~new_n49608_ & ~new_n49614_;
  assign new_n49616_ = ~\b[50]  & ~new_n49615_;
  assign new_n49617_ = ~new_n48880_ & ~new_n49571_;
  assign new_n49618_ = ~new_n48890_ & new_n49538_;
  assign new_n49619_ = ~new_n49534_ & new_n49618_;
  assign new_n49620_ = ~new_n49535_ & ~new_n49538_;
  assign new_n49621_ = ~new_n49619_ & ~new_n49620_;
  assign new_n49622_ = new_n21537_ & ~new_n49621_;
  assign new_n49623_ = ~new_n49570_ & new_n49622_;
  assign new_n49624_ = ~new_n49617_ & ~new_n49623_;
  assign new_n49625_ = ~\b[49]  & ~new_n49624_;
  assign new_n49626_ = ~new_n48889_ & ~new_n49571_;
  assign new_n49627_ = ~new_n48899_ & new_n49533_;
  assign new_n49628_ = ~new_n49529_ & new_n49627_;
  assign new_n49629_ = ~new_n49530_ & ~new_n49533_;
  assign new_n49630_ = ~new_n49628_ & ~new_n49629_;
  assign new_n49631_ = new_n21537_ & ~new_n49630_;
  assign new_n49632_ = ~new_n49570_ & new_n49631_;
  assign new_n49633_ = ~new_n49626_ & ~new_n49632_;
  assign new_n49634_ = ~\b[48]  & ~new_n49633_;
  assign new_n49635_ = ~new_n48898_ & ~new_n49571_;
  assign new_n49636_ = ~new_n48908_ & new_n49528_;
  assign new_n49637_ = ~new_n49524_ & new_n49636_;
  assign new_n49638_ = ~new_n49525_ & ~new_n49528_;
  assign new_n49639_ = ~new_n49637_ & ~new_n49638_;
  assign new_n49640_ = new_n21537_ & ~new_n49639_;
  assign new_n49641_ = ~new_n49570_ & new_n49640_;
  assign new_n49642_ = ~new_n49635_ & ~new_n49641_;
  assign new_n49643_ = ~\b[47]  & ~new_n49642_;
  assign new_n49644_ = ~new_n48907_ & ~new_n49571_;
  assign new_n49645_ = ~new_n48917_ & new_n49523_;
  assign new_n49646_ = ~new_n49519_ & new_n49645_;
  assign new_n49647_ = ~new_n49520_ & ~new_n49523_;
  assign new_n49648_ = ~new_n49646_ & ~new_n49647_;
  assign new_n49649_ = new_n21537_ & ~new_n49648_;
  assign new_n49650_ = ~new_n49570_ & new_n49649_;
  assign new_n49651_ = ~new_n49644_ & ~new_n49650_;
  assign new_n49652_ = ~\b[46]  & ~new_n49651_;
  assign new_n49653_ = ~new_n48916_ & ~new_n49571_;
  assign new_n49654_ = ~new_n48926_ & new_n49518_;
  assign new_n49655_ = ~new_n49514_ & new_n49654_;
  assign new_n49656_ = ~new_n49515_ & ~new_n49518_;
  assign new_n49657_ = ~new_n49655_ & ~new_n49656_;
  assign new_n49658_ = new_n21537_ & ~new_n49657_;
  assign new_n49659_ = ~new_n49570_ & new_n49658_;
  assign new_n49660_ = ~new_n49653_ & ~new_n49659_;
  assign new_n49661_ = ~\b[45]  & ~new_n49660_;
  assign new_n49662_ = ~new_n48925_ & ~new_n49571_;
  assign new_n49663_ = ~new_n48935_ & new_n49513_;
  assign new_n49664_ = ~new_n49509_ & new_n49663_;
  assign new_n49665_ = ~new_n49510_ & ~new_n49513_;
  assign new_n49666_ = ~new_n49664_ & ~new_n49665_;
  assign new_n49667_ = new_n21537_ & ~new_n49666_;
  assign new_n49668_ = ~new_n49570_ & new_n49667_;
  assign new_n49669_ = ~new_n49662_ & ~new_n49668_;
  assign new_n49670_ = ~\b[44]  & ~new_n49669_;
  assign new_n49671_ = ~new_n48934_ & ~new_n49571_;
  assign new_n49672_ = ~new_n48944_ & new_n49508_;
  assign new_n49673_ = ~new_n49504_ & new_n49672_;
  assign new_n49674_ = ~new_n49505_ & ~new_n49508_;
  assign new_n49675_ = ~new_n49673_ & ~new_n49674_;
  assign new_n49676_ = new_n21537_ & ~new_n49675_;
  assign new_n49677_ = ~new_n49570_ & new_n49676_;
  assign new_n49678_ = ~new_n49671_ & ~new_n49677_;
  assign new_n49679_ = ~\b[43]  & ~new_n49678_;
  assign new_n49680_ = ~new_n48943_ & ~new_n49571_;
  assign new_n49681_ = ~new_n48953_ & new_n49503_;
  assign new_n49682_ = ~new_n49499_ & new_n49681_;
  assign new_n49683_ = ~new_n49500_ & ~new_n49503_;
  assign new_n49684_ = ~new_n49682_ & ~new_n49683_;
  assign new_n49685_ = new_n21537_ & ~new_n49684_;
  assign new_n49686_ = ~new_n49570_ & new_n49685_;
  assign new_n49687_ = ~new_n49680_ & ~new_n49686_;
  assign new_n49688_ = ~\b[42]  & ~new_n49687_;
  assign new_n49689_ = ~new_n48952_ & ~new_n49571_;
  assign new_n49690_ = ~new_n48962_ & new_n49498_;
  assign new_n49691_ = ~new_n49494_ & new_n49690_;
  assign new_n49692_ = ~new_n49495_ & ~new_n49498_;
  assign new_n49693_ = ~new_n49691_ & ~new_n49692_;
  assign new_n49694_ = new_n21537_ & ~new_n49693_;
  assign new_n49695_ = ~new_n49570_ & new_n49694_;
  assign new_n49696_ = ~new_n49689_ & ~new_n49695_;
  assign new_n49697_ = ~\b[41]  & ~new_n49696_;
  assign new_n49698_ = ~new_n48961_ & ~new_n49571_;
  assign new_n49699_ = ~new_n48971_ & new_n49493_;
  assign new_n49700_ = ~new_n49489_ & new_n49699_;
  assign new_n49701_ = ~new_n49490_ & ~new_n49493_;
  assign new_n49702_ = ~new_n49700_ & ~new_n49701_;
  assign new_n49703_ = new_n21537_ & ~new_n49702_;
  assign new_n49704_ = ~new_n49570_ & new_n49703_;
  assign new_n49705_ = ~new_n49698_ & ~new_n49704_;
  assign new_n49706_ = ~\b[40]  & ~new_n49705_;
  assign new_n49707_ = ~new_n48970_ & ~new_n49571_;
  assign new_n49708_ = ~new_n48980_ & new_n49488_;
  assign new_n49709_ = ~new_n49484_ & new_n49708_;
  assign new_n49710_ = ~new_n49485_ & ~new_n49488_;
  assign new_n49711_ = ~new_n49709_ & ~new_n49710_;
  assign new_n49712_ = new_n21537_ & ~new_n49711_;
  assign new_n49713_ = ~new_n49570_ & new_n49712_;
  assign new_n49714_ = ~new_n49707_ & ~new_n49713_;
  assign new_n49715_ = ~\b[39]  & ~new_n49714_;
  assign new_n49716_ = ~new_n48979_ & ~new_n49571_;
  assign new_n49717_ = ~new_n48989_ & new_n49483_;
  assign new_n49718_ = ~new_n49479_ & new_n49717_;
  assign new_n49719_ = ~new_n49480_ & ~new_n49483_;
  assign new_n49720_ = ~new_n49718_ & ~new_n49719_;
  assign new_n49721_ = new_n21537_ & ~new_n49720_;
  assign new_n49722_ = ~new_n49570_ & new_n49721_;
  assign new_n49723_ = ~new_n49716_ & ~new_n49722_;
  assign new_n49724_ = ~\b[38]  & ~new_n49723_;
  assign new_n49725_ = ~new_n48988_ & ~new_n49571_;
  assign new_n49726_ = ~new_n48998_ & new_n49478_;
  assign new_n49727_ = ~new_n49474_ & new_n49726_;
  assign new_n49728_ = ~new_n49475_ & ~new_n49478_;
  assign new_n49729_ = ~new_n49727_ & ~new_n49728_;
  assign new_n49730_ = new_n21537_ & ~new_n49729_;
  assign new_n49731_ = ~new_n49570_ & new_n49730_;
  assign new_n49732_ = ~new_n49725_ & ~new_n49731_;
  assign new_n49733_ = ~\b[37]  & ~new_n49732_;
  assign new_n49734_ = ~new_n48997_ & ~new_n49571_;
  assign new_n49735_ = ~new_n49007_ & new_n49473_;
  assign new_n49736_ = ~new_n49469_ & new_n49735_;
  assign new_n49737_ = ~new_n49470_ & ~new_n49473_;
  assign new_n49738_ = ~new_n49736_ & ~new_n49737_;
  assign new_n49739_ = new_n21537_ & ~new_n49738_;
  assign new_n49740_ = ~new_n49570_ & new_n49739_;
  assign new_n49741_ = ~new_n49734_ & ~new_n49740_;
  assign new_n49742_ = ~\b[36]  & ~new_n49741_;
  assign new_n49743_ = ~new_n49006_ & ~new_n49571_;
  assign new_n49744_ = ~new_n49016_ & new_n49468_;
  assign new_n49745_ = ~new_n49464_ & new_n49744_;
  assign new_n49746_ = ~new_n49465_ & ~new_n49468_;
  assign new_n49747_ = ~new_n49745_ & ~new_n49746_;
  assign new_n49748_ = new_n21537_ & ~new_n49747_;
  assign new_n49749_ = ~new_n49570_ & new_n49748_;
  assign new_n49750_ = ~new_n49743_ & ~new_n49749_;
  assign new_n49751_ = ~\b[35]  & ~new_n49750_;
  assign new_n49752_ = ~new_n49015_ & ~new_n49571_;
  assign new_n49753_ = ~new_n49025_ & new_n49463_;
  assign new_n49754_ = ~new_n49459_ & new_n49753_;
  assign new_n49755_ = ~new_n49460_ & ~new_n49463_;
  assign new_n49756_ = ~new_n49754_ & ~new_n49755_;
  assign new_n49757_ = new_n21537_ & ~new_n49756_;
  assign new_n49758_ = ~new_n49570_ & new_n49757_;
  assign new_n49759_ = ~new_n49752_ & ~new_n49758_;
  assign new_n49760_ = ~\b[34]  & ~new_n49759_;
  assign new_n49761_ = ~new_n49024_ & ~new_n49571_;
  assign new_n49762_ = ~new_n49034_ & new_n49458_;
  assign new_n49763_ = ~new_n49454_ & new_n49762_;
  assign new_n49764_ = ~new_n49455_ & ~new_n49458_;
  assign new_n49765_ = ~new_n49763_ & ~new_n49764_;
  assign new_n49766_ = new_n21537_ & ~new_n49765_;
  assign new_n49767_ = ~new_n49570_ & new_n49766_;
  assign new_n49768_ = ~new_n49761_ & ~new_n49767_;
  assign new_n49769_ = ~\b[33]  & ~new_n49768_;
  assign new_n49770_ = ~new_n49033_ & ~new_n49571_;
  assign new_n49771_ = ~new_n49043_ & new_n49453_;
  assign new_n49772_ = ~new_n49449_ & new_n49771_;
  assign new_n49773_ = ~new_n49450_ & ~new_n49453_;
  assign new_n49774_ = ~new_n49772_ & ~new_n49773_;
  assign new_n49775_ = new_n21537_ & ~new_n49774_;
  assign new_n49776_ = ~new_n49570_ & new_n49775_;
  assign new_n49777_ = ~new_n49770_ & ~new_n49776_;
  assign new_n49778_ = ~\b[32]  & ~new_n49777_;
  assign new_n49779_ = ~new_n49042_ & ~new_n49571_;
  assign new_n49780_ = ~new_n49052_ & new_n49448_;
  assign new_n49781_ = ~new_n49444_ & new_n49780_;
  assign new_n49782_ = ~new_n49445_ & ~new_n49448_;
  assign new_n49783_ = ~new_n49781_ & ~new_n49782_;
  assign new_n49784_ = new_n21537_ & ~new_n49783_;
  assign new_n49785_ = ~new_n49570_ & new_n49784_;
  assign new_n49786_ = ~new_n49779_ & ~new_n49785_;
  assign new_n49787_ = ~\b[31]  & ~new_n49786_;
  assign new_n49788_ = ~new_n49051_ & ~new_n49571_;
  assign new_n49789_ = ~new_n49061_ & new_n49443_;
  assign new_n49790_ = ~new_n49439_ & new_n49789_;
  assign new_n49791_ = ~new_n49440_ & ~new_n49443_;
  assign new_n49792_ = ~new_n49790_ & ~new_n49791_;
  assign new_n49793_ = new_n21537_ & ~new_n49792_;
  assign new_n49794_ = ~new_n49570_ & new_n49793_;
  assign new_n49795_ = ~new_n49788_ & ~new_n49794_;
  assign new_n49796_ = ~\b[30]  & ~new_n49795_;
  assign new_n49797_ = ~new_n49060_ & ~new_n49571_;
  assign new_n49798_ = ~new_n49070_ & new_n49438_;
  assign new_n49799_ = ~new_n49434_ & new_n49798_;
  assign new_n49800_ = ~new_n49435_ & ~new_n49438_;
  assign new_n49801_ = ~new_n49799_ & ~new_n49800_;
  assign new_n49802_ = new_n21537_ & ~new_n49801_;
  assign new_n49803_ = ~new_n49570_ & new_n49802_;
  assign new_n49804_ = ~new_n49797_ & ~new_n49803_;
  assign new_n49805_ = ~\b[29]  & ~new_n49804_;
  assign new_n49806_ = ~new_n49069_ & ~new_n49571_;
  assign new_n49807_ = ~new_n49079_ & new_n49433_;
  assign new_n49808_ = ~new_n49429_ & new_n49807_;
  assign new_n49809_ = ~new_n49430_ & ~new_n49433_;
  assign new_n49810_ = ~new_n49808_ & ~new_n49809_;
  assign new_n49811_ = new_n21537_ & ~new_n49810_;
  assign new_n49812_ = ~new_n49570_ & new_n49811_;
  assign new_n49813_ = ~new_n49806_ & ~new_n49812_;
  assign new_n49814_ = ~\b[28]  & ~new_n49813_;
  assign new_n49815_ = ~new_n49078_ & ~new_n49571_;
  assign new_n49816_ = ~new_n49088_ & new_n49428_;
  assign new_n49817_ = ~new_n49424_ & new_n49816_;
  assign new_n49818_ = ~new_n49425_ & ~new_n49428_;
  assign new_n49819_ = ~new_n49817_ & ~new_n49818_;
  assign new_n49820_ = new_n21537_ & ~new_n49819_;
  assign new_n49821_ = ~new_n49570_ & new_n49820_;
  assign new_n49822_ = ~new_n49815_ & ~new_n49821_;
  assign new_n49823_ = ~\b[27]  & ~new_n49822_;
  assign new_n49824_ = ~new_n49087_ & ~new_n49571_;
  assign new_n49825_ = ~new_n49097_ & new_n49423_;
  assign new_n49826_ = ~new_n49419_ & new_n49825_;
  assign new_n49827_ = ~new_n49420_ & ~new_n49423_;
  assign new_n49828_ = ~new_n49826_ & ~new_n49827_;
  assign new_n49829_ = new_n21537_ & ~new_n49828_;
  assign new_n49830_ = ~new_n49570_ & new_n49829_;
  assign new_n49831_ = ~new_n49824_ & ~new_n49830_;
  assign new_n49832_ = ~\b[26]  & ~new_n49831_;
  assign new_n49833_ = ~new_n49096_ & ~new_n49571_;
  assign new_n49834_ = ~new_n49106_ & new_n49418_;
  assign new_n49835_ = ~new_n49414_ & new_n49834_;
  assign new_n49836_ = ~new_n49415_ & ~new_n49418_;
  assign new_n49837_ = ~new_n49835_ & ~new_n49836_;
  assign new_n49838_ = new_n21537_ & ~new_n49837_;
  assign new_n49839_ = ~new_n49570_ & new_n49838_;
  assign new_n49840_ = ~new_n49833_ & ~new_n49839_;
  assign new_n49841_ = ~\b[25]  & ~new_n49840_;
  assign new_n49842_ = ~new_n49105_ & ~new_n49571_;
  assign new_n49843_ = ~new_n49115_ & new_n49413_;
  assign new_n49844_ = ~new_n49409_ & new_n49843_;
  assign new_n49845_ = ~new_n49410_ & ~new_n49413_;
  assign new_n49846_ = ~new_n49844_ & ~new_n49845_;
  assign new_n49847_ = new_n21537_ & ~new_n49846_;
  assign new_n49848_ = ~new_n49570_ & new_n49847_;
  assign new_n49849_ = ~new_n49842_ & ~new_n49848_;
  assign new_n49850_ = ~\b[24]  & ~new_n49849_;
  assign new_n49851_ = ~new_n49114_ & ~new_n49571_;
  assign new_n49852_ = ~new_n49124_ & new_n49408_;
  assign new_n49853_ = ~new_n49404_ & new_n49852_;
  assign new_n49854_ = ~new_n49405_ & ~new_n49408_;
  assign new_n49855_ = ~new_n49853_ & ~new_n49854_;
  assign new_n49856_ = new_n21537_ & ~new_n49855_;
  assign new_n49857_ = ~new_n49570_ & new_n49856_;
  assign new_n49858_ = ~new_n49851_ & ~new_n49857_;
  assign new_n49859_ = ~\b[23]  & ~new_n49858_;
  assign new_n49860_ = ~new_n49123_ & ~new_n49571_;
  assign new_n49861_ = ~new_n49133_ & new_n49403_;
  assign new_n49862_ = ~new_n49399_ & new_n49861_;
  assign new_n49863_ = ~new_n49400_ & ~new_n49403_;
  assign new_n49864_ = ~new_n49862_ & ~new_n49863_;
  assign new_n49865_ = new_n21537_ & ~new_n49864_;
  assign new_n49866_ = ~new_n49570_ & new_n49865_;
  assign new_n49867_ = ~new_n49860_ & ~new_n49866_;
  assign new_n49868_ = ~\b[22]  & ~new_n49867_;
  assign new_n49869_ = ~new_n49132_ & ~new_n49571_;
  assign new_n49870_ = ~new_n49142_ & new_n49398_;
  assign new_n49871_ = ~new_n49394_ & new_n49870_;
  assign new_n49872_ = ~new_n49395_ & ~new_n49398_;
  assign new_n49873_ = ~new_n49871_ & ~new_n49872_;
  assign new_n49874_ = new_n21537_ & ~new_n49873_;
  assign new_n49875_ = ~new_n49570_ & new_n49874_;
  assign new_n49876_ = ~new_n49869_ & ~new_n49875_;
  assign new_n49877_ = ~\b[21]  & ~new_n49876_;
  assign new_n49878_ = ~new_n49141_ & ~new_n49571_;
  assign new_n49879_ = ~new_n49151_ & new_n49393_;
  assign new_n49880_ = ~new_n49389_ & new_n49879_;
  assign new_n49881_ = ~new_n49390_ & ~new_n49393_;
  assign new_n49882_ = ~new_n49880_ & ~new_n49881_;
  assign new_n49883_ = new_n21537_ & ~new_n49882_;
  assign new_n49884_ = ~new_n49570_ & new_n49883_;
  assign new_n49885_ = ~new_n49878_ & ~new_n49884_;
  assign new_n49886_ = ~\b[20]  & ~new_n49885_;
  assign new_n49887_ = ~new_n49150_ & ~new_n49571_;
  assign new_n49888_ = ~new_n49160_ & new_n49388_;
  assign new_n49889_ = ~new_n49384_ & new_n49888_;
  assign new_n49890_ = ~new_n49385_ & ~new_n49388_;
  assign new_n49891_ = ~new_n49889_ & ~new_n49890_;
  assign new_n49892_ = new_n21537_ & ~new_n49891_;
  assign new_n49893_ = ~new_n49570_ & new_n49892_;
  assign new_n49894_ = ~new_n49887_ & ~new_n49893_;
  assign new_n49895_ = ~\b[19]  & ~new_n49894_;
  assign new_n49896_ = ~new_n49159_ & ~new_n49571_;
  assign new_n49897_ = ~new_n49169_ & new_n49383_;
  assign new_n49898_ = ~new_n49379_ & new_n49897_;
  assign new_n49899_ = ~new_n49380_ & ~new_n49383_;
  assign new_n49900_ = ~new_n49898_ & ~new_n49899_;
  assign new_n49901_ = new_n21537_ & ~new_n49900_;
  assign new_n49902_ = ~new_n49570_ & new_n49901_;
  assign new_n49903_ = ~new_n49896_ & ~new_n49902_;
  assign new_n49904_ = ~\b[18]  & ~new_n49903_;
  assign new_n49905_ = ~new_n49168_ & ~new_n49571_;
  assign new_n49906_ = ~new_n49178_ & new_n49378_;
  assign new_n49907_ = ~new_n49374_ & new_n49906_;
  assign new_n49908_ = ~new_n49375_ & ~new_n49378_;
  assign new_n49909_ = ~new_n49907_ & ~new_n49908_;
  assign new_n49910_ = new_n21537_ & ~new_n49909_;
  assign new_n49911_ = ~new_n49570_ & new_n49910_;
  assign new_n49912_ = ~new_n49905_ & ~new_n49911_;
  assign new_n49913_ = ~\b[17]  & ~new_n49912_;
  assign new_n49914_ = ~new_n49177_ & ~new_n49571_;
  assign new_n49915_ = ~new_n49187_ & new_n49373_;
  assign new_n49916_ = ~new_n49369_ & new_n49915_;
  assign new_n49917_ = ~new_n49370_ & ~new_n49373_;
  assign new_n49918_ = ~new_n49916_ & ~new_n49917_;
  assign new_n49919_ = new_n21537_ & ~new_n49918_;
  assign new_n49920_ = ~new_n49570_ & new_n49919_;
  assign new_n49921_ = ~new_n49914_ & ~new_n49920_;
  assign new_n49922_ = ~\b[16]  & ~new_n49921_;
  assign new_n49923_ = ~new_n49186_ & ~new_n49571_;
  assign new_n49924_ = ~new_n49196_ & new_n49368_;
  assign new_n49925_ = ~new_n49364_ & new_n49924_;
  assign new_n49926_ = ~new_n49365_ & ~new_n49368_;
  assign new_n49927_ = ~new_n49925_ & ~new_n49926_;
  assign new_n49928_ = new_n21537_ & ~new_n49927_;
  assign new_n49929_ = ~new_n49570_ & new_n49928_;
  assign new_n49930_ = ~new_n49923_ & ~new_n49929_;
  assign new_n49931_ = ~\b[15]  & ~new_n49930_;
  assign new_n49932_ = ~new_n49195_ & ~new_n49571_;
  assign new_n49933_ = ~new_n49205_ & new_n49363_;
  assign new_n49934_ = ~new_n49359_ & new_n49933_;
  assign new_n49935_ = ~new_n49360_ & ~new_n49363_;
  assign new_n49936_ = ~new_n49934_ & ~new_n49935_;
  assign new_n49937_ = new_n21537_ & ~new_n49936_;
  assign new_n49938_ = ~new_n49570_ & new_n49937_;
  assign new_n49939_ = ~new_n49932_ & ~new_n49938_;
  assign new_n49940_ = ~\b[14]  & ~new_n49939_;
  assign new_n49941_ = ~new_n49204_ & ~new_n49571_;
  assign new_n49942_ = ~new_n49214_ & new_n49358_;
  assign new_n49943_ = ~new_n49354_ & new_n49942_;
  assign new_n49944_ = ~new_n49355_ & ~new_n49358_;
  assign new_n49945_ = ~new_n49943_ & ~new_n49944_;
  assign new_n49946_ = new_n21537_ & ~new_n49945_;
  assign new_n49947_ = ~new_n49570_ & new_n49946_;
  assign new_n49948_ = ~new_n49941_ & ~new_n49947_;
  assign new_n49949_ = ~\b[13]  & ~new_n49948_;
  assign new_n49950_ = ~new_n49213_ & ~new_n49571_;
  assign new_n49951_ = ~new_n49223_ & new_n49353_;
  assign new_n49952_ = ~new_n49349_ & new_n49951_;
  assign new_n49953_ = ~new_n49350_ & ~new_n49353_;
  assign new_n49954_ = ~new_n49952_ & ~new_n49953_;
  assign new_n49955_ = new_n21537_ & ~new_n49954_;
  assign new_n49956_ = ~new_n49570_ & new_n49955_;
  assign new_n49957_ = ~new_n49950_ & ~new_n49956_;
  assign new_n49958_ = ~\b[12]  & ~new_n49957_;
  assign new_n49959_ = ~new_n49222_ & ~new_n49571_;
  assign new_n49960_ = ~new_n49232_ & new_n49348_;
  assign new_n49961_ = ~new_n49344_ & new_n49960_;
  assign new_n49962_ = ~new_n49345_ & ~new_n49348_;
  assign new_n49963_ = ~new_n49961_ & ~new_n49962_;
  assign new_n49964_ = new_n21537_ & ~new_n49963_;
  assign new_n49965_ = ~new_n49570_ & new_n49964_;
  assign new_n49966_ = ~new_n49959_ & ~new_n49965_;
  assign new_n49967_ = ~\b[11]  & ~new_n49966_;
  assign new_n49968_ = ~new_n49231_ & ~new_n49571_;
  assign new_n49969_ = ~new_n49241_ & new_n49343_;
  assign new_n49970_ = ~new_n49339_ & new_n49969_;
  assign new_n49971_ = ~new_n49340_ & ~new_n49343_;
  assign new_n49972_ = ~new_n49970_ & ~new_n49971_;
  assign new_n49973_ = new_n21537_ & ~new_n49972_;
  assign new_n49974_ = ~new_n49570_ & new_n49973_;
  assign new_n49975_ = ~new_n49968_ & ~new_n49974_;
  assign new_n49976_ = ~\b[10]  & ~new_n49975_;
  assign new_n49977_ = ~new_n49240_ & ~new_n49571_;
  assign new_n49978_ = ~new_n49250_ & new_n49338_;
  assign new_n49979_ = ~new_n49334_ & new_n49978_;
  assign new_n49980_ = ~new_n49335_ & ~new_n49338_;
  assign new_n49981_ = ~new_n49979_ & ~new_n49980_;
  assign new_n49982_ = new_n21537_ & ~new_n49981_;
  assign new_n49983_ = ~new_n49570_ & new_n49982_;
  assign new_n49984_ = ~new_n49977_ & ~new_n49983_;
  assign new_n49985_ = ~\b[9]  & ~new_n49984_;
  assign new_n49986_ = ~new_n49249_ & ~new_n49571_;
  assign new_n49987_ = ~new_n49259_ & new_n49333_;
  assign new_n49988_ = ~new_n49329_ & new_n49987_;
  assign new_n49989_ = ~new_n49330_ & ~new_n49333_;
  assign new_n49990_ = ~new_n49988_ & ~new_n49989_;
  assign new_n49991_ = new_n21537_ & ~new_n49990_;
  assign new_n49992_ = ~new_n49570_ & new_n49991_;
  assign new_n49993_ = ~new_n49986_ & ~new_n49992_;
  assign new_n49994_ = ~\b[8]  & ~new_n49993_;
  assign new_n49995_ = ~new_n49258_ & ~new_n49571_;
  assign new_n49996_ = ~new_n49268_ & new_n49328_;
  assign new_n49997_ = ~new_n49324_ & new_n49996_;
  assign new_n49998_ = ~new_n49325_ & ~new_n49328_;
  assign new_n49999_ = ~new_n49997_ & ~new_n49998_;
  assign new_n50000_ = new_n21537_ & ~new_n49999_;
  assign new_n50001_ = ~new_n49570_ & new_n50000_;
  assign new_n50002_ = ~new_n49995_ & ~new_n50001_;
  assign new_n50003_ = ~\b[7]  & ~new_n50002_;
  assign new_n50004_ = ~new_n49267_ & ~new_n49571_;
  assign new_n50005_ = ~new_n49277_ & new_n49323_;
  assign new_n50006_ = ~new_n49319_ & new_n50005_;
  assign new_n50007_ = ~new_n49320_ & ~new_n49323_;
  assign new_n50008_ = ~new_n50006_ & ~new_n50007_;
  assign new_n50009_ = new_n21537_ & ~new_n50008_;
  assign new_n50010_ = ~new_n49570_ & new_n50009_;
  assign new_n50011_ = ~new_n50004_ & ~new_n50010_;
  assign new_n50012_ = ~\b[6]  & ~new_n50011_;
  assign new_n50013_ = ~new_n49276_ & ~new_n49571_;
  assign new_n50014_ = ~new_n49286_ & new_n49318_;
  assign new_n50015_ = ~new_n49314_ & new_n50014_;
  assign new_n50016_ = ~new_n49315_ & ~new_n49318_;
  assign new_n50017_ = ~new_n50015_ & ~new_n50016_;
  assign new_n50018_ = new_n21537_ & ~new_n50017_;
  assign new_n50019_ = ~new_n49570_ & new_n50018_;
  assign new_n50020_ = ~new_n50013_ & ~new_n50019_;
  assign new_n50021_ = ~\b[5]  & ~new_n50020_;
  assign new_n50022_ = ~new_n49285_ & ~new_n49571_;
  assign new_n50023_ = ~new_n49294_ & new_n49313_;
  assign new_n50024_ = ~new_n49309_ & new_n50023_;
  assign new_n50025_ = ~new_n49310_ & ~new_n49313_;
  assign new_n50026_ = ~new_n50024_ & ~new_n50025_;
  assign new_n50027_ = new_n21537_ & ~new_n50026_;
  assign new_n50028_ = ~new_n49570_ & new_n50027_;
  assign new_n50029_ = ~new_n50022_ & ~new_n50028_;
  assign new_n50030_ = ~\b[4]  & ~new_n50029_;
  assign new_n50031_ = ~new_n49293_ & ~new_n49571_;
  assign new_n50032_ = ~new_n49304_ & new_n49308_;
  assign new_n50033_ = ~new_n49303_ & new_n50032_;
  assign new_n50034_ = ~new_n49305_ & ~new_n49308_;
  assign new_n50035_ = ~new_n50033_ & ~new_n50034_;
  assign new_n50036_ = new_n21537_ & ~new_n50035_;
  assign new_n50037_ = ~new_n49570_ & new_n50036_;
  assign new_n50038_ = ~new_n50031_ & ~new_n50037_;
  assign new_n50039_ = ~\b[3]  & ~new_n50038_;
  assign new_n50040_ = ~new_n49298_ & ~new_n49571_;
  assign new_n50041_ = new_n21267_ & ~new_n49301_;
  assign new_n50042_ = ~new_n49299_ & new_n50041_;
  assign new_n50043_ = new_n21537_ & ~new_n50042_;
  assign new_n50044_ = ~new_n49303_ & new_n50043_;
  assign new_n50045_ = ~new_n49570_ & new_n50044_;
  assign new_n50046_ = ~new_n50040_ & ~new_n50045_;
  assign new_n50047_ = ~\b[2]  & ~new_n50046_;
  assign new_n50048_ = new_n22017_ & ~new_n49570_;
  assign new_n50049_ = \a[9]  & ~new_n50048_;
  assign new_n50050_ = new_n22022_ & ~new_n49570_;
  assign new_n50051_ = ~new_n50049_ & ~new_n50050_;
  assign new_n50052_ = \b[1]  & ~new_n50051_;
  assign new_n50053_ = ~\b[1]  & ~new_n50050_;
  assign new_n50054_ = ~new_n50049_ & new_n50053_;
  assign new_n50055_ = ~new_n50052_ & ~new_n50054_;
  assign new_n50056_ = ~new_n22029_ & ~new_n50055_;
  assign new_n50057_ = ~\b[1]  & ~new_n50051_;
  assign new_n50058_ = ~new_n50056_ & ~new_n50057_;
  assign new_n50059_ = \b[2]  & ~new_n50045_;
  assign new_n50060_ = ~new_n50040_ & new_n50059_;
  assign new_n50061_ = ~new_n50047_ & ~new_n50060_;
  assign new_n50062_ = ~new_n50058_ & new_n50061_;
  assign new_n50063_ = ~new_n50047_ & ~new_n50062_;
  assign new_n50064_ = \b[3]  & ~new_n50037_;
  assign new_n50065_ = ~new_n50031_ & new_n50064_;
  assign new_n50066_ = ~new_n50039_ & ~new_n50065_;
  assign new_n50067_ = ~new_n50063_ & new_n50066_;
  assign new_n50068_ = ~new_n50039_ & ~new_n50067_;
  assign new_n50069_ = \b[4]  & ~new_n50028_;
  assign new_n50070_ = ~new_n50022_ & new_n50069_;
  assign new_n50071_ = ~new_n50030_ & ~new_n50070_;
  assign new_n50072_ = ~new_n50068_ & new_n50071_;
  assign new_n50073_ = ~new_n50030_ & ~new_n50072_;
  assign new_n50074_ = \b[5]  & ~new_n50019_;
  assign new_n50075_ = ~new_n50013_ & new_n50074_;
  assign new_n50076_ = ~new_n50021_ & ~new_n50075_;
  assign new_n50077_ = ~new_n50073_ & new_n50076_;
  assign new_n50078_ = ~new_n50021_ & ~new_n50077_;
  assign new_n50079_ = \b[6]  & ~new_n50010_;
  assign new_n50080_ = ~new_n50004_ & new_n50079_;
  assign new_n50081_ = ~new_n50012_ & ~new_n50080_;
  assign new_n50082_ = ~new_n50078_ & new_n50081_;
  assign new_n50083_ = ~new_n50012_ & ~new_n50082_;
  assign new_n50084_ = \b[7]  & ~new_n50001_;
  assign new_n50085_ = ~new_n49995_ & new_n50084_;
  assign new_n50086_ = ~new_n50003_ & ~new_n50085_;
  assign new_n50087_ = ~new_n50083_ & new_n50086_;
  assign new_n50088_ = ~new_n50003_ & ~new_n50087_;
  assign new_n50089_ = \b[8]  & ~new_n49992_;
  assign new_n50090_ = ~new_n49986_ & new_n50089_;
  assign new_n50091_ = ~new_n49994_ & ~new_n50090_;
  assign new_n50092_ = ~new_n50088_ & new_n50091_;
  assign new_n50093_ = ~new_n49994_ & ~new_n50092_;
  assign new_n50094_ = \b[9]  & ~new_n49983_;
  assign new_n50095_ = ~new_n49977_ & new_n50094_;
  assign new_n50096_ = ~new_n49985_ & ~new_n50095_;
  assign new_n50097_ = ~new_n50093_ & new_n50096_;
  assign new_n50098_ = ~new_n49985_ & ~new_n50097_;
  assign new_n50099_ = \b[10]  & ~new_n49974_;
  assign new_n50100_ = ~new_n49968_ & new_n50099_;
  assign new_n50101_ = ~new_n49976_ & ~new_n50100_;
  assign new_n50102_ = ~new_n50098_ & new_n50101_;
  assign new_n50103_ = ~new_n49976_ & ~new_n50102_;
  assign new_n50104_ = \b[11]  & ~new_n49965_;
  assign new_n50105_ = ~new_n49959_ & new_n50104_;
  assign new_n50106_ = ~new_n49967_ & ~new_n50105_;
  assign new_n50107_ = ~new_n50103_ & new_n50106_;
  assign new_n50108_ = ~new_n49967_ & ~new_n50107_;
  assign new_n50109_ = \b[12]  & ~new_n49956_;
  assign new_n50110_ = ~new_n49950_ & new_n50109_;
  assign new_n50111_ = ~new_n49958_ & ~new_n50110_;
  assign new_n50112_ = ~new_n50108_ & new_n50111_;
  assign new_n50113_ = ~new_n49958_ & ~new_n50112_;
  assign new_n50114_ = \b[13]  & ~new_n49947_;
  assign new_n50115_ = ~new_n49941_ & new_n50114_;
  assign new_n50116_ = ~new_n49949_ & ~new_n50115_;
  assign new_n50117_ = ~new_n50113_ & new_n50116_;
  assign new_n50118_ = ~new_n49949_ & ~new_n50117_;
  assign new_n50119_ = \b[14]  & ~new_n49938_;
  assign new_n50120_ = ~new_n49932_ & new_n50119_;
  assign new_n50121_ = ~new_n49940_ & ~new_n50120_;
  assign new_n50122_ = ~new_n50118_ & new_n50121_;
  assign new_n50123_ = ~new_n49940_ & ~new_n50122_;
  assign new_n50124_ = \b[15]  & ~new_n49929_;
  assign new_n50125_ = ~new_n49923_ & new_n50124_;
  assign new_n50126_ = ~new_n49931_ & ~new_n50125_;
  assign new_n50127_ = ~new_n50123_ & new_n50126_;
  assign new_n50128_ = ~new_n49931_ & ~new_n50127_;
  assign new_n50129_ = \b[16]  & ~new_n49920_;
  assign new_n50130_ = ~new_n49914_ & new_n50129_;
  assign new_n50131_ = ~new_n49922_ & ~new_n50130_;
  assign new_n50132_ = ~new_n50128_ & new_n50131_;
  assign new_n50133_ = ~new_n49922_ & ~new_n50132_;
  assign new_n50134_ = \b[17]  & ~new_n49911_;
  assign new_n50135_ = ~new_n49905_ & new_n50134_;
  assign new_n50136_ = ~new_n49913_ & ~new_n50135_;
  assign new_n50137_ = ~new_n50133_ & new_n50136_;
  assign new_n50138_ = ~new_n49913_ & ~new_n50137_;
  assign new_n50139_ = \b[18]  & ~new_n49902_;
  assign new_n50140_ = ~new_n49896_ & new_n50139_;
  assign new_n50141_ = ~new_n49904_ & ~new_n50140_;
  assign new_n50142_ = ~new_n50138_ & new_n50141_;
  assign new_n50143_ = ~new_n49904_ & ~new_n50142_;
  assign new_n50144_ = \b[19]  & ~new_n49893_;
  assign new_n50145_ = ~new_n49887_ & new_n50144_;
  assign new_n50146_ = ~new_n49895_ & ~new_n50145_;
  assign new_n50147_ = ~new_n50143_ & new_n50146_;
  assign new_n50148_ = ~new_n49895_ & ~new_n50147_;
  assign new_n50149_ = \b[20]  & ~new_n49884_;
  assign new_n50150_ = ~new_n49878_ & new_n50149_;
  assign new_n50151_ = ~new_n49886_ & ~new_n50150_;
  assign new_n50152_ = ~new_n50148_ & new_n50151_;
  assign new_n50153_ = ~new_n49886_ & ~new_n50152_;
  assign new_n50154_ = \b[21]  & ~new_n49875_;
  assign new_n50155_ = ~new_n49869_ & new_n50154_;
  assign new_n50156_ = ~new_n49877_ & ~new_n50155_;
  assign new_n50157_ = ~new_n50153_ & new_n50156_;
  assign new_n50158_ = ~new_n49877_ & ~new_n50157_;
  assign new_n50159_ = \b[22]  & ~new_n49866_;
  assign new_n50160_ = ~new_n49860_ & new_n50159_;
  assign new_n50161_ = ~new_n49868_ & ~new_n50160_;
  assign new_n50162_ = ~new_n50158_ & new_n50161_;
  assign new_n50163_ = ~new_n49868_ & ~new_n50162_;
  assign new_n50164_ = \b[23]  & ~new_n49857_;
  assign new_n50165_ = ~new_n49851_ & new_n50164_;
  assign new_n50166_ = ~new_n49859_ & ~new_n50165_;
  assign new_n50167_ = ~new_n50163_ & new_n50166_;
  assign new_n50168_ = ~new_n49859_ & ~new_n50167_;
  assign new_n50169_ = \b[24]  & ~new_n49848_;
  assign new_n50170_ = ~new_n49842_ & new_n50169_;
  assign new_n50171_ = ~new_n49850_ & ~new_n50170_;
  assign new_n50172_ = ~new_n50168_ & new_n50171_;
  assign new_n50173_ = ~new_n49850_ & ~new_n50172_;
  assign new_n50174_ = \b[25]  & ~new_n49839_;
  assign new_n50175_ = ~new_n49833_ & new_n50174_;
  assign new_n50176_ = ~new_n49841_ & ~new_n50175_;
  assign new_n50177_ = ~new_n50173_ & new_n50176_;
  assign new_n50178_ = ~new_n49841_ & ~new_n50177_;
  assign new_n50179_ = \b[26]  & ~new_n49830_;
  assign new_n50180_ = ~new_n49824_ & new_n50179_;
  assign new_n50181_ = ~new_n49832_ & ~new_n50180_;
  assign new_n50182_ = ~new_n50178_ & new_n50181_;
  assign new_n50183_ = ~new_n49832_ & ~new_n50182_;
  assign new_n50184_ = \b[27]  & ~new_n49821_;
  assign new_n50185_ = ~new_n49815_ & new_n50184_;
  assign new_n50186_ = ~new_n49823_ & ~new_n50185_;
  assign new_n50187_ = ~new_n50183_ & new_n50186_;
  assign new_n50188_ = ~new_n49823_ & ~new_n50187_;
  assign new_n50189_ = \b[28]  & ~new_n49812_;
  assign new_n50190_ = ~new_n49806_ & new_n50189_;
  assign new_n50191_ = ~new_n49814_ & ~new_n50190_;
  assign new_n50192_ = ~new_n50188_ & new_n50191_;
  assign new_n50193_ = ~new_n49814_ & ~new_n50192_;
  assign new_n50194_ = \b[29]  & ~new_n49803_;
  assign new_n50195_ = ~new_n49797_ & new_n50194_;
  assign new_n50196_ = ~new_n49805_ & ~new_n50195_;
  assign new_n50197_ = ~new_n50193_ & new_n50196_;
  assign new_n50198_ = ~new_n49805_ & ~new_n50197_;
  assign new_n50199_ = \b[30]  & ~new_n49794_;
  assign new_n50200_ = ~new_n49788_ & new_n50199_;
  assign new_n50201_ = ~new_n49796_ & ~new_n50200_;
  assign new_n50202_ = ~new_n50198_ & new_n50201_;
  assign new_n50203_ = ~new_n49796_ & ~new_n50202_;
  assign new_n50204_ = \b[31]  & ~new_n49785_;
  assign new_n50205_ = ~new_n49779_ & new_n50204_;
  assign new_n50206_ = ~new_n49787_ & ~new_n50205_;
  assign new_n50207_ = ~new_n50203_ & new_n50206_;
  assign new_n50208_ = ~new_n49787_ & ~new_n50207_;
  assign new_n50209_ = \b[32]  & ~new_n49776_;
  assign new_n50210_ = ~new_n49770_ & new_n50209_;
  assign new_n50211_ = ~new_n49778_ & ~new_n50210_;
  assign new_n50212_ = ~new_n50208_ & new_n50211_;
  assign new_n50213_ = ~new_n49778_ & ~new_n50212_;
  assign new_n50214_ = \b[33]  & ~new_n49767_;
  assign new_n50215_ = ~new_n49761_ & new_n50214_;
  assign new_n50216_ = ~new_n49769_ & ~new_n50215_;
  assign new_n50217_ = ~new_n50213_ & new_n50216_;
  assign new_n50218_ = ~new_n49769_ & ~new_n50217_;
  assign new_n50219_ = \b[34]  & ~new_n49758_;
  assign new_n50220_ = ~new_n49752_ & new_n50219_;
  assign new_n50221_ = ~new_n49760_ & ~new_n50220_;
  assign new_n50222_ = ~new_n50218_ & new_n50221_;
  assign new_n50223_ = ~new_n49760_ & ~new_n50222_;
  assign new_n50224_ = \b[35]  & ~new_n49749_;
  assign new_n50225_ = ~new_n49743_ & new_n50224_;
  assign new_n50226_ = ~new_n49751_ & ~new_n50225_;
  assign new_n50227_ = ~new_n50223_ & new_n50226_;
  assign new_n50228_ = ~new_n49751_ & ~new_n50227_;
  assign new_n50229_ = \b[36]  & ~new_n49740_;
  assign new_n50230_ = ~new_n49734_ & new_n50229_;
  assign new_n50231_ = ~new_n49742_ & ~new_n50230_;
  assign new_n50232_ = ~new_n50228_ & new_n50231_;
  assign new_n50233_ = ~new_n49742_ & ~new_n50232_;
  assign new_n50234_ = \b[37]  & ~new_n49731_;
  assign new_n50235_ = ~new_n49725_ & new_n50234_;
  assign new_n50236_ = ~new_n49733_ & ~new_n50235_;
  assign new_n50237_ = ~new_n50233_ & new_n50236_;
  assign new_n50238_ = ~new_n49733_ & ~new_n50237_;
  assign new_n50239_ = \b[38]  & ~new_n49722_;
  assign new_n50240_ = ~new_n49716_ & new_n50239_;
  assign new_n50241_ = ~new_n49724_ & ~new_n50240_;
  assign new_n50242_ = ~new_n50238_ & new_n50241_;
  assign new_n50243_ = ~new_n49724_ & ~new_n50242_;
  assign new_n50244_ = \b[39]  & ~new_n49713_;
  assign new_n50245_ = ~new_n49707_ & new_n50244_;
  assign new_n50246_ = ~new_n49715_ & ~new_n50245_;
  assign new_n50247_ = ~new_n50243_ & new_n50246_;
  assign new_n50248_ = ~new_n49715_ & ~new_n50247_;
  assign new_n50249_ = \b[40]  & ~new_n49704_;
  assign new_n50250_ = ~new_n49698_ & new_n50249_;
  assign new_n50251_ = ~new_n49706_ & ~new_n50250_;
  assign new_n50252_ = ~new_n50248_ & new_n50251_;
  assign new_n50253_ = ~new_n49706_ & ~new_n50252_;
  assign new_n50254_ = \b[41]  & ~new_n49695_;
  assign new_n50255_ = ~new_n49689_ & new_n50254_;
  assign new_n50256_ = ~new_n49697_ & ~new_n50255_;
  assign new_n50257_ = ~new_n50253_ & new_n50256_;
  assign new_n50258_ = ~new_n49697_ & ~new_n50257_;
  assign new_n50259_ = \b[42]  & ~new_n49686_;
  assign new_n50260_ = ~new_n49680_ & new_n50259_;
  assign new_n50261_ = ~new_n49688_ & ~new_n50260_;
  assign new_n50262_ = ~new_n50258_ & new_n50261_;
  assign new_n50263_ = ~new_n49688_ & ~new_n50262_;
  assign new_n50264_ = \b[43]  & ~new_n49677_;
  assign new_n50265_ = ~new_n49671_ & new_n50264_;
  assign new_n50266_ = ~new_n49679_ & ~new_n50265_;
  assign new_n50267_ = ~new_n50263_ & new_n50266_;
  assign new_n50268_ = ~new_n49679_ & ~new_n50267_;
  assign new_n50269_ = \b[44]  & ~new_n49668_;
  assign new_n50270_ = ~new_n49662_ & new_n50269_;
  assign new_n50271_ = ~new_n49670_ & ~new_n50270_;
  assign new_n50272_ = ~new_n50268_ & new_n50271_;
  assign new_n50273_ = ~new_n49670_ & ~new_n50272_;
  assign new_n50274_ = \b[45]  & ~new_n49659_;
  assign new_n50275_ = ~new_n49653_ & new_n50274_;
  assign new_n50276_ = ~new_n49661_ & ~new_n50275_;
  assign new_n50277_ = ~new_n50273_ & new_n50276_;
  assign new_n50278_ = ~new_n49661_ & ~new_n50277_;
  assign new_n50279_ = \b[46]  & ~new_n49650_;
  assign new_n50280_ = ~new_n49644_ & new_n50279_;
  assign new_n50281_ = ~new_n49652_ & ~new_n50280_;
  assign new_n50282_ = ~new_n50278_ & new_n50281_;
  assign new_n50283_ = ~new_n49652_ & ~new_n50282_;
  assign new_n50284_ = \b[47]  & ~new_n49641_;
  assign new_n50285_ = ~new_n49635_ & new_n50284_;
  assign new_n50286_ = ~new_n49643_ & ~new_n50285_;
  assign new_n50287_ = ~new_n50283_ & new_n50286_;
  assign new_n50288_ = ~new_n49643_ & ~new_n50287_;
  assign new_n50289_ = \b[48]  & ~new_n49632_;
  assign new_n50290_ = ~new_n49626_ & new_n50289_;
  assign new_n50291_ = ~new_n49634_ & ~new_n50290_;
  assign new_n50292_ = ~new_n50288_ & new_n50291_;
  assign new_n50293_ = ~new_n49634_ & ~new_n50292_;
  assign new_n50294_ = \b[49]  & ~new_n49623_;
  assign new_n50295_ = ~new_n49617_ & new_n50294_;
  assign new_n50296_ = ~new_n49625_ & ~new_n50295_;
  assign new_n50297_ = ~new_n50293_ & new_n50296_;
  assign new_n50298_ = ~new_n49625_ & ~new_n50297_;
  assign new_n50299_ = \b[50]  & ~new_n49614_;
  assign new_n50300_ = ~new_n49608_ & new_n50299_;
  assign new_n50301_ = ~new_n49616_ & ~new_n50300_;
  assign new_n50302_ = ~new_n50298_ & new_n50301_;
  assign new_n50303_ = ~new_n49616_ & ~new_n50302_;
  assign new_n50304_ = \b[51]  & ~new_n49605_;
  assign new_n50305_ = ~new_n49599_ & new_n50304_;
  assign new_n50306_ = ~new_n49607_ & ~new_n50305_;
  assign new_n50307_ = ~new_n50303_ & new_n50306_;
  assign new_n50308_ = ~new_n49607_ & ~new_n50307_;
  assign new_n50309_ = \b[52]  & ~new_n49596_;
  assign new_n50310_ = ~new_n49590_ & new_n50309_;
  assign new_n50311_ = ~new_n49598_ & ~new_n50310_;
  assign new_n50312_ = ~new_n50308_ & new_n50311_;
  assign new_n50313_ = ~new_n49598_ & ~new_n50312_;
  assign new_n50314_ = \b[53]  & ~new_n49587_;
  assign new_n50315_ = ~new_n49581_ & new_n50314_;
  assign new_n50316_ = ~new_n49589_ & ~new_n50315_;
  assign new_n50317_ = ~new_n50313_ & new_n50316_;
  assign new_n50318_ = ~new_n49589_ & ~new_n50317_;
  assign new_n50319_ = \b[54]  & ~new_n49578_;
  assign new_n50320_ = ~new_n49572_ & new_n50319_;
  assign new_n50321_ = ~new_n49580_ & ~new_n50320_;
  assign new_n50322_ = ~new_n50318_ & new_n50321_;
  assign new_n50323_ = ~new_n49580_ & ~new_n50322_;
  assign new_n50324_ = ~new_n48834_ & ~new_n49571_;
  assign new_n50325_ = ~new_n48836_ & new_n49568_;
  assign new_n50326_ = ~new_n49564_ & new_n50325_;
  assign new_n50327_ = ~new_n49565_ & ~new_n49568_;
  assign new_n50328_ = ~new_n50326_ & ~new_n50327_;
  assign new_n50329_ = new_n49571_ & ~new_n50328_;
  assign new_n50330_ = ~new_n50324_ & ~new_n50329_;
  assign new_n50331_ = ~\b[55]  & ~new_n50330_;
  assign new_n50332_ = \b[55]  & ~new_n50324_;
  assign new_n50333_ = ~new_n50329_ & new_n50332_;
  assign new_n50334_ = new_n337_ & ~new_n50333_;
  assign new_n50335_ = ~new_n50331_ & new_n50334_;
  assign new_n50336_ = ~new_n50323_ & new_n50335_;
  assign new_n50337_ = new_n21537_ & ~new_n50330_;
  assign new_n50338_ = ~new_n50336_ & ~new_n50337_;
  assign new_n50339_ = ~new_n49589_ & new_n50321_;
  assign new_n50340_ = ~new_n50317_ & new_n50339_;
  assign new_n50341_ = ~new_n50318_ & ~new_n50321_;
  assign new_n50342_ = ~new_n50340_ & ~new_n50341_;
  assign new_n50343_ = ~new_n50338_ & ~new_n50342_;
  assign new_n50344_ = ~new_n49579_ & ~new_n50337_;
  assign new_n50345_ = ~new_n50336_ & new_n50344_;
  assign new_n50346_ = ~new_n50343_ & ~new_n50345_;
  assign new_n50347_ = ~\b[55]  & ~new_n50346_;
  assign new_n50348_ = ~new_n49598_ & new_n50316_;
  assign new_n50349_ = ~new_n50312_ & new_n50348_;
  assign new_n50350_ = ~new_n50313_ & ~new_n50316_;
  assign new_n50351_ = ~new_n50349_ & ~new_n50350_;
  assign new_n50352_ = ~new_n50338_ & ~new_n50351_;
  assign new_n50353_ = ~new_n49588_ & ~new_n50337_;
  assign new_n50354_ = ~new_n50336_ & new_n50353_;
  assign new_n50355_ = ~new_n50352_ & ~new_n50354_;
  assign new_n50356_ = ~\b[54]  & ~new_n50355_;
  assign new_n50357_ = ~new_n49607_ & new_n50311_;
  assign new_n50358_ = ~new_n50307_ & new_n50357_;
  assign new_n50359_ = ~new_n50308_ & ~new_n50311_;
  assign new_n50360_ = ~new_n50358_ & ~new_n50359_;
  assign new_n50361_ = ~new_n50338_ & ~new_n50360_;
  assign new_n50362_ = ~new_n49597_ & ~new_n50337_;
  assign new_n50363_ = ~new_n50336_ & new_n50362_;
  assign new_n50364_ = ~new_n50361_ & ~new_n50363_;
  assign new_n50365_ = ~\b[53]  & ~new_n50364_;
  assign new_n50366_ = ~new_n49616_ & new_n50306_;
  assign new_n50367_ = ~new_n50302_ & new_n50366_;
  assign new_n50368_ = ~new_n50303_ & ~new_n50306_;
  assign new_n50369_ = ~new_n50367_ & ~new_n50368_;
  assign new_n50370_ = ~new_n50338_ & ~new_n50369_;
  assign new_n50371_ = ~new_n49606_ & ~new_n50337_;
  assign new_n50372_ = ~new_n50336_ & new_n50371_;
  assign new_n50373_ = ~new_n50370_ & ~new_n50372_;
  assign new_n50374_ = ~\b[52]  & ~new_n50373_;
  assign new_n50375_ = ~new_n49625_ & new_n50301_;
  assign new_n50376_ = ~new_n50297_ & new_n50375_;
  assign new_n50377_ = ~new_n50298_ & ~new_n50301_;
  assign new_n50378_ = ~new_n50376_ & ~new_n50377_;
  assign new_n50379_ = ~new_n50338_ & ~new_n50378_;
  assign new_n50380_ = ~new_n49615_ & ~new_n50337_;
  assign new_n50381_ = ~new_n50336_ & new_n50380_;
  assign new_n50382_ = ~new_n50379_ & ~new_n50381_;
  assign new_n50383_ = ~\b[51]  & ~new_n50382_;
  assign new_n50384_ = ~new_n49634_ & new_n50296_;
  assign new_n50385_ = ~new_n50292_ & new_n50384_;
  assign new_n50386_ = ~new_n50293_ & ~new_n50296_;
  assign new_n50387_ = ~new_n50385_ & ~new_n50386_;
  assign new_n50388_ = ~new_n50338_ & ~new_n50387_;
  assign new_n50389_ = ~new_n49624_ & ~new_n50337_;
  assign new_n50390_ = ~new_n50336_ & new_n50389_;
  assign new_n50391_ = ~new_n50388_ & ~new_n50390_;
  assign new_n50392_ = ~\b[50]  & ~new_n50391_;
  assign new_n50393_ = ~new_n49643_ & new_n50291_;
  assign new_n50394_ = ~new_n50287_ & new_n50393_;
  assign new_n50395_ = ~new_n50288_ & ~new_n50291_;
  assign new_n50396_ = ~new_n50394_ & ~new_n50395_;
  assign new_n50397_ = ~new_n50338_ & ~new_n50396_;
  assign new_n50398_ = ~new_n49633_ & ~new_n50337_;
  assign new_n50399_ = ~new_n50336_ & new_n50398_;
  assign new_n50400_ = ~new_n50397_ & ~new_n50399_;
  assign new_n50401_ = ~\b[49]  & ~new_n50400_;
  assign new_n50402_ = ~new_n49652_ & new_n50286_;
  assign new_n50403_ = ~new_n50282_ & new_n50402_;
  assign new_n50404_ = ~new_n50283_ & ~new_n50286_;
  assign new_n50405_ = ~new_n50403_ & ~new_n50404_;
  assign new_n50406_ = ~new_n50338_ & ~new_n50405_;
  assign new_n50407_ = ~new_n49642_ & ~new_n50337_;
  assign new_n50408_ = ~new_n50336_ & new_n50407_;
  assign new_n50409_ = ~new_n50406_ & ~new_n50408_;
  assign new_n50410_ = ~\b[48]  & ~new_n50409_;
  assign new_n50411_ = ~new_n49661_ & new_n50281_;
  assign new_n50412_ = ~new_n50277_ & new_n50411_;
  assign new_n50413_ = ~new_n50278_ & ~new_n50281_;
  assign new_n50414_ = ~new_n50412_ & ~new_n50413_;
  assign new_n50415_ = ~new_n50338_ & ~new_n50414_;
  assign new_n50416_ = ~new_n49651_ & ~new_n50337_;
  assign new_n50417_ = ~new_n50336_ & new_n50416_;
  assign new_n50418_ = ~new_n50415_ & ~new_n50417_;
  assign new_n50419_ = ~\b[47]  & ~new_n50418_;
  assign new_n50420_ = ~new_n49670_ & new_n50276_;
  assign new_n50421_ = ~new_n50272_ & new_n50420_;
  assign new_n50422_ = ~new_n50273_ & ~new_n50276_;
  assign new_n50423_ = ~new_n50421_ & ~new_n50422_;
  assign new_n50424_ = ~new_n50338_ & ~new_n50423_;
  assign new_n50425_ = ~new_n49660_ & ~new_n50337_;
  assign new_n50426_ = ~new_n50336_ & new_n50425_;
  assign new_n50427_ = ~new_n50424_ & ~new_n50426_;
  assign new_n50428_ = ~\b[46]  & ~new_n50427_;
  assign new_n50429_ = ~new_n49679_ & new_n50271_;
  assign new_n50430_ = ~new_n50267_ & new_n50429_;
  assign new_n50431_ = ~new_n50268_ & ~new_n50271_;
  assign new_n50432_ = ~new_n50430_ & ~new_n50431_;
  assign new_n50433_ = ~new_n50338_ & ~new_n50432_;
  assign new_n50434_ = ~new_n49669_ & ~new_n50337_;
  assign new_n50435_ = ~new_n50336_ & new_n50434_;
  assign new_n50436_ = ~new_n50433_ & ~new_n50435_;
  assign new_n50437_ = ~\b[45]  & ~new_n50436_;
  assign new_n50438_ = ~new_n49688_ & new_n50266_;
  assign new_n50439_ = ~new_n50262_ & new_n50438_;
  assign new_n50440_ = ~new_n50263_ & ~new_n50266_;
  assign new_n50441_ = ~new_n50439_ & ~new_n50440_;
  assign new_n50442_ = ~new_n50338_ & ~new_n50441_;
  assign new_n50443_ = ~new_n49678_ & ~new_n50337_;
  assign new_n50444_ = ~new_n50336_ & new_n50443_;
  assign new_n50445_ = ~new_n50442_ & ~new_n50444_;
  assign new_n50446_ = ~\b[44]  & ~new_n50445_;
  assign new_n50447_ = ~new_n49697_ & new_n50261_;
  assign new_n50448_ = ~new_n50257_ & new_n50447_;
  assign new_n50449_ = ~new_n50258_ & ~new_n50261_;
  assign new_n50450_ = ~new_n50448_ & ~new_n50449_;
  assign new_n50451_ = ~new_n50338_ & ~new_n50450_;
  assign new_n50452_ = ~new_n49687_ & ~new_n50337_;
  assign new_n50453_ = ~new_n50336_ & new_n50452_;
  assign new_n50454_ = ~new_n50451_ & ~new_n50453_;
  assign new_n50455_ = ~\b[43]  & ~new_n50454_;
  assign new_n50456_ = ~new_n49706_ & new_n50256_;
  assign new_n50457_ = ~new_n50252_ & new_n50456_;
  assign new_n50458_ = ~new_n50253_ & ~new_n50256_;
  assign new_n50459_ = ~new_n50457_ & ~new_n50458_;
  assign new_n50460_ = ~new_n50338_ & ~new_n50459_;
  assign new_n50461_ = ~new_n49696_ & ~new_n50337_;
  assign new_n50462_ = ~new_n50336_ & new_n50461_;
  assign new_n50463_ = ~new_n50460_ & ~new_n50462_;
  assign new_n50464_ = ~\b[42]  & ~new_n50463_;
  assign new_n50465_ = ~new_n49715_ & new_n50251_;
  assign new_n50466_ = ~new_n50247_ & new_n50465_;
  assign new_n50467_ = ~new_n50248_ & ~new_n50251_;
  assign new_n50468_ = ~new_n50466_ & ~new_n50467_;
  assign new_n50469_ = ~new_n50338_ & ~new_n50468_;
  assign new_n50470_ = ~new_n49705_ & ~new_n50337_;
  assign new_n50471_ = ~new_n50336_ & new_n50470_;
  assign new_n50472_ = ~new_n50469_ & ~new_n50471_;
  assign new_n50473_ = ~\b[41]  & ~new_n50472_;
  assign new_n50474_ = ~new_n49724_ & new_n50246_;
  assign new_n50475_ = ~new_n50242_ & new_n50474_;
  assign new_n50476_ = ~new_n50243_ & ~new_n50246_;
  assign new_n50477_ = ~new_n50475_ & ~new_n50476_;
  assign new_n50478_ = ~new_n50338_ & ~new_n50477_;
  assign new_n50479_ = ~new_n49714_ & ~new_n50337_;
  assign new_n50480_ = ~new_n50336_ & new_n50479_;
  assign new_n50481_ = ~new_n50478_ & ~new_n50480_;
  assign new_n50482_ = ~\b[40]  & ~new_n50481_;
  assign new_n50483_ = ~new_n49733_ & new_n50241_;
  assign new_n50484_ = ~new_n50237_ & new_n50483_;
  assign new_n50485_ = ~new_n50238_ & ~new_n50241_;
  assign new_n50486_ = ~new_n50484_ & ~new_n50485_;
  assign new_n50487_ = ~new_n50338_ & ~new_n50486_;
  assign new_n50488_ = ~new_n49723_ & ~new_n50337_;
  assign new_n50489_ = ~new_n50336_ & new_n50488_;
  assign new_n50490_ = ~new_n50487_ & ~new_n50489_;
  assign new_n50491_ = ~\b[39]  & ~new_n50490_;
  assign new_n50492_ = ~new_n49742_ & new_n50236_;
  assign new_n50493_ = ~new_n50232_ & new_n50492_;
  assign new_n50494_ = ~new_n50233_ & ~new_n50236_;
  assign new_n50495_ = ~new_n50493_ & ~new_n50494_;
  assign new_n50496_ = ~new_n50338_ & ~new_n50495_;
  assign new_n50497_ = ~new_n49732_ & ~new_n50337_;
  assign new_n50498_ = ~new_n50336_ & new_n50497_;
  assign new_n50499_ = ~new_n50496_ & ~new_n50498_;
  assign new_n50500_ = ~\b[38]  & ~new_n50499_;
  assign new_n50501_ = ~new_n49751_ & new_n50231_;
  assign new_n50502_ = ~new_n50227_ & new_n50501_;
  assign new_n50503_ = ~new_n50228_ & ~new_n50231_;
  assign new_n50504_ = ~new_n50502_ & ~new_n50503_;
  assign new_n50505_ = ~new_n50338_ & ~new_n50504_;
  assign new_n50506_ = ~new_n49741_ & ~new_n50337_;
  assign new_n50507_ = ~new_n50336_ & new_n50506_;
  assign new_n50508_ = ~new_n50505_ & ~new_n50507_;
  assign new_n50509_ = ~\b[37]  & ~new_n50508_;
  assign new_n50510_ = ~new_n49760_ & new_n50226_;
  assign new_n50511_ = ~new_n50222_ & new_n50510_;
  assign new_n50512_ = ~new_n50223_ & ~new_n50226_;
  assign new_n50513_ = ~new_n50511_ & ~new_n50512_;
  assign new_n50514_ = ~new_n50338_ & ~new_n50513_;
  assign new_n50515_ = ~new_n49750_ & ~new_n50337_;
  assign new_n50516_ = ~new_n50336_ & new_n50515_;
  assign new_n50517_ = ~new_n50514_ & ~new_n50516_;
  assign new_n50518_ = ~\b[36]  & ~new_n50517_;
  assign new_n50519_ = ~new_n49769_ & new_n50221_;
  assign new_n50520_ = ~new_n50217_ & new_n50519_;
  assign new_n50521_ = ~new_n50218_ & ~new_n50221_;
  assign new_n50522_ = ~new_n50520_ & ~new_n50521_;
  assign new_n50523_ = ~new_n50338_ & ~new_n50522_;
  assign new_n50524_ = ~new_n49759_ & ~new_n50337_;
  assign new_n50525_ = ~new_n50336_ & new_n50524_;
  assign new_n50526_ = ~new_n50523_ & ~new_n50525_;
  assign new_n50527_ = ~\b[35]  & ~new_n50526_;
  assign new_n50528_ = ~new_n49778_ & new_n50216_;
  assign new_n50529_ = ~new_n50212_ & new_n50528_;
  assign new_n50530_ = ~new_n50213_ & ~new_n50216_;
  assign new_n50531_ = ~new_n50529_ & ~new_n50530_;
  assign new_n50532_ = ~new_n50338_ & ~new_n50531_;
  assign new_n50533_ = ~new_n49768_ & ~new_n50337_;
  assign new_n50534_ = ~new_n50336_ & new_n50533_;
  assign new_n50535_ = ~new_n50532_ & ~new_n50534_;
  assign new_n50536_ = ~\b[34]  & ~new_n50535_;
  assign new_n50537_ = ~new_n49787_ & new_n50211_;
  assign new_n50538_ = ~new_n50207_ & new_n50537_;
  assign new_n50539_ = ~new_n50208_ & ~new_n50211_;
  assign new_n50540_ = ~new_n50538_ & ~new_n50539_;
  assign new_n50541_ = ~new_n50338_ & ~new_n50540_;
  assign new_n50542_ = ~new_n49777_ & ~new_n50337_;
  assign new_n50543_ = ~new_n50336_ & new_n50542_;
  assign new_n50544_ = ~new_n50541_ & ~new_n50543_;
  assign new_n50545_ = ~\b[33]  & ~new_n50544_;
  assign new_n50546_ = ~new_n49796_ & new_n50206_;
  assign new_n50547_ = ~new_n50202_ & new_n50546_;
  assign new_n50548_ = ~new_n50203_ & ~new_n50206_;
  assign new_n50549_ = ~new_n50547_ & ~new_n50548_;
  assign new_n50550_ = ~new_n50338_ & ~new_n50549_;
  assign new_n50551_ = ~new_n49786_ & ~new_n50337_;
  assign new_n50552_ = ~new_n50336_ & new_n50551_;
  assign new_n50553_ = ~new_n50550_ & ~new_n50552_;
  assign new_n50554_ = ~\b[32]  & ~new_n50553_;
  assign new_n50555_ = ~new_n49805_ & new_n50201_;
  assign new_n50556_ = ~new_n50197_ & new_n50555_;
  assign new_n50557_ = ~new_n50198_ & ~new_n50201_;
  assign new_n50558_ = ~new_n50556_ & ~new_n50557_;
  assign new_n50559_ = ~new_n50338_ & ~new_n50558_;
  assign new_n50560_ = ~new_n49795_ & ~new_n50337_;
  assign new_n50561_ = ~new_n50336_ & new_n50560_;
  assign new_n50562_ = ~new_n50559_ & ~new_n50561_;
  assign new_n50563_ = ~\b[31]  & ~new_n50562_;
  assign new_n50564_ = ~new_n49814_ & new_n50196_;
  assign new_n50565_ = ~new_n50192_ & new_n50564_;
  assign new_n50566_ = ~new_n50193_ & ~new_n50196_;
  assign new_n50567_ = ~new_n50565_ & ~new_n50566_;
  assign new_n50568_ = ~new_n50338_ & ~new_n50567_;
  assign new_n50569_ = ~new_n49804_ & ~new_n50337_;
  assign new_n50570_ = ~new_n50336_ & new_n50569_;
  assign new_n50571_ = ~new_n50568_ & ~new_n50570_;
  assign new_n50572_ = ~\b[30]  & ~new_n50571_;
  assign new_n50573_ = ~new_n49823_ & new_n50191_;
  assign new_n50574_ = ~new_n50187_ & new_n50573_;
  assign new_n50575_ = ~new_n50188_ & ~new_n50191_;
  assign new_n50576_ = ~new_n50574_ & ~new_n50575_;
  assign new_n50577_ = ~new_n50338_ & ~new_n50576_;
  assign new_n50578_ = ~new_n49813_ & ~new_n50337_;
  assign new_n50579_ = ~new_n50336_ & new_n50578_;
  assign new_n50580_ = ~new_n50577_ & ~new_n50579_;
  assign new_n50581_ = ~\b[29]  & ~new_n50580_;
  assign new_n50582_ = ~new_n49832_ & new_n50186_;
  assign new_n50583_ = ~new_n50182_ & new_n50582_;
  assign new_n50584_ = ~new_n50183_ & ~new_n50186_;
  assign new_n50585_ = ~new_n50583_ & ~new_n50584_;
  assign new_n50586_ = ~new_n50338_ & ~new_n50585_;
  assign new_n50587_ = ~new_n49822_ & ~new_n50337_;
  assign new_n50588_ = ~new_n50336_ & new_n50587_;
  assign new_n50589_ = ~new_n50586_ & ~new_n50588_;
  assign new_n50590_ = ~\b[28]  & ~new_n50589_;
  assign new_n50591_ = ~new_n49841_ & new_n50181_;
  assign new_n50592_ = ~new_n50177_ & new_n50591_;
  assign new_n50593_ = ~new_n50178_ & ~new_n50181_;
  assign new_n50594_ = ~new_n50592_ & ~new_n50593_;
  assign new_n50595_ = ~new_n50338_ & ~new_n50594_;
  assign new_n50596_ = ~new_n49831_ & ~new_n50337_;
  assign new_n50597_ = ~new_n50336_ & new_n50596_;
  assign new_n50598_ = ~new_n50595_ & ~new_n50597_;
  assign new_n50599_ = ~\b[27]  & ~new_n50598_;
  assign new_n50600_ = ~new_n49850_ & new_n50176_;
  assign new_n50601_ = ~new_n50172_ & new_n50600_;
  assign new_n50602_ = ~new_n50173_ & ~new_n50176_;
  assign new_n50603_ = ~new_n50601_ & ~new_n50602_;
  assign new_n50604_ = ~new_n50338_ & ~new_n50603_;
  assign new_n50605_ = ~new_n49840_ & ~new_n50337_;
  assign new_n50606_ = ~new_n50336_ & new_n50605_;
  assign new_n50607_ = ~new_n50604_ & ~new_n50606_;
  assign new_n50608_ = ~\b[26]  & ~new_n50607_;
  assign new_n50609_ = ~new_n49859_ & new_n50171_;
  assign new_n50610_ = ~new_n50167_ & new_n50609_;
  assign new_n50611_ = ~new_n50168_ & ~new_n50171_;
  assign new_n50612_ = ~new_n50610_ & ~new_n50611_;
  assign new_n50613_ = ~new_n50338_ & ~new_n50612_;
  assign new_n50614_ = ~new_n49849_ & ~new_n50337_;
  assign new_n50615_ = ~new_n50336_ & new_n50614_;
  assign new_n50616_ = ~new_n50613_ & ~new_n50615_;
  assign new_n50617_ = ~\b[25]  & ~new_n50616_;
  assign new_n50618_ = ~new_n49868_ & new_n50166_;
  assign new_n50619_ = ~new_n50162_ & new_n50618_;
  assign new_n50620_ = ~new_n50163_ & ~new_n50166_;
  assign new_n50621_ = ~new_n50619_ & ~new_n50620_;
  assign new_n50622_ = ~new_n50338_ & ~new_n50621_;
  assign new_n50623_ = ~new_n49858_ & ~new_n50337_;
  assign new_n50624_ = ~new_n50336_ & new_n50623_;
  assign new_n50625_ = ~new_n50622_ & ~new_n50624_;
  assign new_n50626_ = ~\b[24]  & ~new_n50625_;
  assign new_n50627_ = ~new_n49877_ & new_n50161_;
  assign new_n50628_ = ~new_n50157_ & new_n50627_;
  assign new_n50629_ = ~new_n50158_ & ~new_n50161_;
  assign new_n50630_ = ~new_n50628_ & ~new_n50629_;
  assign new_n50631_ = ~new_n50338_ & ~new_n50630_;
  assign new_n50632_ = ~new_n49867_ & ~new_n50337_;
  assign new_n50633_ = ~new_n50336_ & new_n50632_;
  assign new_n50634_ = ~new_n50631_ & ~new_n50633_;
  assign new_n50635_ = ~\b[23]  & ~new_n50634_;
  assign new_n50636_ = ~new_n49886_ & new_n50156_;
  assign new_n50637_ = ~new_n50152_ & new_n50636_;
  assign new_n50638_ = ~new_n50153_ & ~new_n50156_;
  assign new_n50639_ = ~new_n50637_ & ~new_n50638_;
  assign new_n50640_ = ~new_n50338_ & ~new_n50639_;
  assign new_n50641_ = ~new_n49876_ & ~new_n50337_;
  assign new_n50642_ = ~new_n50336_ & new_n50641_;
  assign new_n50643_ = ~new_n50640_ & ~new_n50642_;
  assign new_n50644_ = ~\b[22]  & ~new_n50643_;
  assign new_n50645_ = ~new_n49895_ & new_n50151_;
  assign new_n50646_ = ~new_n50147_ & new_n50645_;
  assign new_n50647_ = ~new_n50148_ & ~new_n50151_;
  assign new_n50648_ = ~new_n50646_ & ~new_n50647_;
  assign new_n50649_ = ~new_n50338_ & ~new_n50648_;
  assign new_n50650_ = ~new_n49885_ & ~new_n50337_;
  assign new_n50651_ = ~new_n50336_ & new_n50650_;
  assign new_n50652_ = ~new_n50649_ & ~new_n50651_;
  assign new_n50653_ = ~\b[21]  & ~new_n50652_;
  assign new_n50654_ = ~new_n49904_ & new_n50146_;
  assign new_n50655_ = ~new_n50142_ & new_n50654_;
  assign new_n50656_ = ~new_n50143_ & ~new_n50146_;
  assign new_n50657_ = ~new_n50655_ & ~new_n50656_;
  assign new_n50658_ = ~new_n50338_ & ~new_n50657_;
  assign new_n50659_ = ~new_n49894_ & ~new_n50337_;
  assign new_n50660_ = ~new_n50336_ & new_n50659_;
  assign new_n50661_ = ~new_n50658_ & ~new_n50660_;
  assign new_n50662_ = ~\b[20]  & ~new_n50661_;
  assign new_n50663_ = ~new_n49913_ & new_n50141_;
  assign new_n50664_ = ~new_n50137_ & new_n50663_;
  assign new_n50665_ = ~new_n50138_ & ~new_n50141_;
  assign new_n50666_ = ~new_n50664_ & ~new_n50665_;
  assign new_n50667_ = ~new_n50338_ & ~new_n50666_;
  assign new_n50668_ = ~new_n49903_ & ~new_n50337_;
  assign new_n50669_ = ~new_n50336_ & new_n50668_;
  assign new_n50670_ = ~new_n50667_ & ~new_n50669_;
  assign new_n50671_ = ~\b[19]  & ~new_n50670_;
  assign new_n50672_ = ~new_n49922_ & new_n50136_;
  assign new_n50673_ = ~new_n50132_ & new_n50672_;
  assign new_n50674_ = ~new_n50133_ & ~new_n50136_;
  assign new_n50675_ = ~new_n50673_ & ~new_n50674_;
  assign new_n50676_ = ~new_n50338_ & ~new_n50675_;
  assign new_n50677_ = ~new_n49912_ & ~new_n50337_;
  assign new_n50678_ = ~new_n50336_ & new_n50677_;
  assign new_n50679_ = ~new_n50676_ & ~new_n50678_;
  assign new_n50680_ = ~\b[18]  & ~new_n50679_;
  assign new_n50681_ = ~new_n49931_ & new_n50131_;
  assign new_n50682_ = ~new_n50127_ & new_n50681_;
  assign new_n50683_ = ~new_n50128_ & ~new_n50131_;
  assign new_n50684_ = ~new_n50682_ & ~new_n50683_;
  assign new_n50685_ = ~new_n50338_ & ~new_n50684_;
  assign new_n50686_ = ~new_n49921_ & ~new_n50337_;
  assign new_n50687_ = ~new_n50336_ & new_n50686_;
  assign new_n50688_ = ~new_n50685_ & ~new_n50687_;
  assign new_n50689_ = ~\b[17]  & ~new_n50688_;
  assign new_n50690_ = ~new_n49940_ & new_n50126_;
  assign new_n50691_ = ~new_n50122_ & new_n50690_;
  assign new_n50692_ = ~new_n50123_ & ~new_n50126_;
  assign new_n50693_ = ~new_n50691_ & ~new_n50692_;
  assign new_n50694_ = ~new_n50338_ & ~new_n50693_;
  assign new_n50695_ = ~new_n49930_ & ~new_n50337_;
  assign new_n50696_ = ~new_n50336_ & new_n50695_;
  assign new_n50697_ = ~new_n50694_ & ~new_n50696_;
  assign new_n50698_ = ~\b[16]  & ~new_n50697_;
  assign new_n50699_ = ~new_n49949_ & new_n50121_;
  assign new_n50700_ = ~new_n50117_ & new_n50699_;
  assign new_n50701_ = ~new_n50118_ & ~new_n50121_;
  assign new_n50702_ = ~new_n50700_ & ~new_n50701_;
  assign new_n50703_ = ~new_n50338_ & ~new_n50702_;
  assign new_n50704_ = ~new_n49939_ & ~new_n50337_;
  assign new_n50705_ = ~new_n50336_ & new_n50704_;
  assign new_n50706_ = ~new_n50703_ & ~new_n50705_;
  assign new_n50707_ = ~\b[15]  & ~new_n50706_;
  assign new_n50708_ = ~new_n49958_ & new_n50116_;
  assign new_n50709_ = ~new_n50112_ & new_n50708_;
  assign new_n50710_ = ~new_n50113_ & ~new_n50116_;
  assign new_n50711_ = ~new_n50709_ & ~new_n50710_;
  assign new_n50712_ = ~new_n50338_ & ~new_n50711_;
  assign new_n50713_ = ~new_n49948_ & ~new_n50337_;
  assign new_n50714_ = ~new_n50336_ & new_n50713_;
  assign new_n50715_ = ~new_n50712_ & ~new_n50714_;
  assign new_n50716_ = ~\b[14]  & ~new_n50715_;
  assign new_n50717_ = ~new_n49967_ & new_n50111_;
  assign new_n50718_ = ~new_n50107_ & new_n50717_;
  assign new_n50719_ = ~new_n50108_ & ~new_n50111_;
  assign new_n50720_ = ~new_n50718_ & ~new_n50719_;
  assign new_n50721_ = ~new_n50338_ & ~new_n50720_;
  assign new_n50722_ = ~new_n49957_ & ~new_n50337_;
  assign new_n50723_ = ~new_n50336_ & new_n50722_;
  assign new_n50724_ = ~new_n50721_ & ~new_n50723_;
  assign new_n50725_ = ~\b[13]  & ~new_n50724_;
  assign new_n50726_ = ~new_n49976_ & new_n50106_;
  assign new_n50727_ = ~new_n50102_ & new_n50726_;
  assign new_n50728_ = ~new_n50103_ & ~new_n50106_;
  assign new_n50729_ = ~new_n50727_ & ~new_n50728_;
  assign new_n50730_ = ~new_n50338_ & ~new_n50729_;
  assign new_n50731_ = ~new_n49966_ & ~new_n50337_;
  assign new_n50732_ = ~new_n50336_ & new_n50731_;
  assign new_n50733_ = ~new_n50730_ & ~new_n50732_;
  assign new_n50734_ = ~\b[12]  & ~new_n50733_;
  assign new_n50735_ = ~new_n49985_ & new_n50101_;
  assign new_n50736_ = ~new_n50097_ & new_n50735_;
  assign new_n50737_ = ~new_n50098_ & ~new_n50101_;
  assign new_n50738_ = ~new_n50736_ & ~new_n50737_;
  assign new_n50739_ = ~new_n50338_ & ~new_n50738_;
  assign new_n50740_ = ~new_n49975_ & ~new_n50337_;
  assign new_n50741_ = ~new_n50336_ & new_n50740_;
  assign new_n50742_ = ~new_n50739_ & ~new_n50741_;
  assign new_n50743_ = ~\b[11]  & ~new_n50742_;
  assign new_n50744_ = ~new_n49994_ & new_n50096_;
  assign new_n50745_ = ~new_n50092_ & new_n50744_;
  assign new_n50746_ = ~new_n50093_ & ~new_n50096_;
  assign new_n50747_ = ~new_n50745_ & ~new_n50746_;
  assign new_n50748_ = ~new_n50338_ & ~new_n50747_;
  assign new_n50749_ = ~new_n49984_ & ~new_n50337_;
  assign new_n50750_ = ~new_n50336_ & new_n50749_;
  assign new_n50751_ = ~new_n50748_ & ~new_n50750_;
  assign new_n50752_ = ~\b[10]  & ~new_n50751_;
  assign new_n50753_ = ~new_n50003_ & new_n50091_;
  assign new_n50754_ = ~new_n50087_ & new_n50753_;
  assign new_n50755_ = ~new_n50088_ & ~new_n50091_;
  assign new_n50756_ = ~new_n50754_ & ~new_n50755_;
  assign new_n50757_ = ~new_n50338_ & ~new_n50756_;
  assign new_n50758_ = ~new_n49993_ & ~new_n50337_;
  assign new_n50759_ = ~new_n50336_ & new_n50758_;
  assign new_n50760_ = ~new_n50757_ & ~new_n50759_;
  assign new_n50761_ = ~\b[9]  & ~new_n50760_;
  assign new_n50762_ = ~new_n50012_ & new_n50086_;
  assign new_n50763_ = ~new_n50082_ & new_n50762_;
  assign new_n50764_ = ~new_n50083_ & ~new_n50086_;
  assign new_n50765_ = ~new_n50763_ & ~new_n50764_;
  assign new_n50766_ = ~new_n50338_ & ~new_n50765_;
  assign new_n50767_ = ~new_n50002_ & ~new_n50337_;
  assign new_n50768_ = ~new_n50336_ & new_n50767_;
  assign new_n50769_ = ~new_n50766_ & ~new_n50768_;
  assign new_n50770_ = ~\b[8]  & ~new_n50769_;
  assign new_n50771_ = ~new_n50021_ & new_n50081_;
  assign new_n50772_ = ~new_n50077_ & new_n50771_;
  assign new_n50773_ = ~new_n50078_ & ~new_n50081_;
  assign new_n50774_ = ~new_n50772_ & ~new_n50773_;
  assign new_n50775_ = ~new_n50338_ & ~new_n50774_;
  assign new_n50776_ = ~new_n50011_ & ~new_n50337_;
  assign new_n50777_ = ~new_n50336_ & new_n50776_;
  assign new_n50778_ = ~new_n50775_ & ~new_n50777_;
  assign new_n50779_ = ~\b[7]  & ~new_n50778_;
  assign new_n50780_ = ~new_n50030_ & new_n50076_;
  assign new_n50781_ = ~new_n50072_ & new_n50780_;
  assign new_n50782_ = ~new_n50073_ & ~new_n50076_;
  assign new_n50783_ = ~new_n50781_ & ~new_n50782_;
  assign new_n50784_ = ~new_n50338_ & ~new_n50783_;
  assign new_n50785_ = ~new_n50020_ & ~new_n50337_;
  assign new_n50786_ = ~new_n50336_ & new_n50785_;
  assign new_n50787_ = ~new_n50784_ & ~new_n50786_;
  assign new_n50788_ = ~\b[6]  & ~new_n50787_;
  assign new_n50789_ = ~new_n50039_ & new_n50071_;
  assign new_n50790_ = ~new_n50067_ & new_n50789_;
  assign new_n50791_ = ~new_n50068_ & ~new_n50071_;
  assign new_n50792_ = ~new_n50790_ & ~new_n50791_;
  assign new_n50793_ = ~new_n50338_ & ~new_n50792_;
  assign new_n50794_ = ~new_n50029_ & ~new_n50337_;
  assign new_n50795_ = ~new_n50336_ & new_n50794_;
  assign new_n50796_ = ~new_n50793_ & ~new_n50795_;
  assign new_n50797_ = ~\b[5]  & ~new_n50796_;
  assign new_n50798_ = ~new_n50047_ & new_n50066_;
  assign new_n50799_ = ~new_n50062_ & new_n50798_;
  assign new_n50800_ = ~new_n50063_ & ~new_n50066_;
  assign new_n50801_ = ~new_n50799_ & ~new_n50800_;
  assign new_n50802_ = ~new_n50338_ & ~new_n50801_;
  assign new_n50803_ = ~new_n50038_ & ~new_n50337_;
  assign new_n50804_ = ~new_n50336_ & new_n50803_;
  assign new_n50805_ = ~new_n50802_ & ~new_n50804_;
  assign new_n50806_ = ~\b[4]  & ~new_n50805_;
  assign new_n50807_ = ~new_n50057_ & new_n50061_;
  assign new_n50808_ = ~new_n50056_ & new_n50807_;
  assign new_n50809_ = ~new_n50058_ & ~new_n50061_;
  assign new_n50810_ = ~new_n50808_ & ~new_n50809_;
  assign new_n50811_ = ~new_n50338_ & ~new_n50810_;
  assign new_n50812_ = ~new_n50046_ & ~new_n50337_;
  assign new_n50813_ = ~new_n50336_ & new_n50812_;
  assign new_n50814_ = ~new_n50811_ & ~new_n50813_;
  assign new_n50815_ = ~\b[3]  & ~new_n50814_;
  assign new_n50816_ = new_n22029_ & ~new_n50054_;
  assign new_n50817_ = ~new_n50052_ & new_n50816_;
  assign new_n50818_ = ~new_n50056_ & ~new_n50817_;
  assign new_n50819_ = ~new_n50338_ & new_n50818_;
  assign new_n50820_ = ~new_n50051_ & ~new_n50337_;
  assign new_n50821_ = ~new_n50336_ & new_n50820_;
  assign new_n50822_ = ~new_n50819_ & ~new_n50821_;
  assign new_n50823_ = ~\b[2]  & ~new_n50822_;
  assign new_n50824_ = \b[0]  & ~new_n50338_;
  assign new_n50825_ = \a[8]  & ~new_n50824_;
  assign new_n50826_ = new_n22029_ & ~new_n50338_;
  assign new_n50827_ = ~new_n50825_ & ~new_n50826_;
  assign new_n50828_ = \b[1]  & ~new_n50827_;
  assign new_n50829_ = ~\b[1]  & ~new_n50826_;
  assign new_n50830_ = ~new_n50825_ & new_n50829_;
  assign new_n50831_ = ~new_n50828_ & ~new_n50830_;
  assign new_n50832_ = ~new_n22806_ & ~new_n50831_;
  assign new_n50833_ = ~\b[1]  & ~new_n50827_;
  assign new_n50834_ = ~new_n50832_ & ~new_n50833_;
  assign new_n50835_ = \b[2]  & ~new_n50821_;
  assign new_n50836_ = ~new_n50819_ & new_n50835_;
  assign new_n50837_ = ~new_n50823_ & ~new_n50836_;
  assign new_n50838_ = ~new_n50834_ & new_n50837_;
  assign new_n50839_ = ~new_n50823_ & ~new_n50838_;
  assign new_n50840_ = \b[3]  & ~new_n50813_;
  assign new_n50841_ = ~new_n50811_ & new_n50840_;
  assign new_n50842_ = ~new_n50815_ & ~new_n50841_;
  assign new_n50843_ = ~new_n50839_ & new_n50842_;
  assign new_n50844_ = ~new_n50815_ & ~new_n50843_;
  assign new_n50845_ = \b[4]  & ~new_n50804_;
  assign new_n50846_ = ~new_n50802_ & new_n50845_;
  assign new_n50847_ = ~new_n50806_ & ~new_n50846_;
  assign new_n50848_ = ~new_n50844_ & new_n50847_;
  assign new_n50849_ = ~new_n50806_ & ~new_n50848_;
  assign new_n50850_ = \b[5]  & ~new_n50795_;
  assign new_n50851_ = ~new_n50793_ & new_n50850_;
  assign new_n50852_ = ~new_n50797_ & ~new_n50851_;
  assign new_n50853_ = ~new_n50849_ & new_n50852_;
  assign new_n50854_ = ~new_n50797_ & ~new_n50853_;
  assign new_n50855_ = \b[6]  & ~new_n50786_;
  assign new_n50856_ = ~new_n50784_ & new_n50855_;
  assign new_n50857_ = ~new_n50788_ & ~new_n50856_;
  assign new_n50858_ = ~new_n50854_ & new_n50857_;
  assign new_n50859_ = ~new_n50788_ & ~new_n50858_;
  assign new_n50860_ = \b[7]  & ~new_n50777_;
  assign new_n50861_ = ~new_n50775_ & new_n50860_;
  assign new_n50862_ = ~new_n50779_ & ~new_n50861_;
  assign new_n50863_ = ~new_n50859_ & new_n50862_;
  assign new_n50864_ = ~new_n50779_ & ~new_n50863_;
  assign new_n50865_ = \b[8]  & ~new_n50768_;
  assign new_n50866_ = ~new_n50766_ & new_n50865_;
  assign new_n50867_ = ~new_n50770_ & ~new_n50866_;
  assign new_n50868_ = ~new_n50864_ & new_n50867_;
  assign new_n50869_ = ~new_n50770_ & ~new_n50868_;
  assign new_n50870_ = \b[9]  & ~new_n50759_;
  assign new_n50871_ = ~new_n50757_ & new_n50870_;
  assign new_n50872_ = ~new_n50761_ & ~new_n50871_;
  assign new_n50873_ = ~new_n50869_ & new_n50872_;
  assign new_n50874_ = ~new_n50761_ & ~new_n50873_;
  assign new_n50875_ = \b[10]  & ~new_n50750_;
  assign new_n50876_ = ~new_n50748_ & new_n50875_;
  assign new_n50877_ = ~new_n50752_ & ~new_n50876_;
  assign new_n50878_ = ~new_n50874_ & new_n50877_;
  assign new_n50879_ = ~new_n50752_ & ~new_n50878_;
  assign new_n50880_ = \b[11]  & ~new_n50741_;
  assign new_n50881_ = ~new_n50739_ & new_n50880_;
  assign new_n50882_ = ~new_n50743_ & ~new_n50881_;
  assign new_n50883_ = ~new_n50879_ & new_n50882_;
  assign new_n50884_ = ~new_n50743_ & ~new_n50883_;
  assign new_n50885_ = \b[12]  & ~new_n50732_;
  assign new_n50886_ = ~new_n50730_ & new_n50885_;
  assign new_n50887_ = ~new_n50734_ & ~new_n50886_;
  assign new_n50888_ = ~new_n50884_ & new_n50887_;
  assign new_n50889_ = ~new_n50734_ & ~new_n50888_;
  assign new_n50890_ = \b[13]  & ~new_n50723_;
  assign new_n50891_ = ~new_n50721_ & new_n50890_;
  assign new_n50892_ = ~new_n50725_ & ~new_n50891_;
  assign new_n50893_ = ~new_n50889_ & new_n50892_;
  assign new_n50894_ = ~new_n50725_ & ~new_n50893_;
  assign new_n50895_ = \b[14]  & ~new_n50714_;
  assign new_n50896_ = ~new_n50712_ & new_n50895_;
  assign new_n50897_ = ~new_n50716_ & ~new_n50896_;
  assign new_n50898_ = ~new_n50894_ & new_n50897_;
  assign new_n50899_ = ~new_n50716_ & ~new_n50898_;
  assign new_n50900_ = \b[15]  & ~new_n50705_;
  assign new_n50901_ = ~new_n50703_ & new_n50900_;
  assign new_n50902_ = ~new_n50707_ & ~new_n50901_;
  assign new_n50903_ = ~new_n50899_ & new_n50902_;
  assign new_n50904_ = ~new_n50707_ & ~new_n50903_;
  assign new_n50905_ = \b[16]  & ~new_n50696_;
  assign new_n50906_ = ~new_n50694_ & new_n50905_;
  assign new_n50907_ = ~new_n50698_ & ~new_n50906_;
  assign new_n50908_ = ~new_n50904_ & new_n50907_;
  assign new_n50909_ = ~new_n50698_ & ~new_n50908_;
  assign new_n50910_ = \b[17]  & ~new_n50687_;
  assign new_n50911_ = ~new_n50685_ & new_n50910_;
  assign new_n50912_ = ~new_n50689_ & ~new_n50911_;
  assign new_n50913_ = ~new_n50909_ & new_n50912_;
  assign new_n50914_ = ~new_n50689_ & ~new_n50913_;
  assign new_n50915_ = \b[18]  & ~new_n50678_;
  assign new_n50916_ = ~new_n50676_ & new_n50915_;
  assign new_n50917_ = ~new_n50680_ & ~new_n50916_;
  assign new_n50918_ = ~new_n50914_ & new_n50917_;
  assign new_n50919_ = ~new_n50680_ & ~new_n50918_;
  assign new_n50920_ = \b[19]  & ~new_n50669_;
  assign new_n50921_ = ~new_n50667_ & new_n50920_;
  assign new_n50922_ = ~new_n50671_ & ~new_n50921_;
  assign new_n50923_ = ~new_n50919_ & new_n50922_;
  assign new_n50924_ = ~new_n50671_ & ~new_n50923_;
  assign new_n50925_ = \b[20]  & ~new_n50660_;
  assign new_n50926_ = ~new_n50658_ & new_n50925_;
  assign new_n50927_ = ~new_n50662_ & ~new_n50926_;
  assign new_n50928_ = ~new_n50924_ & new_n50927_;
  assign new_n50929_ = ~new_n50662_ & ~new_n50928_;
  assign new_n50930_ = \b[21]  & ~new_n50651_;
  assign new_n50931_ = ~new_n50649_ & new_n50930_;
  assign new_n50932_ = ~new_n50653_ & ~new_n50931_;
  assign new_n50933_ = ~new_n50929_ & new_n50932_;
  assign new_n50934_ = ~new_n50653_ & ~new_n50933_;
  assign new_n50935_ = \b[22]  & ~new_n50642_;
  assign new_n50936_ = ~new_n50640_ & new_n50935_;
  assign new_n50937_ = ~new_n50644_ & ~new_n50936_;
  assign new_n50938_ = ~new_n50934_ & new_n50937_;
  assign new_n50939_ = ~new_n50644_ & ~new_n50938_;
  assign new_n50940_ = \b[23]  & ~new_n50633_;
  assign new_n50941_ = ~new_n50631_ & new_n50940_;
  assign new_n50942_ = ~new_n50635_ & ~new_n50941_;
  assign new_n50943_ = ~new_n50939_ & new_n50942_;
  assign new_n50944_ = ~new_n50635_ & ~new_n50943_;
  assign new_n50945_ = \b[24]  & ~new_n50624_;
  assign new_n50946_ = ~new_n50622_ & new_n50945_;
  assign new_n50947_ = ~new_n50626_ & ~new_n50946_;
  assign new_n50948_ = ~new_n50944_ & new_n50947_;
  assign new_n50949_ = ~new_n50626_ & ~new_n50948_;
  assign new_n50950_ = \b[25]  & ~new_n50615_;
  assign new_n50951_ = ~new_n50613_ & new_n50950_;
  assign new_n50952_ = ~new_n50617_ & ~new_n50951_;
  assign new_n50953_ = ~new_n50949_ & new_n50952_;
  assign new_n50954_ = ~new_n50617_ & ~new_n50953_;
  assign new_n50955_ = \b[26]  & ~new_n50606_;
  assign new_n50956_ = ~new_n50604_ & new_n50955_;
  assign new_n50957_ = ~new_n50608_ & ~new_n50956_;
  assign new_n50958_ = ~new_n50954_ & new_n50957_;
  assign new_n50959_ = ~new_n50608_ & ~new_n50958_;
  assign new_n50960_ = \b[27]  & ~new_n50597_;
  assign new_n50961_ = ~new_n50595_ & new_n50960_;
  assign new_n50962_ = ~new_n50599_ & ~new_n50961_;
  assign new_n50963_ = ~new_n50959_ & new_n50962_;
  assign new_n50964_ = ~new_n50599_ & ~new_n50963_;
  assign new_n50965_ = \b[28]  & ~new_n50588_;
  assign new_n50966_ = ~new_n50586_ & new_n50965_;
  assign new_n50967_ = ~new_n50590_ & ~new_n50966_;
  assign new_n50968_ = ~new_n50964_ & new_n50967_;
  assign new_n50969_ = ~new_n50590_ & ~new_n50968_;
  assign new_n50970_ = \b[29]  & ~new_n50579_;
  assign new_n50971_ = ~new_n50577_ & new_n50970_;
  assign new_n50972_ = ~new_n50581_ & ~new_n50971_;
  assign new_n50973_ = ~new_n50969_ & new_n50972_;
  assign new_n50974_ = ~new_n50581_ & ~new_n50973_;
  assign new_n50975_ = \b[30]  & ~new_n50570_;
  assign new_n50976_ = ~new_n50568_ & new_n50975_;
  assign new_n50977_ = ~new_n50572_ & ~new_n50976_;
  assign new_n50978_ = ~new_n50974_ & new_n50977_;
  assign new_n50979_ = ~new_n50572_ & ~new_n50978_;
  assign new_n50980_ = \b[31]  & ~new_n50561_;
  assign new_n50981_ = ~new_n50559_ & new_n50980_;
  assign new_n50982_ = ~new_n50563_ & ~new_n50981_;
  assign new_n50983_ = ~new_n50979_ & new_n50982_;
  assign new_n50984_ = ~new_n50563_ & ~new_n50983_;
  assign new_n50985_ = \b[32]  & ~new_n50552_;
  assign new_n50986_ = ~new_n50550_ & new_n50985_;
  assign new_n50987_ = ~new_n50554_ & ~new_n50986_;
  assign new_n50988_ = ~new_n50984_ & new_n50987_;
  assign new_n50989_ = ~new_n50554_ & ~new_n50988_;
  assign new_n50990_ = \b[33]  & ~new_n50543_;
  assign new_n50991_ = ~new_n50541_ & new_n50990_;
  assign new_n50992_ = ~new_n50545_ & ~new_n50991_;
  assign new_n50993_ = ~new_n50989_ & new_n50992_;
  assign new_n50994_ = ~new_n50545_ & ~new_n50993_;
  assign new_n50995_ = \b[34]  & ~new_n50534_;
  assign new_n50996_ = ~new_n50532_ & new_n50995_;
  assign new_n50997_ = ~new_n50536_ & ~new_n50996_;
  assign new_n50998_ = ~new_n50994_ & new_n50997_;
  assign new_n50999_ = ~new_n50536_ & ~new_n50998_;
  assign new_n51000_ = \b[35]  & ~new_n50525_;
  assign new_n51001_ = ~new_n50523_ & new_n51000_;
  assign new_n51002_ = ~new_n50527_ & ~new_n51001_;
  assign new_n51003_ = ~new_n50999_ & new_n51002_;
  assign new_n51004_ = ~new_n50527_ & ~new_n51003_;
  assign new_n51005_ = \b[36]  & ~new_n50516_;
  assign new_n51006_ = ~new_n50514_ & new_n51005_;
  assign new_n51007_ = ~new_n50518_ & ~new_n51006_;
  assign new_n51008_ = ~new_n51004_ & new_n51007_;
  assign new_n51009_ = ~new_n50518_ & ~new_n51008_;
  assign new_n51010_ = \b[37]  & ~new_n50507_;
  assign new_n51011_ = ~new_n50505_ & new_n51010_;
  assign new_n51012_ = ~new_n50509_ & ~new_n51011_;
  assign new_n51013_ = ~new_n51009_ & new_n51012_;
  assign new_n51014_ = ~new_n50509_ & ~new_n51013_;
  assign new_n51015_ = \b[38]  & ~new_n50498_;
  assign new_n51016_ = ~new_n50496_ & new_n51015_;
  assign new_n51017_ = ~new_n50500_ & ~new_n51016_;
  assign new_n51018_ = ~new_n51014_ & new_n51017_;
  assign new_n51019_ = ~new_n50500_ & ~new_n51018_;
  assign new_n51020_ = \b[39]  & ~new_n50489_;
  assign new_n51021_ = ~new_n50487_ & new_n51020_;
  assign new_n51022_ = ~new_n50491_ & ~new_n51021_;
  assign new_n51023_ = ~new_n51019_ & new_n51022_;
  assign new_n51024_ = ~new_n50491_ & ~new_n51023_;
  assign new_n51025_ = \b[40]  & ~new_n50480_;
  assign new_n51026_ = ~new_n50478_ & new_n51025_;
  assign new_n51027_ = ~new_n50482_ & ~new_n51026_;
  assign new_n51028_ = ~new_n51024_ & new_n51027_;
  assign new_n51029_ = ~new_n50482_ & ~new_n51028_;
  assign new_n51030_ = \b[41]  & ~new_n50471_;
  assign new_n51031_ = ~new_n50469_ & new_n51030_;
  assign new_n51032_ = ~new_n50473_ & ~new_n51031_;
  assign new_n51033_ = ~new_n51029_ & new_n51032_;
  assign new_n51034_ = ~new_n50473_ & ~new_n51033_;
  assign new_n51035_ = \b[42]  & ~new_n50462_;
  assign new_n51036_ = ~new_n50460_ & new_n51035_;
  assign new_n51037_ = ~new_n50464_ & ~new_n51036_;
  assign new_n51038_ = ~new_n51034_ & new_n51037_;
  assign new_n51039_ = ~new_n50464_ & ~new_n51038_;
  assign new_n51040_ = \b[43]  & ~new_n50453_;
  assign new_n51041_ = ~new_n50451_ & new_n51040_;
  assign new_n51042_ = ~new_n50455_ & ~new_n51041_;
  assign new_n51043_ = ~new_n51039_ & new_n51042_;
  assign new_n51044_ = ~new_n50455_ & ~new_n51043_;
  assign new_n51045_ = \b[44]  & ~new_n50444_;
  assign new_n51046_ = ~new_n50442_ & new_n51045_;
  assign new_n51047_ = ~new_n50446_ & ~new_n51046_;
  assign new_n51048_ = ~new_n51044_ & new_n51047_;
  assign new_n51049_ = ~new_n50446_ & ~new_n51048_;
  assign new_n51050_ = \b[45]  & ~new_n50435_;
  assign new_n51051_ = ~new_n50433_ & new_n51050_;
  assign new_n51052_ = ~new_n50437_ & ~new_n51051_;
  assign new_n51053_ = ~new_n51049_ & new_n51052_;
  assign new_n51054_ = ~new_n50437_ & ~new_n51053_;
  assign new_n51055_ = \b[46]  & ~new_n50426_;
  assign new_n51056_ = ~new_n50424_ & new_n51055_;
  assign new_n51057_ = ~new_n50428_ & ~new_n51056_;
  assign new_n51058_ = ~new_n51054_ & new_n51057_;
  assign new_n51059_ = ~new_n50428_ & ~new_n51058_;
  assign new_n51060_ = \b[47]  & ~new_n50417_;
  assign new_n51061_ = ~new_n50415_ & new_n51060_;
  assign new_n51062_ = ~new_n50419_ & ~new_n51061_;
  assign new_n51063_ = ~new_n51059_ & new_n51062_;
  assign new_n51064_ = ~new_n50419_ & ~new_n51063_;
  assign new_n51065_ = \b[48]  & ~new_n50408_;
  assign new_n51066_ = ~new_n50406_ & new_n51065_;
  assign new_n51067_ = ~new_n50410_ & ~new_n51066_;
  assign new_n51068_ = ~new_n51064_ & new_n51067_;
  assign new_n51069_ = ~new_n50410_ & ~new_n51068_;
  assign new_n51070_ = \b[49]  & ~new_n50399_;
  assign new_n51071_ = ~new_n50397_ & new_n51070_;
  assign new_n51072_ = ~new_n50401_ & ~new_n51071_;
  assign new_n51073_ = ~new_n51069_ & new_n51072_;
  assign new_n51074_ = ~new_n50401_ & ~new_n51073_;
  assign new_n51075_ = \b[50]  & ~new_n50390_;
  assign new_n51076_ = ~new_n50388_ & new_n51075_;
  assign new_n51077_ = ~new_n50392_ & ~new_n51076_;
  assign new_n51078_ = ~new_n51074_ & new_n51077_;
  assign new_n51079_ = ~new_n50392_ & ~new_n51078_;
  assign new_n51080_ = \b[51]  & ~new_n50381_;
  assign new_n51081_ = ~new_n50379_ & new_n51080_;
  assign new_n51082_ = ~new_n50383_ & ~new_n51081_;
  assign new_n51083_ = ~new_n51079_ & new_n51082_;
  assign new_n51084_ = ~new_n50383_ & ~new_n51083_;
  assign new_n51085_ = \b[52]  & ~new_n50372_;
  assign new_n51086_ = ~new_n50370_ & new_n51085_;
  assign new_n51087_ = ~new_n50374_ & ~new_n51086_;
  assign new_n51088_ = ~new_n51084_ & new_n51087_;
  assign new_n51089_ = ~new_n50374_ & ~new_n51088_;
  assign new_n51090_ = \b[53]  & ~new_n50363_;
  assign new_n51091_ = ~new_n50361_ & new_n51090_;
  assign new_n51092_ = ~new_n50365_ & ~new_n51091_;
  assign new_n51093_ = ~new_n51089_ & new_n51092_;
  assign new_n51094_ = ~new_n50365_ & ~new_n51093_;
  assign new_n51095_ = \b[54]  & ~new_n50354_;
  assign new_n51096_ = ~new_n50352_ & new_n51095_;
  assign new_n51097_ = ~new_n50356_ & ~new_n51096_;
  assign new_n51098_ = ~new_n51094_ & new_n51097_;
  assign new_n51099_ = ~new_n50356_ & ~new_n51098_;
  assign new_n51100_ = \b[55]  & ~new_n50345_;
  assign new_n51101_ = ~new_n50343_ & new_n51100_;
  assign new_n51102_ = ~new_n50347_ & ~new_n51101_;
  assign new_n51103_ = ~new_n51099_ & new_n51102_;
  assign new_n51104_ = ~new_n50347_ & ~new_n51103_;
  assign new_n51105_ = ~new_n49580_ & ~new_n50333_;
  assign new_n51106_ = ~new_n50331_ & new_n51105_;
  assign new_n51107_ = ~new_n50322_ & new_n51106_;
  assign new_n51108_ = ~new_n50331_ & ~new_n50333_;
  assign new_n51109_ = ~new_n50323_ & ~new_n51108_;
  assign new_n51110_ = ~new_n51107_ & ~new_n51109_;
  assign new_n51111_ = ~new_n50338_ & ~new_n51110_;
  assign new_n51112_ = ~new_n50330_ & ~new_n50337_;
  assign new_n51113_ = ~new_n50336_ & new_n51112_;
  assign new_n51114_ = ~new_n51111_ & ~new_n51113_;
  assign new_n51115_ = ~\b[56]  & ~new_n51114_;
  assign new_n51116_ = \b[56]  & ~new_n51113_;
  assign new_n51117_ = ~new_n51111_ & new_n51116_;
  assign new_n51118_ = new_n407_ & ~new_n51117_;
  assign new_n51119_ = ~new_n51115_ & new_n51118_;
  assign new_n51120_ = ~new_n51104_ & new_n51119_;
  assign new_n51121_ = new_n337_ & ~new_n51114_;
  assign new_n51122_ = ~new_n51120_ & ~new_n51121_;
  assign new_n51123_ = ~new_n50356_ & new_n51102_;
  assign new_n51124_ = ~new_n51098_ & new_n51123_;
  assign new_n51125_ = ~new_n51099_ & ~new_n51102_;
  assign new_n51126_ = ~new_n51124_ & ~new_n51125_;
  assign new_n51127_ = ~new_n51122_ & ~new_n51126_;
  assign new_n51128_ = ~new_n50346_ & ~new_n51121_;
  assign new_n51129_ = ~new_n51120_ & new_n51128_;
  assign new_n51130_ = ~new_n51127_ & ~new_n51129_;
  assign new_n51131_ = ~new_n50347_ & ~new_n51117_;
  assign new_n51132_ = ~new_n51115_ & new_n51131_;
  assign new_n51133_ = ~new_n51103_ & new_n51132_;
  assign new_n51134_ = ~new_n51115_ & ~new_n51117_;
  assign new_n51135_ = ~new_n51104_ & ~new_n51134_;
  assign new_n51136_ = ~new_n51133_ & ~new_n51135_;
  assign new_n51137_ = ~new_n51122_ & ~new_n51136_;
  assign new_n51138_ = ~new_n51114_ & ~new_n51121_;
  assign new_n51139_ = ~new_n51120_ & new_n51138_;
  assign new_n51140_ = ~new_n51137_ & ~new_n51139_;
  assign new_n51141_ = ~\b[57]  & ~new_n51140_;
  assign new_n51142_ = ~\b[56]  & ~new_n51130_;
  assign new_n51143_ = ~new_n50365_ & new_n51097_;
  assign new_n51144_ = ~new_n51093_ & new_n51143_;
  assign new_n51145_ = ~new_n51094_ & ~new_n51097_;
  assign new_n51146_ = ~new_n51144_ & ~new_n51145_;
  assign new_n51147_ = ~new_n51122_ & ~new_n51146_;
  assign new_n51148_ = ~new_n50355_ & ~new_n51121_;
  assign new_n51149_ = ~new_n51120_ & new_n51148_;
  assign new_n51150_ = ~new_n51147_ & ~new_n51149_;
  assign new_n51151_ = ~\b[55]  & ~new_n51150_;
  assign new_n51152_ = ~new_n50374_ & new_n51092_;
  assign new_n51153_ = ~new_n51088_ & new_n51152_;
  assign new_n51154_ = ~new_n51089_ & ~new_n51092_;
  assign new_n51155_ = ~new_n51153_ & ~new_n51154_;
  assign new_n51156_ = ~new_n51122_ & ~new_n51155_;
  assign new_n51157_ = ~new_n50364_ & ~new_n51121_;
  assign new_n51158_ = ~new_n51120_ & new_n51157_;
  assign new_n51159_ = ~new_n51156_ & ~new_n51158_;
  assign new_n51160_ = ~\b[54]  & ~new_n51159_;
  assign new_n51161_ = ~new_n50383_ & new_n51087_;
  assign new_n51162_ = ~new_n51083_ & new_n51161_;
  assign new_n51163_ = ~new_n51084_ & ~new_n51087_;
  assign new_n51164_ = ~new_n51162_ & ~new_n51163_;
  assign new_n51165_ = ~new_n51122_ & ~new_n51164_;
  assign new_n51166_ = ~new_n50373_ & ~new_n51121_;
  assign new_n51167_ = ~new_n51120_ & new_n51166_;
  assign new_n51168_ = ~new_n51165_ & ~new_n51167_;
  assign new_n51169_ = ~\b[53]  & ~new_n51168_;
  assign new_n51170_ = ~new_n50392_ & new_n51082_;
  assign new_n51171_ = ~new_n51078_ & new_n51170_;
  assign new_n51172_ = ~new_n51079_ & ~new_n51082_;
  assign new_n51173_ = ~new_n51171_ & ~new_n51172_;
  assign new_n51174_ = ~new_n51122_ & ~new_n51173_;
  assign new_n51175_ = ~new_n50382_ & ~new_n51121_;
  assign new_n51176_ = ~new_n51120_ & new_n51175_;
  assign new_n51177_ = ~new_n51174_ & ~new_n51176_;
  assign new_n51178_ = ~\b[52]  & ~new_n51177_;
  assign new_n51179_ = ~new_n50401_ & new_n51077_;
  assign new_n51180_ = ~new_n51073_ & new_n51179_;
  assign new_n51181_ = ~new_n51074_ & ~new_n51077_;
  assign new_n51182_ = ~new_n51180_ & ~new_n51181_;
  assign new_n51183_ = ~new_n51122_ & ~new_n51182_;
  assign new_n51184_ = ~new_n50391_ & ~new_n51121_;
  assign new_n51185_ = ~new_n51120_ & new_n51184_;
  assign new_n51186_ = ~new_n51183_ & ~new_n51185_;
  assign new_n51187_ = ~\b[51]  & ~new_n51186_;
  assign new_n51188_ = ~new_n50410_ & new_n51072_;
  assign new_n51189_ = ~new_n51068_ & new_n51188_;
  assign new_n51190_ = ~new_n51069_ & ~new_n51072_;
  assign new_n51191_ = ~new_n51189_ & ~new_n51190_;
  assign new_n51192_ = ~new_n51122_ & ~new_n51191_;
  assign new_n51193_ = ~new_n50400_ & ~new_n51121_;
  assign new_n51194_ = ~new_n51120_ & new_n51193_;
  assign new_n51195_ = ~new_n51192_ & ~new_n51194_;
  assign new_n51196_ = ~\b[50]  & ~new_n51195_;
  assign new_n51197_ = ~new_n50419_ & new_n51067_;
  assign new_n51198_ = ~new_n51063_ & new_n51197_;
  assign new_n51199_ = ~new_n51064_ & ~new_n51067_;
  assign new_n51200_ = ~new_n51198_ & ~new_n51199_;
  assign new_n51201_ = ~new_n51122_ & ~new_n51200_;
  assign new_n51202_ = ~new_n50409_ & ~new_n51121_;
  assign new_n51203_ = ~new_n51120_ & new_n51202_;
  assign new_n51204_ = ~new_n51201_ & ~new_n51203_;
  assign new_n51205_ = ~\b[49]  & ~new_n51204_;
  assign new_n51206_ = ~new_n50428_ & new_n51062_;
  assign new_n51207_ = ~new_n51058_ & new_n51206_;
  assign new_n51208_ = ~new_n51059_ & ~new_n51062_;
  assign new_n51209_ = ~new_n51207_ & ~new_n51208_;
  assign new_n51210_ = ~new_n51122_ & ~new_n51209_;
  assign new_n51211_ = ~new_n50418_ & ~new_n51121_;
  assign new_n51212_ = ~new_n51120_ & new_n51211_;
  assign new_n51213_ = ~new_n51210_ & ~new_n51212_;
  assign new_n51214_ = ~\b[48]  & ~new_n51213_;
  assign new_n51215_ = ~new_n50437_ & new_n51057_;
  assign new_n51216_ = ~new_n51053_ & new_n51215_;
  assign new_n51217_ = ~new_n51054_ & ~new_n51057_;
  assign new_n51218_ = ~new_n51216_ & ~new_n51217_;
  assign new_n51219_ = ~new_n51122_ & ~new_n51218_;
  assign new_n51220_ = ~new_n50427_ & ~new_n51121_;
  assign new_n51221_ = ~new_n51120_ & new_n51220_;
  assign new_n51222_ = ~new_n51219_ & ~new_n51221_;
  assign new_n51223_ = ~\b[47]  & ~new_n51222_;
  assign new_n51224_ = ~new_n50446_ & new_n51052_;
  assign new_n51225_ = ~new_n51048_ & new_n51224_;
  assign new_n51226_ = ~new_n51049_ & ~new_n51052_;
  assign new_n51227_ = ~new_n51225_ & ~new_n51226_;
  assign new_n51228_ = ~new_n51122_ & ~new_n51227_;
  assign new_n51229_ = ~new_n50436_ & ~new_n51121_;
  assign new_n51230_ = ~new_n51120_ & new_n51229_;
  assign new_n51231_ = ~new_n51228_ & ~new_n51230_;
  assign new_n51232_ = ~\b[46]  & ~new_n51231_;
  assign new_n51233_ = ~new_n50455_ & new_n51047_;
  assign new_n51234_ = ~new_n51043_ & new_n51233_;
  assign new_n51235_ = ~new_n51044_ & ~new_n51047_;
  assign new_n51236_ = ~new_n51234_ & ~new_n51235_;
  assign new_n51237_ = ~new_n51122_ & ~new_n51236_;
  assign new_n51238_ = ~new_n50445_ & ~new_n51121_;
  assign new_n51239_ = ~new_n51120_ & new_n51238_;
  assign new_n51240_ = ~new_n51237_ & ~new_n51239_;
  assign new_n51241_ = ~\b[45]  & ~new_n51240_;
  assign new_n51242_ = ~new_n50464_ & new_n51042_;
  assign new_n51243_ = ~new_n51038_ & new_n51242_;
  assign new_n51244_ = ~new_n51039_ & ~new_n51042_;
  assign new_n51245_ = ~new_n51243_ & ~new_n51244_;
  assign new_n51246_ = ~new_n51122_ & ~new_n51245_;
  assign new_n51247_ = ~new_n50454_ & ~new_n51121_;
  assign new_n51248_ = ~new_n51120_ & new_n51247_;
  assign new_n51249_ = ~new_n51246_ & ~new_n51248_;
  assign new_n51250_ = ~\b[44]  & ~new_n51249_;
  assign new_n51251_ = ~new_n50473_ & new_n51037_;
  assign new_n51252_ = ~new_n51033_ & new_n51251_;
  assign new_n51253_ = ~new_n51034_ & ~new_n51037_;
  assign new_n51254_ = ~new_n51252_ & ~new_n51253_;
  assign new_n51255_ = ~new_n51122_ & ~new_n51254_;
  assign new_n51256_ = ~new_n50463_ & ~new_n51121_;
  assign new_n51257_ = ~new_n51120_ & new_n51256_;
  assign new_n51258_ = ~new_n51255_ & ~new_n51257_;
  assign new_n51259_ = ~\b[43]  & ~new_n51258_;
  assign new_n51260_ = ~new_n50482_ & new_n51032_;
  assign new_n51261_ = ~new_n51028_ & new_n51260_;
  assign new_n51262_ = ~new_n51029_ & ~new_n51032_;
  assign new_n51263_ = ~new_n51261_ & ~new_n51262_;
  assign new_n51264_ = ~new_n51122_ & ~new_n51263_;
  assign new_n51265_ = ~new_n50472_ & ~new_n51121_;
  assign new_n51266_ = ~new_n51120_ & new_n51265_;
  assign new_n51267_ = ~new_n51264_ & ~new_n51266_;
  assign new_n51268_ = ~\b[42]  & ~new_n51267_;
  assign new_n51269_ = ~new_n50491_ & new_n51027_;
  assign new_n51270_ = ~new_n51023_ & new_n51269_;
  assign new_n51271_ = ~new_n51024_ & ~new_n51027_;
  assign new_n51272_ = ~new_n51270_ & ~new_n51271_;
  assign new_n51273_ = ~new_n51122_ & ~new_n51272_;
  assign new_n51274_ = ~new_n50481_ & ~new_n51121_;
  assign new_n51275_ = ~new_n51120_ & new_n51274_;
  assign new_n51276_ = ~new_n51273_ & ~new_n51275_;
  assign new_n51277_ = ~\b[41]  & ~new_n51276_;
  assign new_n51278_ = ~new_n50500_ & new_n51022_;
  assign new_n51279_ = ~new_n51018_ & new_n51278_;
  assign new_n51280_ = ~new_n51019_ & ~new_n51022_;
  assign new_n51281_ = ~new_n51279_ & ~new_n51280_;
  assign new_n51282_ = ~new_n51122_ & ~new_n51281_;
  assign new_n51283_ = ~new_n50490_ & ~new_n51121_;
  assign new_n51284_ = ~new_n51120_ & new_n51283_;
  assign new_n51285_ = ~new_n51282_ & ~new_n51284_;
  assign new_n51286_ = ~\b[40]  & ~new_n51285_;
  assign new_n51287_ = ~new_n50509_ & new_n51017_;
  assign new_n51288_ = ~new_n51013_ & new_n51287_;
  assign new_n51289_ = ~new_n51014_ & ~new_n51017_;
  assign new_n51290_ = ~new_n51288_ & ~new_n51289_;
  assign new_n51291_ = ~new_n51122_ & ~new_n51290_;
  assign new_n51292_ = ~new_n50499_ & ~new_n51121_;
  assign new_n51293_ = ~new_n51120_ & new_n51292_;
  assign new_n51294_ = ~new_n51291_ & ~new_n51293_;
  assign new_n51295_ = ~\b[39]  & ~new_n51294_;
  assign new_n51296_ = ~new_n50518_ & new_n51012_;
  assign new_n51297_ = ~new_n51008_ & new_n51296_;
  assign new_n51298_ = ~new_n51009_ & ~new_n51012_;
  assign new_n51299_ = ~new_n51297_ & ~new_n51298_;
  assign new_n51300_ = ~new_n51122_ & ~new_n51299_;
  assign new_n51301_ = ~new_n50508_ & ~new_n51121_;
  assign new_n51302_ = ~new_n51120_ & new_n51301_;
  assign new_n51303_ = ~new_n51300_ & ~new_n51302_;
  assign new_n51304_ = ~\b[38]  & ~new_n51303_;
  assign new_n51305_ = ~new_n50527_ & new_n51007_;
  assign new_n51306_ = ~new_n51003_ & new_n51305_;
  assign new_n51307_ = ~new_n51004_ & ~new_n51007_;
  assign new_n51308_ = ~new_n51306_ & ~new_n51307_;
  assign new_n51309_ = ~new_n51122_ & ~new_n51308_;
  assign new_n51310_ = ~new_n50517_ & ~new_n51121_;
  assign new_n51311_ = ~new_n51120_ & new_n51310_;
  assign new_n51312_ = ~new_n51309_ & ~new_n51311_;
  assign new_n51313_ = ~\b[37]  & ~new_n51312_;
  assign new_n51314_ = ~new_n50536_ & new_n51002_;
  assign new_n51315_ = ~new_n50998_ & new_n51314_;
  assign new_n51316_ = ~new_n50999_ & ~new_n51002_;
  assign new_n51317_ = ~new_n51315_ & ~new_n51316_;
  assign new_n51318_ = ~new_n51122_ & ~new_n51317_;
  assign new_n51319_ = ~new_n50526_ & ~new_n51121_;
  assign new_n51320_ = ~new_n51120_ & new_n51319_;
  assign new_n51321_ = ~new_n51318_ & ~new_n51320_;
  assign new_n51322_ = ~\b[36]  & ~new_n51321_;
  assign new_n51323_ = ~new_n50545_ & new_n50997_;
  assign new_n51324_ = ~new_n50993_ & new_n51323_;
  assign new_n51325_ = ~new_n50994_ & ~new_n50997_;
  assign new_n51326_ = ~new_n51324_ & ~new_n51325_;
  assign new_n51327_ = ~new_n51122_ & ~new_n51326_;
  assign new_n51328_ = ~new_n50535_ & ~new_n51121_;
  assign new_n51329_ = ~new_n51120_ & new_n51328_;
  assign new_n51330_ = ~new_n51327_ & ~new_n51329_;
  assign new_n51331_ = ~\b[35]  & ~new_n51330_;
  assign new_n51332_ = ~new_n50554_ & new_n50992_;
  assign new_n51333_ = ~new_n50988_ & new_n51332_;
  assign new_n51334_ = ~new_n50989_ & ~new_n50992_;
  assign new_n51335_ = ~new_n51333_ & ~new_n51334_;
  assign new_n51336_ = ~new_n51122_ & ~new_n51335_;
  assign new_n51337_ = ~new_n50544_ & ~new_n51121_;
  assign new_n51338_ = ~new_n51120_ & new_n51337_;
  assign new_n51339_ = ~new_n51336_ & ~new_n51338_;
  assign new_n51340_ = ~\b[34]  & ~new_n51339_;
  assign new_n51341_ = ~new_n50563_ & new_n50987_;
  assign new_n51342_ = ~new_n50983_ & new_n51341_;
  assign new_n51343_ = ~new_n50984_ & ~new_n50987_;
  assign new_n51344_ = ~new_n51342_ & ~new_n51343_;
  assign new_n51345_ = ~new_n51122_ & ~new_n51344_;
  assign new_n51346_ = ~new_n50553_ & ~new_n51121_;
  assign new_n51347_ = ~new_n51120_ & new_n51346_;
  assign new_n51348_ = ~new_n51345_ & ~new_n51347_;
  assign new_n51349_ = ~\b[33]  & ~new_n51348_;
  assign new_n51350_ = ~new_n50572_ & new_n50982_;
  assign new_n51351_ = ~new_n50978_ & new_n51350_;
  assign new_n51352_ = ~new_n50979_ & ~new_n50982_;
  assign new_n51353_ = ~new_n51351_ & ~new_n51352_;
  assign new_n51354_ = ~new_n51122_ & ~new_n51353_;
  assign new_n51355_ = ~new_n50562_ & ~new_n51121_;
  assign new_n51356_ = ~new_n51120_ & new_n51355_;
  assign new_n51357_ = ~new_n51354_ & ~new_n51356_;
  assign new_n51358_ = ~\b[32]  & ~new_n51357_;
  assign new_n51359_ = ~new_n50581_ & new_n50977_;
  assign new_n51360_ = ~new_n50973_ & new_n51359_;
  assign new_n51361_ = ~new_n50974_ & ~new_n50977_;
  assign new_n51362_ = ~new_n51360_ & ~new_n51361_;
  assign new_n51363_ = ~new_n51122_ & ~new_n51362_;
  assign new_n51364_ = ~new_n50571_ & ~new_n51121_;
  assign new_n51365_ = ~new_n51120_ & new_n51364_;
  assign new_n51366_ = ~new_n51363_ & ~new_n51365_;
  assign new_n51367_ = ~\b[31]  & ~new_n51366_;
  assign new_n51368_ = ~new_n50590_ & new_n50972_;
  assign new_n51369_ = ~new_n50968_ & new_n51368_;
  assign new_n51370_ = ~new_n50969_ & ~new_n50972_;
  assign new_n51371_ = ~new_n51369_ & ~new_n51370_;
  assign new_n51372_ = ~new_n51122_ & ~new_n51371_;
  assign new_n51373_ = ~new_n50580_ & ~new_n51121_;
  assign new_n51374_ = ~new_n51120_ & new_n51373_;
  assign new_n51375_ = ~new_n51372_ & ~new_n51374_;
  assign new_n51376_ = ~\b[30]  & ~new_n51375_;
  assign new_n51377_ = ~new_n50599_ & new_n50967_;
  assign new_n51378_ = ~new_n50963_ & new_n51377_;
  assign new_n51379_ = ~new_n50964_ & ~new_n50967_;
  assign new_n51380_ = ~new_n51378_ & ~new_n51379_;
  assign new_n51381_ = ~new_n51122_ & ~new_n51380_;
  assign new_n51382_ = ~new_n50589_ & ~new_n51121_;
  assign new_n51383_ = ~new_n51120_ & new_n51382_;
  assign new_n51384_ = ~new_n51381_ & ~new_n51383_;
  assign new_n51385_ = ~\b[29]  & ~new_n51384_;
  assign new_n51386_ = ~new_n50608_ & new_n50962_;
  assign new_n51387_ = ~new_n50958_ & new_n51386_;
  assign new_n51388_ = ~new_n50959_ & ~new_n50962_;
  assign new_n51389_ = ~new_n51387_ & ~new_n51388_;
  assign new_n51390_ = ~new_n51122_ & ~new_n51389_;
  assign new_n51391_ = ~new_n50598_ & ~new_n51121_;
  assign new_n51392_ = ~new_n51120_ & new_n51391_;
  assign new_n51393_ = ~new_n51390_ & ~new_n51392_;
  assign new_n51394_ = ~\b[28]  & ~new_n51393_;
  assign new_n51395_ = ~new_n50617_ & new_n50957_;
  assign new_n51396_ = ~new_n50953_ & new_n51395_;
  assign new_n51397_ = ~new_n50954_ & ~new_n50957_;
  assign new_n51398_ = ~new_n51396_ & ~new_n51397_;
  assign new_n51399_ = ~new_n51122_ & ~new_n51398_;
  assign new_n51400_ = ~new_n50607_ & ~new_n51121_;
  assign new_n51401_ = ~new_n51120_ & new_n51400_;
  assign new_n51402_ = ~new_n51399_ & ~new_n51401_;
  assign new_n51403_ = ~\b[27]  & ~new_n51402_;
  assign new_n51404_ = ~new_n50626_ & new_n50952_;
  assign new_n51405_ = ~new_n50948_ & new_n51404_;
  assign new_n51406_ = ~new_n50949_ & ~new_n50952_;
  assign new_n51407_ = ~new_n51405_ & ~new_n51406_;
  assign new_n51408_ = ~new_n51122_ & ~new_n51407_;
  assign new_n51409_ = ~new_n50616_ & ~new_n51121_;
  assign new_n51410_ = ~new_n51120_ & new_n51409_;
  assign new_n51411_ = ~new_n51408_ & ~new_n51410_;
  assign new_n51412_ = ~\b[26]  & ~new_n51411_;
  assign new_n51413_ = ~new_n50635_ & new_n50947_;
  assign new_n51414_ = ~new_n50943_ & new_n51413_;
  assign new_n51415_ = ~new_n50944_ & ~new_n50947_;
  assign new_n51416_ = ~new_n51414_ & ~new_n51415_;
  assign new_n51417_ = ~new_n51122_ & ~new_n51416_;
  assign new_n51418_ = ~new_n50625_ & ~new_n51121_;
  assign new_n51419_ = ~new_n51120_ & new_n51418_;
  assign new_n51420_ = ~new_n51417_ & ~new_n51419_;
  assign new_n51421_ = ~\b[25]  & ~new_n51420_;
  assign new_n51422_ = ~new_n50644_ & new_n50942_;
  assign new_n51423_ = ~new_n50938_ & new_n51422_;
  assign new_n51424_ = ~new_n50939_ & ~new_n50942_;
  assign new_n51425_ = ~new_n51423_ & ~new_n51424_;
  assign new_n51426_ = ~new_n51122_ & ~new_n51425_;
  assign new_n51427_ = ~new_n50634_ & ~new_n51121_;
  assign new_n51428_ = ~new_n51120_ & new_n51427_;
  assign new_n51429_ = ~new_n51426_ & ~new_n51428_;
  assign new_n51430_ = ~\b[24]  & ~new_n51429_;
  assign new_n51431_ = ~new_n50653_ & new_n50937_;
  assign new_n51432_ = ~new_n50933_ & new_n51431_;
  assign new_n51433_ = ~new_n50934_ & ~new_n50937_;
  assign new_n51434_ = ~new_n51432_ & ~new_n51433_;
  assign new_n51435_ = ~new_n51122_ & ~new_n51434_;
  assign new_n51436_ = ~new_n50643_ & ~new_n51121_;
  assign new_n51437_ = ~new_n51120_ & new_n51436_;
  assign new_n51438_ = ~new_n51435_ & ~new_n51437_;
  assign new_n51439_ = ~\b[23]  & ~new_n51438_;
  assign new_n51440_ = ~new_n50662_ & new_n50932_;
  assign new_n51441_ = ~new_n50928_ & new_n51440_;
  assign new_n51442_ = ~new_n50929_ & ~new_n50932_;
  assign new_n51443_ = ~new_n51441_ & ~new_n51442_;
  assign new_n51444_ = ~new_n51122_ & ~new_n51443_;
  assign new_n51445_ = ~new_n50652_ & ~new_n51121_;
  assign new_n51446_ = ~new_n51120_ & new_n51445_;
  assign new_n51447_ = ~new_n51444_ & ~new_n51446_;
  assign new_n51448_ = ~\b[22]  & ~new_n51447_;
  assign new_n51449_ = ~new_n50671_ & new_n50927_;
  assign new_n51450_ = ~new_n50923_ & new_n51449_;
  assign new_n51451_ = ~new_n50924_ & ~new_n50927_;
  assign new_n51452_ = ~new_n51450_ & ~new_n51451_;
  assign new_n51453_ = ~new_n51122_ & ~new_n51452_;
  assign new_n51454_ = ~new_n50661_ & ~new_n51121_;
  assign new_n51455_ = ~new_n51120_ & new_n51454_;
  assign new_n51456_ = ~new_n51453_ & ~new_n51455_;
  assign new_n51457_ = ~\b[21]  & ~new_n51456_;
  assign new_n51458_ = ~new_n50680_ & new_n50922_;
  assign new_n51459_ = ~new_n50918_ & new_n51458_;
  assign new_n51460_ = ~new_n50919_ & ~new_n50922_;
  assign new_n51461_ = ~new_n51459_ & ~new_n51460_;
  assign new_n51462_ = ~new_n51122_ & ~new_n51461_;
  assign new_n51463_ = ~new_n50670_ & ~new_n51121_;
  assign new_n51464_ = ~new_n51120_ & new_n51463_;
  assign new_n51465_ = ~new_n51462_ & ~new_n51464_;
  assign new_n51466_ = ~\b[20]  & ~new_n51465_;
  assign new_n51467_ = ~new_n50689_ & new_n50917_;
  assign new_n51468_ = ~new_n50913_ & new_n51467_;
  assign new_n51469_ = ~new_n50914_ & ~new_n50917_;
  assign new_n51470_ = ~new_n51468_ & ~new_n51469_;
  assign new_n51471_ = ~new_n51122_ & ~new_n51470_;
  assign new_n51472_ = ~new_n50679_ & ~new_n51121_;
  assign new_n51473_ = ~new_n51120_ & new_n51472_;
  assign new_n51474_ = ~new_n51471_ & ~new_n51473_;
  assign new_n51475_ = ~\b[19]  & ~new_n51474_;
  assign new_n51476_ = ~new_n50698_ & new_n50912_;
  assign new_n51477_ = ~new_n50908_ & new_n51476_;
  assign new_n51478_ = ~new_n50909_ & ~new_n50912_;
  assign new_n51479_ = ~new_n51477_ & ~new_n51478_;
  assign new_n51480_ = ~new_n51122_ & ~new_n51479_;
  assign new_n51481_ = ~new_n50688_ & ~new_n51121_;
  assign new_n51482_ = ~new_n51120_ & new_n51481_;
  assign new_n51483_ = ~new_n51480_ & ~new_n51482_;
  assign new_n51484_ = ~\b[18]  & ~new_n51483_;
  assign new_n51485_ = ~new_n50707_ & new_n50907_;
  assign new_n51486_ = ~new_n50903_ & new_n51485_;
  assign new_n51487_ = ~new_n50904_ & ~new_n50907_;
  assign new_n51488_ = ~new_n51486_ & ~new_n51487_;
  assign new_n51489_ = ~new_n51122_ & ~new_n51488_;
  assign new_n51490_ = ~new_n50697_ & ~new_n51121_;
  assign new_n51491_ = ~new_n51120_ & new_n51490_;
  assign new_n51492_ = ~new_n51489_ & ~new_n51491_;
  assign new_n51493_ = ~\b[17]  & ~new_n51492_;
  assign new_n51494_ = ~new_n50716_ & new_n50902_;
  assign new_n51495_ = ~new_n50898_ & new_n51494_;
  assign new_n51496_ = ~new_n50899_ & ~new_n50902_;
  assign new_n51497_ = ~new_n51495_ & ~new_n51496_;
  assign new_n51498_ = ~new_n51122_ & ~new_n51497_;
  assign new_n51499_ = ~new_n50706_ & ~new_n51121_;
  assign new_n51500_ = ~new_n51120_ & new_n51499_;
  assign new_n51501_ = ~new_n51498_ & ~new_n51500_;
  assign new_n51502_ = ~\b[16]  & ~new_n51501_;
  assign new_n51503_ = ~new_n50725_ & new_n50897_;
  assign new_n51504_ = ~new_n50893_ & new_n51503_;
  assign new_n51505_ = ~new_n50894_ & ~new_n50897_;
  assign new_n51506_ = ~new_n51504_ & ~new_n51505_;
  assign new_n51507_ = ~new_n51122_ & ~new_n51506_;
  assign new_n51508_ = ~new_n50715_ & ~new_n51121_;
  assign new_n51509_ = ~new_n51120_ & new_n51508_;
  assign new_n51510_ = ~new_n51507_ & ~new_n51509_;
  assign new_n51511_ = ~\b[15]  & ~new_n51510_;
  assign new_n51512_ = ~new_n50734_ & new_n50892_;
  assign new_n51513_ = ~new_n50888_ & new_n51512_;
  assign new_n51514_ = ~new_n50889_ & ~new_n50892_;
  assign new_n51515_ = ~new_n51513_ & ~new_n51514_;
  assign new_n51516_ = ~new_n51122_ & ~new_n51515_;
  assign new_n51517_ = ~new_n50724_ & ~new_n51121_;
  assign new_n51518_ = ~new_n51120_ & new_n51517_;
  assign new_n51519_ = ~new_n51516_ & ~new_n51518_;
  assign new_n51520_ = ~\b[14]  & ~new_n51519_;
  assign new_n51521_ = ~new_n50743_ & new_n50887_;
  assign new_n51522_ = ~new_n50883_ & new_n51521_;
  assign new_n51523_ = ~new_n50884_ & ~new_n50887_;
  assign new_n51524_ = ~new_n51522_ & ~new_n51523_;
  assign new_n51525_ = ~new_n51122_ & ~new_n51524_;
  assign new_n51526_ = ~new_n50733_ & ~new_n51121_;
  assign new_n51527_ = ~new_n51120_ & new_n51526_;
  assign new_n51528_ = ~new_n51525_ & ~new_n51527_;
  assign new_n51529_ = ~\b[13]  & ~new_n51528_;
  assign new_n51530_ = ~new_n50752_ & new_n50882_;
  assign new_n51531_ = ~new_n50878_ & new_n51530_;
  assign new_n51532_ = ~new_n50879_ & ~new_n50882_;
  assign new_n51533_ = ~new_n51531_ & ~new_n51532_;
  assign new_n51534_ = ~new_n51122_ & ~new_n51533_;
  assign new_n51535_ = ~new_n50742_ & ~new_n51121_;
  assign new_n51536_ = ~new_n51120_ & new_n51535_;
  assign new_n51537_ = ~new_n51534_ & ~new_n51536_;
  assign new_n51538_ = ~\b[12]  & ~new_n51537_;
  assign new_n51539_ = ~new_n50761_ & new_n50877_;
  assign new_n51540_ = ~new_n50873_ & new_n51539_;
  assign new_n51541_ = ~new_n50874_ & ~new_n50877_;
  assign new_n51542_ = ~new_n51540_ & ~new_n51541_;
  assign new_n51543_ = ~new_n51122_ & ~new_n51542_;
  assign new_n51544_ = ~new_n50751_ & ~new_n51121_;
  assign new_n51545_ = ~new_n51120_ & new_n51544_;
  assign new_n51546_ = ~new_n51543_ & ~new_n51545_;
  assign new_n51547_ = ~\b[11]  & ~new_n51546_;
  assign new_n51548_ = ~new_n50770_ & new_n50872_;
  assign new_n51549_ = ~new_n50868_ & new_n51548_;
  assign new_n51550_ = ~new_n50869_ & ~new_n50872_;
  assign new_n51551_ = ~new_n51549_ & ~new_n51550_;
  assign new_n51552_ = ~new_n51122_ & ~new_n51551_;
  assign new_n51553_ = ~new_n50760_ & ~new_n51121_;
  assign new_n51554_ = ~new_n51120_ & new_n51553_;
  assign new_n51555_ = ~new_n51552_ & ~new_n51554_;
  assign new_n51556_ = ~\b[10]  & ~new_n51555_;
  assign new_n51557_ = ~new_n50779_ & new_n50867_;
  assign new_n51558_ = ~new_n50863_ & new_n51557_;
  assign new_n51559_ = ~new_n50864_ & ~new_n50867_;
  assign new_n51560_ = ~new_n51558_ & ~new_n51559_;
  assign new_n51561_ = ~new_n51122_ & ~new_n51560_;
  assign new_n51562_ = ~new_n50769_ & ~new_n51121_;
  assign new_n51563_ = ~new_n51120_ & new_n51562_;
  assign new_n51564_ = ~new_n51561_ & ~new_n51563_;
  assign new_n51565_ = ~\b[9]  & ~new_n51564_;
  assign new_n51566_ = ~new_n50788_ & new_n50862_;
  assign new_n51567_ = ~new_n50858_ & new_n51566_;
  assign new_n51568_ = ~new_n50859_ & ~new_n50862_;
  assign new_n51569_ = ~new_n51567_ & ~new_n51568_;
  assign new_n51570_ = ~new_n51122_ & ~new_n51569_;
  assign new_n51571_ = ~new_n50778_ & ~new_n51121_;
  assign new_n51572_ = ~new_n51120_ & new_n51571_;
  assign new_n51573_ = ~new_n51570_ & ~new_n51572_;
  assign new_n51574_ = ~\b[8]  & ~new_n51573_;
  assign new_n51575_ = ~new_n50797_ & new_n50857_;
  assign new_n51576_ = ~new_n50853_ & new_n51575_;
  assign new_n51577_ = ~new_n50854_ & ~new_n50857_;
  assign new_n51578_ = ~new_n51576_ & ~new_n51577_;
  assign new_n51579_ = ~new_n51122_ & ~new_n51578_;
  assign new_n51580_ = ~new_n50787_ & ~new_n51121_;
  assign new_n51581_ = ~new_n51120_ & new_n51580_;
  assign new_n51582_ = ~new_n51579_ & ~new_n51581_;
  assign new_n51583_ = ~\b[7]  & ~new_n51582_;
  assign new_n51584_ = ~new_n50806_ & new_n50852_;
  assign new_n51585_ = ~new_n50848_ & new_n51584_;
  assign new_n51586_ = ~new_n50849_ & ~new_n50852_;
  assign new_n51587_ = ~new_n51585_ & ~new_n51586_;
  assign new_n51588_ = ~new_n51122_ & ~new_n51587_;
  assign new_n51589_ = ~new_n50796_ & ~new_n51121_;
  assign new_n51590_ = ~new_n51120_ & new_n51589_;
  assign new_n51591_ = ~new_n51588_ & ~new_n51590_;
  assign new_n51592_ = ~\b[6]  & ~new_n51591_;
  assign new_n51593_ = ~new_n50815_ & new_n50847_;
  assign new_n51594_ = ~new_n50843_ & new_n51593_;
  assign new_n51595_ = ~new_n50844_ & ~new_n50847_;
  assign new_n51596_ = ~new_n51594_ & ~new_n51595_;
  assign new_n51597_ = ~new_n51122_ & ~new_n51596_;
  assign new_n51598_ = ~new_n50805_ & ~new_n51121_;
  assign new_n51599_ = ~new_n51120_ & new_n51598_;
  assign new_n51600_ = ~new_n51597_ & ~new_n51599_;
  assign new_n51601_ = ~\b[5]  & ~new_n51600_;
  assign new_n51602_ = ~new_n50823_ & new_n50842_;
  assign new_n51603_ = ~new_n50838_ & new_n51602_;
  assign new_n51604_ = ~new_n50839_ & ~new_n50842_;
  assign new_n51605_ = ~new_n51603_ & ~new_n51604_;
  assign new_n51606_ = ~new_n51122_ & ~new_n51605_;
  assign new_n51607_ = ~new_n50814_ & ~new_n51121_;
  assign new_n51608_ = ~new_n51120_ & new_n51607_;
  assign new_n51609_ = ~new_n51606_ & ~new_n51608_;
  assign new_n51610_ = ~\b[4]  & ~new_n51609_;
  assign new_n51611_ = ~new_n50833_ & new_n50837_;
  assign new_n51612_ = ~new_n50832_ & new_n51611_;
  assign new_n51613_ = ~new_n50834_ & ~new_n50837_;
  assign new_n51614_ = ~new_n51612_ & ~new_n51613_;
  assign new_n51615_ = ~new_n51122_ & ~new_n51614_;
  assign new_n51616_ = ~new_n50822_ & ~new_n51121_;
  assign new_n51617_ = ~new_n51120_ & new_n51616_;
  assign new_n51618_ = ~new_n51615_ & ~new_n51617_;
  assign new_n51619_ = ~\b[3]  & ~new_n51618_;
  assign new_n51620_ = new_n22806_ & ~new_n50830_;
  assign new_n51621_ = ~new_n50828_ & new_n51620_;
  assign new_n51622_ = ~new_n50832_ & ~new_n51621_;
  assign new_n51623_ = ~new_n51122_ & new_n51622_;
  assign new_n51624_ = ~new_n50827_ & ~new_n51121_;
  assign new_n51625_ = ~new_n51120_ & new_n51624_;
  assign new_n51626_ = ~new_n51623_ & ~new_n51625_;
  assign new_n51627_ = ~\b[2]  & ~new_n51626_;
  assign new_n51628_ = \b[0]  & ~new_n51122_;
  assign new_n51629_ = \a[7]  & ~new_n51628_;
  assign new_n51630_ = new_n22806_ & ~new_n51122_;
  assign new_n51631_ = ~new_n51629_ & ~new_n51630_;
  assign new_n51632_ = \b[1]  & ~new_n51631_;
  assign new_n51633_ = ~\b[1]  & ~new_n51630_;
  assign new_n51634_ = ~new_n51629_ & new_n51633_;
  assign new_n51635_ = ~new_n51632_ & ~new_n51634_;
  assign new_n51636_ = ~new_n23611_ & ~new_n51635_;
  assign new_n51637_ = ~\b[1]  & ~new_n51631_;
  assign new_n51638_ = ~new_n51636_ & ~new_n51637_;
  assign new_n51639_ = \b[2]  & ~new_n51625_;
  assign new_n51640_ = ~new_n51623_ & new_n51639_;
  assign new_n51641_ = ~new_n51627_ & ~new_n51640_;
  assign new_n51642_ = ~new_n51638_ & new_n51641_;
  assign new_n51643_ = ~new_n51627_ & ~new_n51642_;
  assign new_n51644_ = \b[3]  & ~new_n51617_;
  assign new_n51645_ = ~new_n51615_ & new_n51644_;
  assign new_n51646_ = ~new_n51619_ & ~new_n51645_;
  assign new_n51647_ = ~new_n51643_ & new_n51646_;
  assign new_n51648_ = ~new_n51619_ & ~new_n51647_;
  assign new_n51649_ = \b[4]  & ~new_n51608_;
  assign new_n51650_ = ~new_n51606_ & new_n51649_;
  assign new_n51651_ = ~new_n51610_ & ~new_n51650_;
  assign new_n51652_ = ~new_n51648_ & new_n51651_;
  assign new_n51653_ = ~new_n51610_ & ~new_n51652_;
  assign new_n51654_ = \b[5]  & ~new_n51599_;
  assign new_n51655_ = ~new_n51597_ & new_n51654_;
  assign new_n51656_ = ~new_n51601_ & ~new_n51655_;
  assign new_n51657_ = ~new_n51653_ & new_n51656_;
  assign new_n51658_ = ~new_n51601_ & ~new_n51657_;
  assign new_n51659_ = \b[6]  & ~new_n51590_;
  assign new_n51660_ = ~new_n51588_ & new_n51659_;
  assign new_n51661_ = ~new_n51592_ & ~new_n51660_;
  assign new_n51662_ = ~new_n51658_ & new_n51661_;
  assign new_n51663_ = ~new_n51592_ & ~new_n51662_;
  assign new_n51664_ = \b[7]  & ~new_n51581_;
  assign new_n51665_ = ~new_n51579_ & new_n51664_;
  assign new_n51666_ = ~new_n51583_ & ~new_n51665_;
  assign new_n51667_ = ~new_n51663_ & new_n51666_;
  assign new_n51668_ = ~new_n51583_ & ~new_n51667_;
  assign new_n51669_ = \b[8]  & ~new_n51572_;
  assign new_n51670_ = ~new_n51570_ & new_n51669_;
  assign new_n51671_ = ~new_n51574_ & ~new_n51670_;
  assign new_n51672_ = ~new_n51668_ & new_n51671_;
  assign new_n51673_ = ~new_n51574_ & ~new_n51672_;
  assign new_n51674_ = \b[9]  & ~new_n51563_;
  assign new_n51675_ = ~new_n51561_ & new_n51674_;
  assign new_n51676_ = ~new_n51565_ & ~new_n51675_;
  assign new_n51677_ = ~new_n51673_ & new_n51676_;
  assign new_n51678_ = ~new_n51565_ & ~new_n51677_;
  assign new_n51679_ = \b[10]  & ~new_n51554_;
  assign new_n51680_ = ~new_n51552_ & new_n51679_;
  assign new_n51681_ = ~new_n51556_ & ~new_n51680_;
  assign new_n51682_ = ~new_n51678_ & new_n51681_;
  assign new_n51683_ = ~new_n51556_ & ~new_n51682_;
  assign new_n51684_ = \b[11]  & ~new_n51545_;
  assign new_n51685_ = ~new_n51543_ & new_n51684_;
  assign new_n51686_ = ~new_n51547_ & ~new_n51685_;
  assign new_n51687_ = ~new_n51683_ & new_n51686_;
  assign new_n51688_ = ~new_n51547_ & ~new_n51687_;
  assign new_n51689_ = \b[12]  & ~new_n51536_;
  assign new_n51690_ = ~new_n51534_ & new_n51689_;
  assign new_n51691_ = ~new_n51538_ & ~new_n51690_;
  assign new_n51692_ = ~new_n51688_ & new_n51691_;
  assign new_n51693_ = ~new_n51538_ & ~new_n51692_;
  assign new_n51694_ = \b[13]  & ~new_n51527_;
  assign new_n51695_ = ~new_n51525_ & new_n51694_;
  assign new_n51696_ = ~new_n51529_ & ~new_n51695_;
  assign new_n51697_ = ~new_n51693_ & new_n51696_;
  assign new_n51698_ = ~new_n51529_ & ~new_n51697_;
  assign new_n51699_ = \b[14]  & ~new_n51518_;
  assign new_n51700_ = ~new_n51516_ & new_n51699_;
  assign new_n51701_ = ~new_n51520_ & ~new_n51700_;
  assign new_n51702_ = ~new_n51698_ & new_n51701_;
  assign new_n51703_ = ~new_n51520_ & ~new_n51702_;
  assign new_n51704_ = \b[15]  & ~new_n51509_;
  assign new_n51705_ = ~new_n51507_ & new_n51704_;
  assign new_n51706_ = ~new_n51511_ & ~new_n51705_;
  assign new_n51707_ = ~new_n51703_ & new_n51706_;
  assign new_n51708_ = ~new_n51511_ & ~new_n51707_;
  assign new_n51709_ = \b[16]  & ~new_n51500_;
  assign new_n51710_ = ~new_n51498_ & new_n51709_;
  assign new_n51711_ = ~new_n51502_ & ~new_n51710_;
  assign new_n51712_ = ~new_n51708_ & new_n51711_;
  assign new_n51713_ = ~new_n51502_ & ~new_n51712_;
  assign new_n51714_ = \b[17]  & ~new_n51491_;
  assign new_n51715_ = ~new_n51489_ & new_n51714_;
  assign new_n51716_ = ~new_n51493_ & ~new_n51715_;
  assign new_n51717_ = ~new_n51713_ & new_n51716_;
  assign new_n51718_ = ~new_n51493_ & ~new_n51717_;
  assign new_n51719_ = \b[18]  & ~new_n51482_;
  assign new_n51720_ = ~new_n51480_ & new_n51719_;
  assign new_n51721_ = ~new_n51484_ & ~new_n51720_;
  assign new_n51722_ = ~new_n51718_ & new_n51721_;
  assign new_n51723_ = ~new_n51484_ & ~new_n51722_;
  assign new_n51724_ = \b[19]  & ~new_n51473_;
  assign new_n51725_ = ~new_n51471_ & new_n51724_;
  assign new_n51726_ = ~new_n51475_ & ~new_n51725_;
  assign new_n51727_ = ~new_n51723_ & new_n51726_;
  assign new_n51728_ = ~new_n51475_ & ~new_n51727_;
  assign new_n51729_ = \b[20]  & ~new_n51464_;
  assign new_n51730_ = ~new_n51462_ & new_n51729_;
  assign new_n51731_ = ~new_n51466_ & ~new_n51730_;
  assign new_n51732_ = ~new_n51728_ & new_n51731_;
  assign new_n51733_ = ~new_n51466_ & ~new_n51732_;
  assign new_n51734_ = \b[21]  & ~new_n51455_;
  assign new_n51735_ = ~new_n51453_ & new_n51734_;
  assign new_n51736_ = ~new_n51457_ & ~new_n51735_;
  assign new_n51737_ = ~new_n51733_ & new_n51736_;
  assign new_n51738_ = ~new_n51457_ & ~new_n51737_;
  assign new_n51739_ = \b[22]  & ~new_n51446_;
  assign new_n51740_ = ~new_n51444_ & new_n51739_;
  assign new_n51741_ = ~new_n51448_ & ~new_n51740_;
  assign new_n51742_ = ~new_n51738_ & new_n51741_;
  assign new_n51743_ = ~new_n51448_ & ~new_n51742_;
  assign new_n51744_ = \b[23]  & ~new_n51437_;
  assign new_n51745_ = ~new_n51435_ & new_n51744_;
  assign new_n51746_ = ~new_n51439_ & ~new_n51745_;
  assign new_n51747_ = ~new_n51743_ & new_n51746_;
  assign new_n51748_ = ~new_n51439_ & ~new_n51747_;
  assign new_n51749_ = \b[24]  & ~new_n51428_;
  assign new_n51750_ = ~new_n51426_ & new_n51749_;
  assign new_n51751_ = ~new_n51430_ & ~new_n51750_;
  assign new_n51752_ = ~new_n51748_ & new_n51751_;
  assign new_n51753_ = ~new_n51430_ & ~new_n51752_;
  assign new_n51754_ = \b[25]  & ~new_n51419_;
  assign new_n51755_ = ~new_n51417_ & new_n51754_;
  assign new_n51756_ = ~new_n51421_ & ~new_n51755_;
  assign new_n51757_ = ~new_n51753_ & new_n51756_;
  assign new_n51758_ = ~new_n51421_ & ~new_n51757_;
  assign new_n51759_ = \b[26]  & ~new_n51410_;
  assign new_n51760_ = ~new_n51408_ & new_n51759_;
  assign new_n51761_ = ~new_n51412_ & ~new_n51760_;
  assign new_n51762_ = ~new_n51758_ & new_n51761_;
  assign new_n51763_ = ~new_n51412_ & ~new_n51762_;
  assign new_n51764_ = \b[27]  & ~new_n51401_;
  assign new_n51765_ = ~new_n51399_ & new_n51764_;
  assign new_n51766_ = ~new_n51403_ & ~new_n51765_;
  assign new_n51767_ = ~new_n51763_ & new_n51766_;
  assign new_n51768_ = ~new_n51403_ & ~new_n51767_;
  assign new_n51769_ = \b[28]  & ~new_n51392_;
  assign new_n51770_ = ~new_n51390_ & new_n51769_;
  assign new_n51771_ = ~new_n51394_ & ~new_n51770_;
  assign new_n51772_ = ~new_n51768_ & new_n51771_;
  assign new_n51773_ = ~new_n51394_ & ~new_n51772_;
  assign new_n51774_ = \b[29]  & ~new_n51383_;
  assign new_n51775_ = ~new_n51381_ & new_n51774_;
  assign new_n51776_ = ~new_n51385_ & ~new_n51775_;
  assign new_n51777_ = ~new_n51773_ & new_n51776_;
  assign new_n51778_ = ~new_n51385_ & ~new_n51777_;
  assign new_n51779_ = \b[30]  & ~new_n51374_;
  assign new_n51780_ = ~new_n51372_ & new_n51779_;
  assign new_n51781_ = ~new_n51376_ & ~new_n51780_;
  assign new_n51782_ = ~new_n51778_ & new_n51781_;
  assign new_n51783_ = ~new_n51376_ & ~new_n51782_;
  assign new_n51784_ = \b[31]  & ~new_n51365_;
  assign new_n51785_ = ~new_n51363_ & new_n51784_;
  assign new_n51786_ = ~new_n51367_ & ~new_n51785_;
  assign new_n51787_ = ~new_n51783_ & new_n51786_;
  assign new_n51788_ = ~new_n51367_ & ~new_n51787_;
  assign new_n51789_ = \b[32]  & ~new_n51356_;
  assign new_n51790_ = ~new_n51354_ & new_n51789_;
  assign new_n51791_ = ~new_n51358_ & ~new_n51790_;
  assign new_n51792_ = ~new_n51788_ & new_n51791_;
  assign new_n51793_ = ~new_n51358_ & ~new_n51792_;
  assign new_n51794_ = \b[33]  & ~new_n51347_;
  assign new_n51795_ = ~new_n51345_ & new_n51794_;
  assign new_n51796_ = ~new_n51349_ & ~new_n51795_;
  assign new_n51797_ = ~new_n51793_ & new_n51796_;
  assign new_n51798_ = ~new_n51349_ & ~new_n51797_;
  assign new_n51799_ = \b[34]  & ~new_n51338_;
  assign new_n51800_ = ~new_n51336_ & new_n51799_;
  assign new_n51801_ = ~new_n51340_ & ~new_n51800_;
  assign new_n51802_ = ~new_n51798_ & new_n51801_;
  assign new_n51803_ = ~new_n51340_ & ~new_n51802_;
  assign new_n51804_ = \b[35]  & ~new_n51329_;
  assign new_n51805_ = ~new_n51327_ & new_n51804_;
  assign new_n51806_ = ~new_n51331_ & ~new_n51805_;
  assign new_n51807_ = ~new_n51803_ & new_n51806_;
  assign new_n51808_ = ~new_n51331_ & ~new_n51807_;
  assign new_n51809_ = \b[36]  & ~new_n51320_;
  assign new_n51810_ = ~new_n51318_ & new_n51809_;
  assign new_n51811_ = ~new_n51322_ & ~new_n51810_;
  assign new_n51812_ = ~new_n51808_ & new_n51811_;
  assign new_n51813_ = ~new_n51322_ & ~new_n51812_;
  assign new_n51814_ = \b[37]  & ~new_n51311_;
  assign new_n51815_ = ~new_n51309_ & new_n51814_;
  assign new_n51816_ = ~new_n51313_ & ~new_n51815_;
  assign new_n51817_ = ~new_n51813_ & new_n51816_;
  assign new_n51818_ = ~new_n51313_ & ~new_n51817_;
  assign new_n51819_ = \b[38]  & ~new_n51302_;
  assign new_n51820_ = ~new_n51300_ & new_n51819_;
  assign new_n51821_ = ~new_n51304_ & ~new_n51820_;
  assign new_n51822_ = ~new_n51818_ & new_n51821_;
  assign new_n51823_ = ~new_n51304_ & ~new_n51822_;
  assign new_n51824_ = \b[39]  & ~new_n51293_;
  assign new_n51825_ = ~new_n51291_ & new_n51824_;
  assign new_n51826_ = ~new_n51295_ & ~new_n51825_;
  assign new_n51827_ = ~new_n51823_ & new_n51826_;
  assign new_n51828_ = ~new_n51295_ & ~new_n51827_;
  assign new_n51829_ = \b[40]  & ~new_n51284_;
  assign new_n51830_ = ~new_n51282_ & new_n51829_;
  assign new_n51831_ = ~new_n51286_ & ~new_n51830_;
  assign new_n51832_ = ~new_n51828_ & new_n51831_;
  assign new_n51833_ = ~new_n51286_ & ~new_n51832_;
  assign new_n51834_ = \b[41]  & ~new_n51275_;
  assign new_n51835_ = ~new_n51273_ & new_n51834_;
  assign new_n51836_ = ~new_n51277_ & ~new_n51835_;
  assign new_n51837_ = ~new_n51833_ & new_n51836_;
  assign new_n51838_ = ~new_n51277_ & ~new_n51837_;
  assign new_n51839_ = \b[42]  & ~new_n51266_;
  assign new_n51840_ = ~new_n51264_ & new_n51839_;
  assign new_n51841_ = ~new_n51268_ & ~new_n51840_;
  assign new_n51842_ = ~new_n51838_ & new_n51841_;
  assign new_n51843_ = ~new_n51268_ & ~new_n51842_;
  assign new_n51844_ = \b[43]  & ~new_n51257_;
  assign new_n51845_ = ~new_n51255_ & new_n51844_;
  assign new_n51846_ = ~new_n51259_ & ~new_n51845_;
  assign new_n51847_ = ~new_n51843_ & new_n51846_;
  assign new_n51848_ = ~new_n51259_ & ~new_n51847_;
  assign new_n51849_ = \b[44]  & ~new_n51248_;
  assign new_n51850_ = ~new_n51246_ & new_n51849_;
  assign new_n51851_ = ~new_n51250_ & ~new_n51850_;
  assign new_n51852_ = ~new_n51848_ & new_n51851_;
  assign new_n51853_ = ~new_n51250_ & ~new_n51852_;
  assign new_n51854_ = \b[45]  & ~new_n51239_;
  assign new_n51855_ = ~new_n51237_ & new_n51854_;
  assign new_n51856_ = ~new_n51241_ & ~new_n51855_;
  assign new_n51857_ = ~new_n51853_ & new_n51856_;
  assign new_n51858_ = ~new_n51241_ & ~new_n51857_;
  assign new_n51859_ = \b[46]  & ~new_n51230_;
  assign new_n51860_ = ~new_n51228_ & new_n51859_;
  assign new_n51861_ = ~new_n51232_ & ~new_n51860_;
  assign new_n51862_ = ~new_n51858_ & new_n51861_;
  assign new_n51863_ = ~new_n51232_ & ~new_n51862_;
  assign new_n51864_ = \b[47]  & ~new_n51221_;
  assign new_n51865_ = ~new_n51219_ & new_n51864_;
  assign new_n51866_ = ~new_n51223_ & ~new_n51865_;
  assign new_n51867_ = ~new_n51863_ & new_n51866_;
  assign new_n51868_ = ~new_n51223_ & ~new_n51867_;
  assign new_n51869_ = \b[48]  & ~new_n51212_;
  assign new_n51870_ = ~new_n51210_ & new_n51869_;
  assign new_n51871_ = ~new_n51214_ & ~new_n51870_;
  assign new_n51872_ = ~new_n51868_ & new_n51871_;
  assign new_n51873_ = ~new_n51214_ & ~new_n51872_;
  assign new_n51874_ = \b[49]  & ~new_n51203_;
  assign new_n51875_ = ~new_n51201_ & new_n51874_;
  assign new_n51876_ = ~new_n51205_ & ~new_n51875_;
  assign new_n51877_ = ~new_n51873_ & new_n51876_;
  assign new_n51878_ = ~new_n51205_ & ~new_n51877_;
  assign new_n51879_ = \b[50]  & ~new_n51194_;
  assign new_n51880_ = ~new_n51192_ & new_n51879_;
  assign new_n51881_ = ~new_n51196_ & ~new_n51880_;
  assign new_n51882_ = ~new_n51878_ & new_n51881_;
  assign new_n51883_ = ~new_n51196_ & ~new_n51882_;
  assign new_n51884_ = \b[51]  & ~new_n51185_;
  assign new_n51885_ = ~new_n51183_ & new_n51884_;
  assign new_n51886_ = ~new_n51187_ & ~new_n51885_;
  assign new_n51887_ = ~new_n51883_ & new_n51886_;
  assign new_n51888_ = ~new_n51187_ & ~new_n51887_;
  assign new_n51889_ = \b[52]  & ~new_n51176_;
  assign new_n51890_ = ~new_n51174_ & new_n51889_;
  assign new_n51891_ = ~new_n51178_ & ~new_n51890_;
  assign new_n51892_ = ~new_n51888_ & new_n51891_;
  assign new_n51893_ = ~new_n51178_ & ~new_n51892_;
  assign new_n51894_ = \b[53]  & ~new_n51167_;
  assign new_n51895_ = ~new_n51165_ & new_n51894_;
  assign new_n51896_ = ~new_n51169_ & ~new_n51895_;
  assign new_n51897_ = ~new_n51893_ & new_n51896_;
  assign new_n51898_ = ~new_n51169_ & ~new_n51897_;
  assign new_n51899_ = \b[54]  & ~new_n51158_;
  assign new_n51900_ = ~new_n51156_ & new_n51899_;
  assign new_n51901_ = ~new_n51160_ & ~new_n51900_;
  assign new_n51902_ = ~new_n51898_ & new_n51901_;
  assign new_n51903_ = ~new_n51160_ & ~new_n51902_;
  assign new_n51904_ = \b[55]  & ~new_n51149_;
  assign new_n51905_ = ~new_n51147_ & new_n51904_;
  assign new_n51906_ = ~new_n51151_ & ~new_n51905_;
  assign new_n51907_ = ~new_n51903_ & new_n51906_;
  assign new_n51908_ = ~new_n51151_ & ~new_n51907_;
  assign new_n51909_ = \b[56]  & ~new_n51129_;
  assign new_n51910_ = ~new_n51127_ & new_n51909_;
  assign new_n51911_ = ~new_n51142_ & ~new_n51910_;
  assign new_n51912_ = ~new_n51908_ & new_n51911_;
  assign new_n51913_ = ~new_n51142_ & ~new_n51912_;
  assign new_n51914_ = \b[57]  & ~new_n51139_;
  assign new_n51915_ = ~new_n51137_ & new_n51914_;
  assign new_n51916_ = ~new_n51141_ & ~new_n51915_;
  assign new_n51917_ = ~new_n51913_ & new_n51916_;
  assign new_n51918_ = ~new_n51141_ & ~new_n51917_;
  assign new_n51919_ = new_n23895_ & ~new_n51918_;
  assign new_n51920_ = ~new_n51130_ & ~new_n51919_;
  assign new_n51921_ = ~new_n51151_ & new_n51911_;
  assign new_n51922_ = ~new_n51907_ & new_n51921_;
  assign new_n51923_ = ~new_n51908_ & ~new_n51911_;
  assign new_n51924_ = ~new_n51922_ & ~new_n51923_;
  assign new_n51925_ = new_n23895_ & ~new_n51924_;
  assign new_n51926_ = ~new_n51918_ & new_n51925_;
  assign new_n51927_ = ~new_n51920_ & ~new_n51926_;
  assign new_n51928_ = ~\b[57]  & ~new_n51927_;
  assign new_n51929_ = ~new_n51150_ & ~new_n51919_;
  assign new_n51930_ = ~new_n51160_ & new_n51906_;
  assign new_n51931_ = ~new_n51902_ & new_n51930_;
  assign new_n51932_ = ~new_n51903_ & ~new_n51906_;
  assign new_n51933_ = ~new_n51931_ & ~new_n51932_;
  assign new_n51934_ = new_n23895_ & ~new_n51933_;
  assign new_n51935_ = ~new_n51918_ & new_n51934_;
  assign new_n51936_ = ~new_n51929_ & ~new_n51935_;
  assign new_n51937_ = ~\b[56]  & ~new_n51936_;
  assign new_n51938_ = ~new_n51159_ & ~new_n51919_;
  assign new_n51939_ = ~new_n51169_ & new_n51901_;
  assign new_n51940_ = ~new_n51897_ & new_n51939_;
  assign new_n51941_ = ~new_n51898_ & ~new_n51901_;
  assign new_n51942_ = ~new_n51940_ & ~new_n51941_;
  assign new_n51943_ = new_n23895_ & ~new_n51942_;
  assign new_n51944_ = ~new_n51918_ & new_n51943_;
  assign new_n51945_ = ~new_n51938_ & ~new_n51944_;
  assign new_n51946_ = ~\b[55]  & ~new_n51945_;
  assign new_n51947_ = ~new_n51168_ & ~new_n51919_;
  assign new_n51948_ = ~new_n51178_ & new_n51896_;
  assign new_n51949_ = ~new_n51892_ & new_n51948_;
  assign new_n51950_ = ~new_n51893_ & ~new_n51896_;
  assign new_n51951_ = ~new_n51949_ & ~new_n51950_;
  assign new_n51952_ = new_n23895_ & ~new_n51951_;
  assign new_n51953_ = ~new_n51918_ & new_n51952_;
  assign new_n51954_ = ~new_n51947_ & ~new_n51953_;
  assign new_n51955_ = ~\b[54]  & ~new_n51954_;
  assign new_n51956_ = ~new_n51177_ & ~new_n51919_;
  assign new_n51957_ = ~new_n51187_ & new_n51891_;
  assign new_n51958_ = ~new_n51887_ & new_n51957_;
  assign new_n51959_ = ~new_n51888_ & ~new_n51891_;
  assign new_n51960_ = ~new_n51958_ & ~new_n51959_;
  assign new_n51961_ = new_n23895_ & ~new_n51960_;
  assign new_n51962_ = ~new_n51918_ & new_n51961_;
  assign new_n51963_ = ~new_n51956_ & ~new_n51962_;
  assign new_n51964_ = ~\b[53]  & ~new_n51963_;
  assign new_n51965_ = ~new_n51186_ & ~new_n51919_;
  assign new_n51966_ = ~new_n51196_ & new_n51886_;
  assign new_n51967_ = ~new_n51882_ & new_n51966_;
  assign new_n51968_ = ~new_n51883_ & ~new_n51886_;
  assign new_n51969_ = ~new_n51967_ & ~new_n51968_;
  assign new_n51970_ = new_n23895_ & ~new_n51969_;
  assign new_n51971_ = ~new_n51918_ & new_n51970_;
  assign new_n51972_ = ~new_n51965_ & ~new_n51971_;
  assign new_n51973_ = ~\b[52]  & ~new_n51972_;
  assign new_n51974_ = ~new_n51195_ & ~new_n51919_;
  assign new_n51975_ = ~new_n51205_ & new_n51881_;
  assign new_n51976_ = ~new_n51877_ & new_n51975_;
  assign new_n51977_ = ~new_n51878_ & ~new_n51881_;
  assign new_n51978_ = ~new_n51976_ & ~new_n51977_;
  assign new_n51979_ = new_n23895_ & ~new_n51978_;
  assign new_n51980_ = ~new_n51918_ & new_n51979_;
  assign new_n51981_ = ~new_n51974_ & ~new_n51980_;
  assign new_n51982_ = ~\b[51]  & ~new_n51981_;
  assign new_n51983_ = ~new_n51204_ & ~new_n51919_;
  assign new_n51984_ = ~new_n51214_ & new_n51876_;
  assign new_n51985_ = ~new_n51872_ & new_n51984_;
  assign new_n51986_ = ~new_n51873_ & ~new_n51876_;
  assign new_n51987_ = ~new_n51985_ & ~new_n51986_;
  assign new_n51988_ = new_n23895_ & ~new_n51987_;
  assign new_n51989_ = ~new_n51918_ & new_n51988_;
  assign new_n51990_ = ~new_n51983_ & ~new_n51989_;
  assign new_n51991_ = ~\b[50]  & ~new_n51990_;
  assign new_n51992_ = ~new_n51213_ & ~new_n51919_;
  assign new_n51993_ = ~new_n51223_ & new_n51871_;
  assign new_n51994_ = ~new_n51867_ & new_n51993_;
  assign new_n51995_ = ~new_n51868_ & ~new_n51871_;
  assign new_n51996_ = ~new_n51994_ & ~new_n51995_;
  assign new_n51997_ = new_n23895_ & ~new_n51996_;
  assign new_n51998_ = ~new_n51918_ & new_n51997_;
  assign new_n51999_ = ~new_n51992_ & ~new_n51998_;
  assign new_n52000_ = ~\b[49]  & ~new_n51999_;
  assign new_n52001_ = ~new_n51222_ & ~new_n51919_;
  assign new_n52002_ = ~new_n51232_ & new_n51866_;
  assign new_n52003_ = ~new_n51862_ & new_n52002_;
  assign new_n52004_ = ~new_n51863_ & ~new_n51866_;
  assign new_n52005_ = ~new_n52003_ & ~new_n52004_;
  assign new_n52006_ = new_n23895_ & ~new_n52005_;
  assign new_n52007_ = ~new_n51918_ & new_n52006_;
  assign new_n52008_ = ~new_n52001_ & ~new_n52007_;
  assign new_n52009_ = ~\b[48]  & ~new_n52008_;
  assign new_n52010_ = ~new_n51231_ & ~new_n51919_;
  assign new_n52011_ = ~new_n51241_ & new_n51861_;
  assign new_n52012_ = ~new_n51857_ & new_n52011_;
  assign new_n52013_ = ~new_n51858_ & ~new_n51861_;
  assign new_n52014_ = ~new_n52012_ & ~new_n52013_;
  assign new_n52015_ = new_n23895_ & ~new_n52014_;
  assign new_n52016_ = ~new_n51918_ & new_n52015_;
  assign new_n52017_ = ~new_n52010_ & ~new_n52016_;
  assign new_n52018_ = ~\b[47]  & ~new_n52017_;
  assign new_n52019_ = ~new_n51240_ & ~new_n51919_;
  assign new_n52020_ = ~new_n51250_ & new_n51856_;
  assign new_n52021_ = ~new_n51852_ & new_n52020_;
  assign new_n52022_ = ~new_n51853_ & ~new_n51856_;
  assign new_n52023_ = ~new_n52021_ & ~new_n52022_;
  assign new_n52024_ = new_n23895_ & ~new_n52023_;
  assign new_n52025_ = ~new_n51918_ & new_n52024_;
  assign new_n52026_ = ~new_n52019_ & ~new_n52025_;
  assign new_n52027_ = ~\b[46]  & ~new_n52026_;
  assign new_n52028_ = ~new_n51249_ & ~new_n51919_;
  assign new_n52029_ = ~new_n51259_ & new_n51851_;
  assign new_n52030_ = ~new_n51847_ & new_n52029_;
  assign new_n52031_ = ~new_n51848_ & ~new_n51851_;
  assign new_n52032_ = ~new_n52030_ & ~new_n52031_;
  assign new_n52033_ = new_n23895_ & ~new_n52032_;
  assign new_n52034_ = ~new_n51918_ & new_n52033_;
  assign new_n52035_ = ~new_n52028_ & ~new_n52034_;
  assign new_n52036_ = ~\b[45]  & ~new_n52035_;
  assign new_n52037_ = ~new_n51258_ & ~new_n51919_;
  assign new_n52038_ = ~new_n51268_ & new_n51846_;
  assign new_n52039_ = ~new_n51842_ & new_n52038_;
  assign new_n52040_ = ~new_n51843_ & ~new_n51846_;
  assign new_n52041_ = ~new_n52039_ & ~new_n52040_;
  assign new_n52042_ = new_n23895_ & ~new_n52041_;
  assign new_n52043_ = ~new_n51918_ & new_n52042_;
  assign new_n52044_ = ~new_n52037_ & ~new_n52043_;
  assign new_n52045_ = ~\b[44]  & ~new_n52044_;
  assign new_n52046_ = ~new_n51267_ & ~new_n51919_;
  assign new_n52047_ = ~new_n51277_ & new_n51841_;
  assign new_n52048_ = ~new_n51837_ & new_n52047_;
  assign new_n52049_ = ~new_n51838_ & ~new_n51841_;
  assign new_n52050_ = ~new_n52048_ & ~new_n52049_;
  assign new_n52051_ = new_n23895_ & ~new_n52050_;
  assign new_n52052_ = ~new_n51918_ & new_n52051_;
  assign new_n52053_ = ~new_n52046_ & ~new_n52052_;
  assign new_n52054_ = ~\b[43]  & ~new_n52053_;
  assign new_n52055_ = ~new_n51276_ & ~new_n51919_;
  assign new_n52056_ = ~new_n51286_ & new_n51836_;
  assign new_n52057_ = ~new_n51832_ & new_n52056_;
  assign new_n52058_ = ~new_n51833_ & ~new_n51836_;
  assign new_n52059_ = ~new_n52057_ & ~new_n52058_;
  assign new_n52060_ = new_n23895_ & ~new_n52059_;
  assign new_n52061_ = ~new_n51918_ & new_n52060_;
  assign new_n52062_ = ~new_n52055_ & ~new_n52061_;
  assign new_n52063_ = ~\b[42]  & ~new_n52062_;
  assign new_n52064_ = ~new_n51285_ & ~new_n51919_;
  assign new_n52065_ = ~new_n51295_ & new_n51831_;
  assign new_n52066_ = ~new_n51827_ & new_n52065_;
  assign new_n52067_ = ~new_n51828_ & ~new_n51831_;
  assign new_n52068_ = ~new_n52066_ & ~new_n52067_;
  assign new_n52069_ = new_n23895_ & ~new_n52068_;
  assign new_n52070_ = ~new_n51918_ & new_n52069_;
  assign new_n52071_ = ~new_n52064_ & ~new_n52070_;
  assign new_n52072_ = ~\b[41]  & ~new_n52071_;
  assign new_n52073_ = ~new_n51294_ & ~new_n51919_;
  assign new_n52074_ = ~new_n51304_ & new_n51826_;
  assign new_n52075_ = ~new_n51822_ & new_n52074_;
  assign new_n52076_ = ~new_n51823_ & ~new_n51826_;
  assign new_n52077_ = ~new_n52075_ & ~new_n52076_;
  assign new_n52078_ = new_n23895_ & ~new_n52077_;
  assign new_n52079_ = ~new_n51918_ & new_n52078_;
  assign new_n52080_ = ~new_n52073_ & ~new_n52079_;
  assign new_n52081_ = ~\b[40]  & ~new_n52080_;
  assign new_n52082_ = ~new_n51303_ & ~new_n51919_;
  assign new_n52083_ = ~new_n51313_ & new_n51821_;
  assign new_n52084_ = ~new_n51817_ & new_n52083_;
  assign new_n52085_ = ~new_n51818_ & ~new_n51821_;
  assign new_n52086_ = ~new_n52084_ & ~new_n52085_;
  assign new_n52087_ = new_n23895_ & ~new_n52086_;
  assign new_n52088_ = ~new_n51918_ & new_n52087_;
  assign new_n52089_ = ~new_n52082_ & ~new_n52088_;
  assign new_n52090_ = ~\b[39]  & ~new_n52089_;
  assign new_n52091_ = ~new_n51312_ & ~new_n51919_;
  assign new_n52092_ = ~new_n51322_ & new_n51816_;
  assign new_n52093_ = ~new_n51812_ & new_n52092_;
  assign new_n52094_ = ~new_n51813_ & ~new_n51816_;
  assign new_n52095_ = ~new_n52093_ & ~new_n52094_;
  assign new_n52096_ = new_n23895_ & ~new_n52095_;
  assign new_n52097_ = ~new_n51918_ & new_n52096_;
  assign new_n52098_ = ~new_n52091_ & ~new_n52097_;
  assign new_n52099_ = ~\b[38]  & ~new_n52098_;
  assign new_n52100_ = ~new_n51321_ & ~new_n51919_;
  assign new_n52101_ = ~new_n51331_ & new_n51811_;
  assign new_n52102_ = ~new_n51807_ & new_n52101_;
  assign new_n52103_ = ~new_n51808_ & ~new_n51811_;
  assign new_n52104_ = ~new_n52102_ & ~new_n52103_;
  assign new_n52105_ = new_n23895_ & ~new_n52104_;
  assign new_n52106_ = ~new_n51918_ & new_n52105_;
  assign new_n52107_ = ~new_n52100_ & ~new_n52106_;
  assign new_n52108_ = ~\b[37]  & ~new_n52107_;
  assign new_n52109_ = ~new_n51330_ & ~new_n51919_;
  assign new_n52110_ = ~new_n51340_ & new_n51806_;
  assign new_n52111_ = ~new_n51802_ & new_n52110_;
  assign new_n52112_ = ~new_n51803_ & ~new_n51806_;
  assign new_n52113_ = ~new_n52111_ & ~new_n52112_;
  assign new_n52114_ = new_n23895_ & ~new_n52113_;
  assign new_n52115_ = ~new_n51918_ & new_n52114_;
  assign new_n52116_ = ~new_n52109_ & ~new_n52115_;
  assign new_n52117_ = ~\b[36]  & ~new_n52116_;
  assign new_n52118_ = ~new_n51339_ & ~new_n51919_;
  assign new_n52119_ = ~new_n51349_ & new_n51801_;
  assign new_n52120_ = ~new_n51797_ & new_n52119_;
  assign new_n52121_ = ~new_n51798_ & ~new_n51801_;
  assign new_n52122_ = ~new_n52120_ & ~new_n52121_;
  assign new_n52123_ = new_n23895_ & ~new_n52122_;
  assign new_n52124_ = ~new_n51918_ & new_n52123_;
  assign new_n52125_ = ~new_n52118_ & ~new_n52124_;
  assign new_n52126_ = ~\b[35]  & ~new_n52125_;
  assign new_n52127_ = ~new_n51348_ & ~new_n51919_;
  assign new_n52128_ = ~new_n51358_ & new_n51796_;
  assign new_n52129_ = ~new_n51792_ & new_n52128_;
  assign new_n52130_ = ~new_n51793_ & ~new_n51796_;
  assign new_n52131_ = ~new_n52129_ & ~new_n52130_;
  assign new_n52132_ = new_n23895_ & ~new_n52131_;
  assign new_n52133_ = ~new_n51918_ & new_n52132_;
  assign new_n52134_ = ~new_n52127_ & ~new_n52133_;
  assign new_n52135_ = ~\b[34]  & ~new_n52134_;
  assign new_n52136_ = ~new_n51357_ & ~new_n51919_;
  assign new_n52137_ = ~new_n51367_ & new_n51791_;
  assign new_n52138_ = ~new_n51787_ & new_n52137_;
  assign new_n52139_ = ~new_n51788_ & ~new_n51791_;
  assign new_n52140_ = ~new_n52138_ & ~new_n52139_;
  assign new_n52141_ = new_n23895_ & ~new_n52140_;
  assign new_n52142_ = ~new_n51918_ & new_n52141_;
  assign new_n52143_ = ~new_n52136_ & ~new_n52142_;
  assign new_n52144_ = ~\b[33]  & ~new_n52143_;
  assign new_n52145_ = ~new_n51366_ & ~new_n51919_;
  assign new_n52146_ = ~new_n51376_ & new_n51786_;
  assign new_n52147_ = ~new_n51782_ & new_n52146_;
  assign new_n52148_ = ~new_n51783_ & ~new_n51786_;
  assign new_n52149_ = ~new_n52147_ & ~new_n52148_;
  assign new_n52150_ = new_n23895_ & ~new_n52149_;
  assign new_n52151_ = ~new_n51918_ & new_n52150_;
  assign new_n52152_ = ~new_n52145_ & ~new_n52151_;
  assign new_n52153_ = ~\b[32]  & ~new_n52152_;
  assign new_n52154_ = ~new_n51375_ & ~new_n51919_;
  assign new_n52155_ = ~new_n51385_ & new_n51781_;
  assign new_n52156_ = ~new_n51777_ & new_n52155_;
  assign new_n52157_ = ~new_n51778_ & ~new_n51781_;
  assign new_n52158_ = ~new_n52156_ & ~new_n52157_;
  assign new_n52159_ = new_n23895_ & ~new_n52158_;
  assign new_n52160_ = ~new_n51918_ & new_n52159_;
  assign new_n52161_ = ~new_n52154_ & ~new_n52160_;
  assign new_n52162_ = ~\b[31]  & ~new_n52161_;
  assign new_n52163_ = ~new_n51384_ & ~new_n51919_;
  assign new_n52164_ = ~new_n51394_ & new_n51776_;
  assign new_n52165_ = ~new_n51772_ & new_n52164_;
  assign new_n52166_ = ~new_n51773_ & ~new_n51776_;
  assign new_n52167_ = ~new_n52165_ & ~new_n52166_;
  assign new_n52168_ = new_n23895_ & ~new_n52167_;
  assign new_n52169_ = ~new_n51918_ & new_n52168_;
  assign new_n52170_ = ~new_n52163_ & ~new_n52169_;
  assign new_n52171_ = ~\b[30]  & ~new_n52170_;
  assign new_n52172_ = ~new_n51393_ & ~new_n51919_;
  assign new_n52173_ = ~new_n51403_ & new_n51771_;
  assign new_n52174_ = ~new_n51767_ & new_n52173_;
  assign new_n52175_ = ~new_n51768_ & ~new_n51771_;
  assign new_n52176_ = ~new_n52174_ & ~new_n52175_;
  assign new_n52177_ = new_n23895_ & ~new_n52176_;
  assign new_n52178_ = ~new_n51918_ & new_n52177_;
  assign new_n52179_ = ~new_n52172_ & ~new_n52178_;
  assign new_n52180_ = ~\b[29]  & ~new_n52179_;
  assign new_n52181_ = ~new_n51402_ & ~new_n51919_;
  assign new_n52182_ = ~new_n51412_ & new_n51766_;
  assign new_n52183_ = ~new_n51762_ & new_n52182_;
  assign new_n52184_ = ~new_n51763_ & ~new_n51766_;
  assign new_n52185_ = ~new_n52183_ & ~new_n52184_;
  assign new_n52186_ = new_n23895_ & ~new_n52185_;
  assign new_n52187_ = ~new_n51918_ & new_n52186_;
  assign new_n52188_ = ~new_n52181_ & ~new_n52187_;
  assign new_n52189_ = ~\b[28]  & ~new_n52188_;
  assign new_n52190_ = ~new_n51411_ & ~new_n51919_;
  assign new_n52191_ = ~new_n51421_ & new_n51761_;
  assign new_n52192_ = ~new_n51757_ & new_n52191_;
  assign new_n52193_ = ~new_n51758_ & ~new_n51761_;
  assign new_n52194_ = ~new_n52192_ & ~new_n52193_;
  assign new_n52195_ = new_n23895_ & ~new_n52194_;
  assign new_n52196_ = ~new_n51918_ & new_n52195_;
  assign new_n52197_ = ~new_n52190_ & ~new_n52196_;
  assign new_n52198_ = ~\b[27]  & ~new_n52197_;
  assign new_n52199_ = ~new_n51420_ & ~new_n51919_;
  assign new_n52200_ = ~new_n51430_ & new_n51756_;
  assign new_n52201_ = ~new_n51752_ & new_n52200_;
  assign new_n52202_ = ~new_n51753_ & ~new_n51756_;
  assign new_n52203_ = ~new_n52201_ & ~new_n52202_;
  assign new_n52204_ = new_n23895_ & ~new_n52203_;
  assign new_n52205_ = ~new_n51918_ & new_n52204_;
  assign new_n52206_ = ~new_n52199_ & ~new_n52205_;
  assign new_n52207_ = ~\b[26]  & ~new_n52206_;
  assign new_n52208_ = ~new_n51429_ & ~new_n51919_;
  assign new_n52209_ = ~new_n51439_ & new_n51751_;
  assign new_n52210_ = ~new_n51747_ & new_n52209_;
  assign new_n52211_ = ~new_n51748_ & ~new_n51751_;
  assign new_n52212_ = ~new_n52210_ & ~new_n52211_;
  assign new_n52213_ = new_n23895_ & ~new_n52212_;
  assign new_n52214_ = ~new_n51918_ & new_n52213_;
  assign new_n52215_ = ~new_n52208_ & ~new_n52214_;
  assign new_n52216_ = ~\b[25]  & ~new_n52215_;
  assign new_n52217_ = ~new_n51438_ & ~new_n51919_;
  assign new_n52218_ = ~new_n51448_ & new_n51746_;
  assign new_n52219_ = ~new_n51742_ & new_n52218_;
  assign new_n52220_ = ~new_n51743_ & ~new_n51746_;
  assign new_n52221_ = ~new_n52219_ & ~new_n52220_;
  assign new_n52222_ = new_n23895_ & ~new_n52221_;
  assign new_n52223_ = ~new_n51918_ & new_n52222_;
  assign new_n52224_ = ~new_n52217_ & ~new_n52223_;
  assign new_n52225_ = ~\b[24]  & ~new_n52224_;
  assign new_n52226_ = ~new_n51447_ & ~new_n51919_;
  assign new_n52227_ = ~new_n51457_ & new_n51741_;
  assign new_n52228_ = ~new_n51737_ & new_n52227_;
  assign new_n52229_ = ~new_n51738_ & ~new_n51741_;
  assign new_n52230_ = ~new_n52228_ & ~new_n52229_;
  assign new_n52231_ = new_n23895_ & ~new_n52230_;
  assign new_n52232_ = ~new_n51918_ & new_n52231_;
  assign new_n52233_ = ~new_n52226_ & ~new_n52232_;
  assign new_n52234_ = ~\b[23]  & ~new_n52233_;
  assign new_n52235_ = ~new_n51456_ & ~new_n51919_;
  assign new_n52236_ = ~new_n51466_ & new_n51736_;
  assign new_n52237_ = ~new_n51732_ & new_n52236_;
  assign new_n52238_ = ~new_n51733_ & ~new_n51736_;
  assign new_n52239_ = ~new_n52237_ & ~new_n52238_;
  assign new_n52240_ = new_n23895_ & ~new_n52239_;
  assign new_n52241_ = ~new_n51918_ & new_n52240_;
  assign new_n52242_ = ~new_n52235_ & ~new_n52241_;
  assign new_n52243_ = ~\b[22]  & ~new_n52242_;
  assign new_n52244_ = ~new_n51465_ & ~new_n51919_;
  assign new_n52245_ = ~new_n51475_ & new_n51731_;
  assign new_n52246_ = ~new_n51727_ & new_n52245_;
  assign new_n52247_ = ~new_n51728_ & ~new_n51731_;
  assign new_n52248_ = ~new_n52246_ & ~new_n52247_;
  assign new_n52249_ = new_n23895_ & ~new_n52248_;
  assign new_n52250_ = ~new_n51918_ & new_n52249_;
  assign new_n52251_ = ~new_n52244_ & ~new_n52250_;
  assign new_n52252_ = ~\b[21]  & ~new_n52251_;
  assign new_n52253_ = ~new_n51474_ & ~new_n51919_;
  assign new_n52254_ = ~new_n51484_ & new_n51726_;
  assign new_n52255_ = ~new_n51722_ & new_n52254_;
  assign new_n52256_ = ~new_n51723_ & ~new_n51726_;
  assign new_n52257_ = ~new_n52255_ & ~new_n52256_;
  assign new_n52258_ = new_n23895_ & ~new_n52257_;
  assign new_n52259_ = ~new_n51918_ & new_n52258_;
  assign new_n52260_ = ~new_n52253_ & ~new_n52259_;
  assign new_n52261_ = ~\b[20]  & ~new_n52260_;
  assign new_n52262_ = ~new_n51483_ & ~new_n51919_;
  assign new_n52263_ = ~new_n51493_ & new_n51721_;
  assign new_n52264_ = ~new_n51717_ & new_n52263_;
  assign new_n52265_ = ~new_n51718_ & ~new_n51721_;
  assign new_n52266_ = ~new_n52264_ & ~new_n52265_;
  assign new_n52267_ = new_n23895_ & ~new_n52266_;
  assign new_n52268_ = ~new_n51918_ & new_n52267_;
  assign new_n52269_ = ~new_n52262_ & ~new_n52268_;
  assign new_n52270_ = ~\b[19]  & ~new_n52269_;
  assign new_n52271_ = ~new_n51492_ & ~new_n51919_;
  assign new_n52272_ = ~new_n51502_ & new_n51716_;
  assign new_n52273_ = ~new_n51712_ & new_n52272_;
  assign new_n52274_ = ~new_n51713_ & ~new_n51716_;
  assign new_n52275_ = ~new_n52273_ & ~new_n52274_;
  assign new_n52276_ = new_n23895_ & ~new_n52275_;
  assign new_n52277_ = ~new_n51918_ & new_n52276_;
  assign new_n52278_ = ~new_n52271_ & ~new_n52277_;
  assign new_n52279_ = ~\b[18]  & ~new_n52278_;
  assign new_n52280_ = ~new_n51501_ & ~new_n51919_;
  assign new_n52281_ = ~new_n51511_ & new_n51711_;
  assign new_n52282_ = ~new_n51707_ & new_n52281_;
  assign new_n52283_ = ~new_n51708_ & ~new_n51711_;
  assign new_n52284_ = ~new_n52282_ & ~new_n52283_;
  assign new_n52285_ = new_n23895_ & ~new_n52284_;
  assign new_n52286_ = ~new_n51918_ & new_n52285_;
  assign new_n52287_ = ~new_n52280_ & ~new_n52286_;
  assign new_n52288_ = ~\b[17]  & ~new_n52287_;
  assign new_n52289_ = ~new_n51510_ & ~new_n51919_;
  assign new_n52290_ = ~new_n51520_ & new_n51706_;
  assign new_n52291_ = ~new_n51702_ & new_n52290_;
  assign new_n52292_ = ~new_n51703_ & ~new_n51706_;
  assign new_n52293_ = ~new_n52291_ & ~new_n52292_;
  assign new_n52294_ = new_n23895_ & ~new_n52293_;
  assign new_n52295_ = ~new_n51918_ & new_n52294_;
  assign new_n52296_ = ~new_n52289_ & ~new_n52295_;
  assign new_n52297_ = ~\b[16]  & ~new_n52296_;
  assign new_n52298_ = ~new_n51519_ & ~new_n51919_;
  assign new_n52299_ = ~new_n51529_ & new_n51701_;
  assign new_n52300_ = ~new_n51697_ & new_n52299_;
  assign new_n52301_ = ~new_n51698_ & ~new_n51701_;
  assign new_n52302_ = ~new_n52300_ & ~new_n52301_;
  assign new_n52303_ = new_n23895_ & ~new_n52302_;
  assign new_n52304_ = ~new_n51918_ & new_n52303_;
  assign new_n52305_ = ~new_n52298_ & ~new_n52304_;
  assign new_n52306_ = ~\b[15]  & ~new_n52305_;
  assign new_n52307_ = ~new_n51528_ & ~new_n51919_;
  assign new_n52308_ = ~new_n51538_ & new_n51696_;
  assign new_n52309_ = ~new_n51692_ & new_n52308_;
  assign new_n52310_ = ~new_n51693_ & ~new_n51696_;
  assign new_n52311_ = ~new_n52309_ & ~new_n52310_;
  assign new_n52312_ = new_n23895_ & ~new_n52311_;
  assign new_n52313_ = ~new_n51918_ & new_n52312_;
  assign new_n52314_ = ~new_n52307_ & ~new_n52313_;
  assign new_n52315_ = ~\b[14]  & ~new_n52314_;
  assign new_n52316_ = ~new_n51537_ & ~new_n51919_;
  assign new_n52317_ = ~new_n51547_ & new_n51691_;
  assign new_n52318_ = ~new_n51687_ & new_n52317_;
  assign new_n52319_ = ~new_n51688_ & ~new_n51691_;
  assign new_n52320_ = ~new_n52318_ & ~new_n52319_;
  assign new_n52321_ = new_n23895_ & ~new_n52320_;
  assign new_n52322_ = ~new_n51918_ & new_n52321_;
  assign new_n52323_ = ~new_n52316_ & ~new_n52322_;
  assign new_n52324_ = ~\b[13]  & ~new_n52323_;
  assign new_n52325_ = ~new_n51546_ & ~new_n51919_;
  assign new_n52326_ = ~new_n51556_ & new_n51686_;
  assign new_n52327_ = ~new_n51682_ & new_n52326_;
  assign new_n52328_ = ~new_n51683_ & ~new_n51686_;
  assign new_n52329_ = ~new_n52327_ & ~new_n52328_;
  assign new_n52330_ = new_n23895_ & ~new_n52329_;
  assign new_n52331_ = ~new_n51918_ & new_n52330_;
  assign new_n52332_ = ~new_n52325_ & ~new_n52331_;
  assign new_n52333_ = ~\b[12]  & ~new_n52332_;
  assign new_n52334_ = ~new_n51555_ & ~new_n51919_;
  assign new_n52335_ = ~new_n51565_ & new_n51681_;
  assign new_n52336_ = ~new_n51677_ & new_n52335_;
  assign new_n52337_ = ~new_n51678_ & ~new_n51681_;
  assign new_n52338_ = ~new_n52336_ & ~new_n52337_;
  assign new_n52339_ = new_n23895_ & ~new_n52338_;
  assign new_n52340_ = ~new_n51918_ & new_n52339_;
  assign new_n52341_ = ~new_n52334_ & ~new_n52340_;
  assign new_n52342_ = ~\b[11]  & ~new_n52341_;
  assign new_n52343_ = ~new_n51564_ & ~new_n51919_;
  assign new_n52344_ = ~new_n51574_ & new_n51676_;
  assign new_n52345_ = ~new_n51672_ & new_n52344_;
  assign new_n52346_ = ~new_n51673_ & ~new_n51676_;
  assign new_n52347_ = ~new_n52345_ & ~new_n52346_;
  assign new_n52348_ = new_n23895_ & ~new_n52347_;
  assign new_n52349_ = ~new_n51918_ & new_n52348_;
  assign new_n52350_ = ~new_n52343_ & ~new_n52349_;
  assign new_n52351_ = ~\b[10]  & ~new_n52350_;
  assign new_n52352_ = ~new_n51573_ & ~new_n51919_;
  assign new_n52353_ = ~new_n51583_ & new_n51671_;
  assign new_n52354_ = ~new_n51667_ & new_n52353_;
  assign new_n52355_ = ~new_n51668_ & ~new_n51671_;
  assign new_n52356_ = ~new_n52354_ & ~new_n52355_;
  assign new_n52357_ = new_n23895_ & ~new_n52356_;
  assign new_n52358_ = ~new_n51918_ & new_n52357_;
  assign new_n52359_ = ~new_n52352_ & ~new_n52358_;
  assign new_n52360_ = ~\b[9]  & ~new_n52359_;
  assign new_n52361_ = ~new_n51582_ & ~new_n51919_;
  assign new_n52362_ = ~new_n51592_ & new_n51666_;
  assign new_n52363_ = ~new_n51662_ & new_n52362_;
  assign new_n52364_ = ~new_n51663_ & ~new_n51666_;
  assign new_n52365_ = ~new_n52363_ & ~new_n52364_;
  assign new_n52366_ = new_n23895_ & ~new_n52365_;
  assign new_n52367_ = ~new_n51918_ & new_n52366_;
  assign new_n52368_ = ~new_n52361_ & ~new_n52367_;
  assign new_n52369_ = ~\b[8]  & ~new_n52368_;
  assign new_n52370_ = ~new_n51591_ & ~new_n51919_;
  assign new_n52371_ = ~new_n51601_ & new_n51661_;
  assign new_n52372_ = ~new_n51657_ & new_n52371_;
  assign new_n52373_ = ~new_n51658_ & ~new_n51661_;
  assign new_n52374_ = ~new_n52372_ & ~new_n52373_;
  assign new_n52375_ = new_n23895_ & ~new_n52374_;
  assign new_n52376_ = ~new_n51918_ & new_n52375_;
  assign new_n52377_ = ~new_n52370_ & ~new_n52376_;
  assign new_n52378_ = ~\b[7]  & ~new_n52377_;
  assign new_n52379_ = ~new_n51600_ & ~new_n51919_;
  assign new_n52380_ = ~new_n51610_ & new_n51656_;
  assign new_n52381_ = ~new_n51652_ & new_n52380_;
  assign new_n52382_ = ~new_n51653_ & ~new_n51656_;
  assign new_n52383_ = ~new_n52381_ & ~new_n52382_;
  assign new_n52384_ = new_n23895_ & ~new_n52383_;
  assign new_n52385_ = ~new_n51918_ & new_n52384_;
  assign new_n52386_ = ~new_n52379_ & ~new_n52385_;
  assign new_n52387_ = ~\b[6]  & ~new_n52386_;
  assign new_n52388_ = ~new_n51609_ & ~new_n51919_;
  assign new_n52389_ = ~new_n51619_ & new_n51651_;
  assign new_n52390_ = ~new_n51647_ & new_n52389_;
  assign new_n52391_ = ~new_n51648_ & ~new_n51651_;
  assign new_n52392_ = ~new_n52390_ & ~new_n52391_;
  assign new_n52393_ = new_n23895_ & ~new_n52392_;
  assign new_n52394_ = ~new_n51918_ & new_n52393_;
  assign new_n52395_ = ~new_n52388_ & ~new_n52394_;
  assign new_n52396_ = ~\b[5]  & ~new_n52395_;
  assign new_n52397_ = ~new_n51618_ & ~new_n51919_;
  assign new_n52398_ = ~new_n51627_ & new_n51646_;
  assign new_n52399_ = ~new_n51642_ & new_n52398_;
  assign new_n52400_ = ~new_n51643_ & ~new_n51646_;
  assign new_n52401_ = ~new_n52399_ & ~new_n52400_;
  assign new_n52402_ = new_n23895_ & ~new_n52401_;
  assign new_n52403_ = ~new_n51918_ & new_n52402_;
  assign new_n52404_ = ~new_n52397_ & ~new_n52403_;
  assign new_n52405_ = ~\b[4]  & ~new_n52404_;
  assign new_n52406_ = ~new_n51626_ & ~new_n51919_;
  assign new_n52407_ = ~new_n51637_ & new_n51641_;
  assign new_n52408_ = ~new_n51636_ & new_n52407_;
  assign new_n52409_ = ~new_n51638_ & ~new_n51641_;
  assign new_n52410_ = ~new_n52408_ & ~new_n52409_;
  assign new_n52411_ = new_n23895_ & ~new_n52410_;
  assign new_n52412_ = ~new_n51918_ & new_n52411_;
  assign new_n52413_ = ~new_n52406_ & ~new_n52412_;
  assign new_n52414_ = ~\b[3]  & ~new_n52413_;
  assign new_n52415_ = ~new_n51631_ & ~new_n51919_;
  assign new_n52416_ = new_n23611_ & ~new_n51634_;
  assign new_n52417_ = ~new_n51632_ & new_n52416_;
  assign new_n52418_ = new_n23895_ & ~new_n52417_;
  assign new_n52419_ = ~new_n51636_ & new_n52418_;
  assign new_n52420_ = ~new_n51918_ & new_n52419_;
  assign new_n52421_ = ~new_n52415_ & ~new_n52420_;
  assign new_n52422_ = ~\b[2]  & ~new_n52421_;
  assign new_n52423_ = new_n24402_ & ~new_n51918_;
  assign new_n52424_ = \a[6]  & ~new_n52423_;
  assign new_n52425_ = new_n24406_ & ~new_n51918_;
  assign new_n52426_ = ~new_n52424_ & ~new_n52425_;
  assign new_n52427_ = \b[1]  & ~new_n52426_;
  assign new_n52428_ = ~\b[1]  & ~new_n52425_;
  assign new_n52429_ = ~new_n52424_ & new_n52428_;
  assign new_n52430_ = ~new_n52427_ & ~new_n52429_;
  assign new_n52431_ = ~new_n24413_ & ~new_n52430_;
  assign new_n52432_ = ~\b[1]  & ~new_n52426_;
  assign new_n52433_ = ~new_n52431_ & ~new_n52432_;
  assign new_n52434_ = \b[2]  & ~new_n52420_;
  assign new_n52435_ = ~new_n52415_ & new_n52434_;
  assign new_n52436_ = ~new_n52422_ & ~new_n52435_;
  assign new_n52437_ = ~new_n52433_ & new_n52436_;
  assign new_n52438_ = ~new_n52422_ & ~new_n52437_;
  assign new_n52439_ = \b[3]  & ~new_n52412_;
  assign new_n52440_ = ~new_n52406_ & new_n52439_;
  assign new_n52441_ = ~new_n52414_ & ~new_n52440_;
  assign new_n52442_ = ~new_n52438_ & new_n52441_;
  assign new_n52443_ = ~new_n52414_ & ~new_n52442_;
  assign new_n52444_ = \b[4]  & ~new_n52403_;
  assign new_n52445_ = ~new_n52397_ & new_n52444_;
  assign new_n52446_ = ~new_n52405_ & ~new_n52445_;
  assign new_n52447_ = ~new_n52443_ & new_n52446_;
  assign new_n52448_ = ~new_n52405_ & ~new_n52447_;
  assign new_n52449_ = \b[5]  & ~new_n52394_;
  assign new_n52450_ = ~new_n52388_ & new_n52449_;
  assign new_n52451_ = ~new_n52396_ & ~new_n52450_;
  assign new_n52452_ = ~new_n52448_ & new_n52451_;
  assign new_n52453_ = ~new_n52396_ & ~new_n52452_;
  assign new_n52454_ = \b[6]  & ~new_n52385_;
  assign new_n52455_ = ~new_n52379_ & new_n52454_;
  assign new_n52456_ = ~new_n52387_ & ~new_n52455_;
  assign new_n52457_ = ~new_n52453_ & new_n52456_;
  assign new_n52458_ = ~new_n52387_ & ~new_n52457_;
  assign new_n52459_ = \b[7]  & ~new_n52376_;
  assign new_n52460_ = ~new_n52370_ & new_n52459_;
  assign new_n52461_ = ~new_n52378_ & ~new_n52460_;
  assign new_n52462_ = ~new_n52458_ & new_n52461_;
  assign new_n52463_ = ~new_n52378_ & ~new_n52462_;
  assign new_n52464_ = \b[8]  & ~new_n52367_;
  assign new_n52465_ = ~new_n52361_ & new_n52464_;
  assign new_n52466_ = ~new_n52369_ & ~new_n52465_;
  assign new_n52467_ = ~new_n52463_ & new_n52466_;
  assign new_n52468_ = ~new_n52369_ & ~new_n52467_;
  assign new_n52469_ = \b[9]  & ~new_n52358_;
  assign new_n52470_ = ~new_n52352_ & new_n52469_;
  assign new_n52471_ = ~new_n52360_ & ~new_n52470_;
  assign new_n52472_ = ~new_n52468_ & new_n52471_;
  assign new_n52473_ = ~new_n52360_ & ~new_n52472_;
  assign new_n52474_ = \b[10]  & ~new_n52349_;
  assign new_n52475_ = ~new_n52343_ & new_n52474_;
  assign new_n52476_ = ~new_n52351_ & ~new_n52475_;
  assign new_n52477_ = ~new_n52473_ & new_n52476_;
  assign new_n52478_ = ~new_n52351_ & ~new_n52477_;
  assign new_n52479_ = \b[11]  & ~new_n52340_;
  assign new_n52480_ = ~new_n52334_ & new_n52479_;
  assign new_n52481_ = ~new_n52342_ & ~new_n52480_;
  assign new_n52482_ = ~new_n52478_ & new_n52481_;
  assign new_n52483_ = ~new_n52342_ & ~new_n52482_;
  assign new_n52484_ = \b[12]  & ~new_n52331_;
  assign new_n52485_ = ~new_n52325_ & new_n52484_;
  assign new_n52486_ = ~new_n52333_ & ~new_n52485_;
  assign new_n52487_ = ~new_n52483_ & new_n52486_;
  assign new_n52488_ = ~new_n52333_ & ~new_n52487_;
  assign new_n52489_ = \b[13]  & ~new_n52322_;
  assign new_n52490_ = ~new_n52316_ & new_n52489_;
  assign new_n52491_ = ~new_n52324_ & ~new_n52490_;
  assign new_n52492_ = ~new_n52488_ & new_n52491_;
  assign new_n52493_ = ~new_n52324_ & ~new_n52492_;
  assign new_n52494_ = \b[14]  & ~new_n52313_;
  assign new_n52495_ = ~new_n52307_ & new_n52494_;
  assign new_n52496_ = ~new_n52315_ & ~new_n52495_;
  assign new_n52497_ = ~new_n52493_ & new_n52496_;
  assign new_n52498_ = ~new_n52315_ & ~new_n52497_;
  assign new_n52499_ = \b[15]  & ~new_n52304_;
  assign new_n52500_ = ~new_n52298_ & new_n52499_;
  assign new_n52501_ = ~new_n52306_ & ~new_n52500_;
  assign new_n52502_ = ~new_n52498_ & new_n52501_;
  assign new_n52503_ = ~new_n52306_ & ~new_n52502_;
  assign new_n52504_ = \b[16]  & ~new_n52295_;
  assign new_n52505_ = ~new_n52289_ & new_n52504_;
  assign new_n52506_ = ~new_n52297_ & ~new_n52505_;
  assign new_n52507_ = ~new_n52503_ & new_n52506_;
  assign new_n52508_ = ~new_n52297_ & ~new_n52507_;
  assign new_n52509_ = \b[17]  & ~new_n52286_;
  assign new_n52510_ = ~new_n52280_ & new_n52509_;
  assign new_n52511_ = ~new_n52288_ & ~new_n52510_;
  assign new_n52512_ = ~new_n52508_ & new_n52511_;
  assign new_n52513_ = ~new_n52288_ & ~new_n52512_;
  assign new_n52514_ = \b[18]  & ~new_n52277_;
  assign new_n52515_ = ~new_n52271_ & new_n52514_;
  assign new_n52516_ = ~new_n52279_ & ~new_n52515_;
  assign new_n52517_ = ~new_n52513_ & new_n52516_;
  assign new_n52518_ = ~new_n52279_ & ~new_n52517_;
  assign new_n52519_ = \b[19]  & ~new_n52268_;
  assign new_n52520_ = ~new_n52262_ & new_n52519_;
  assign new_n52521_ = ~new_n52270_ & ~new_n52520_;
  assign new_n52522_ = ~new_n52518_ & new_n52521_;
  assign new_n52523_ = ~new_n52270_ & ~new_n52522_;
  assign new_n52524_ = \b[20]  & ~new_n52259_;
  assign new_n52525_ = ~new_n52253_ & new_n52524_;
  assign new_n52526_ = ~new_n52261_ & ~new_n52525_;
  assign new_n52527_ = ~new_n52523_ & new_n52526_;
  assign new_n52528_ = ~new_n52261_ & ~new_n52527_;
  assign new_n52529_ = \b[21]  & ~new_n52250_;
  assign new_n52530_ = ~new_n52244_ & new_n52529_;
  assign new_n52531_ = ~new_n52252_ & ~new_n52530_;
  assign new_n52532_ = ~new_n52528_ & new_n52531_;
  assign new_n52533_ = ~new_n52252_ & ~new_n52532_;
  assign new_n52534_ = \b[22]  & ~new_n52241_;
  assign new_n52535_ = ~new_n52235_ & new_n52534_;
  assign new_n52536_ = ~new_n52243_ & ~new_n52535_;
  assign new_n52537_ = ~new_n52533_ & new_n52536_;
  assign new_n52538_ = ~new_n52243_ & ~new_n52537_;
  assign new_n52539_ = \b[23]  & ~new_n52232_;
  assign new_n52540_ = ~new_n52226_ & new_n52539_;
  assign new_n52541_ = ~new_n52234_ & ~new_n52540_;
  assign new_n52542_ = ~new_n52538_ & new_n52541_;
  assign new_n52543_ = ~new_n52234_ & ~new_n52542_;
  assign new_n52544_ = \b[24]  & ~new_n52223_;
  assign new_n52545_ = ~new_n52217_ & new_n52544_;
  assign new_n52546_ = ~new_n52225_ & ~new_n52545_;
  assign new_n52547_ = ~new_n52543_ & new_n52546_;
  assign new_n52548_ = ~new_n52225_ & ~new_n52547_;
  assign new_n52549_ = \b[25]  & ~new_n52214_;
  assign new_n52550_ = ~new_n52208_ & new_n52549_;
  assign new_n52551_ = ~new_n52216_ & ~new_n52550_;
  assign new_n52552_ = ~new_n52548_ & new_n52551_;
  assign new_n52553_ = ~new_n52216_ & ~new_n52552_;
  assign new_n52554_ = \b[26]  & ~new_n52205_;
  assign new_n52555_ = ~new_n52199_ & new_n52554_;
  assign new_n52556_ = ~new_n52207_ & ~new_n52555_;
  assign new_n52557_ = ~new_n52553_ & new_n52556_;
  assign new_n52558_ = ~new_n52207_ & ~new_n52557_;
  assign new_n52559_ = \b[27]  & ~new_n52196_;
  assign new_n52560_ = ~new_n52190_ & new_n52559_;
  assign new_n52561_ = ~new_n52198_ & ~new_n52560_;
  assign new_n52562_ = ~new_n52558_ & new_n52561_;
  assign new_n52563_ = ~new_n52198_ & ~new_n52562_;
  assign new_n52564_ = \b[28]  & ~new_n52187_;
  assign new_n52565_ = ~new_n52181_ & new_n52564_;
  assign new_n52566_ = ~new_n52189_ & ~new_n52565_;
  assign new_n52567_ = ~new_n52563_ & new_n52566_;
  assign new_n52568_ = ~new_n52189_ & ~new_n52567_;
  assign new_n52569_ = \b[29]  & ~new_n52178_;
  assign new_n52570_ = ~new_n52172_ & new_n52569_;
  assign new_n52571_ = ~new_n52180_ & ~new_n52570_;
  assign new_n52572_ = ~new_n52568_ & new_n52571_;
  assign new_n52573_ = ~new_n52180_ & ~new_n52572_;
  assign new_n52574_ = \b[30]  & ~new_n52169_;
  assign new_n52575_ = ~new_n52163_ & new_n52574_;
  assign new_n52576_ = ~new_n52171_ & ~new_n52575_;
  assign new_n52577_ = ~new_n52573_ & new_n52576_;
  assign new_n52578_ = ~new_n52171_ & ~new_n52577_;
  assign new_n52579_ = \b[31]  & ~new_n52160_;
  assign new_n52580_ = ~new_n52154_ & new_n52579_;
  assign new_n52581_ = ~new_n52162_ & ~new_n52580_;
  assign new_n52582_ = ~new_n52578_ & new_n52581_;
  assign new_n52583_ = ~new_n52162_ & ~new_n52582_;
  assign new_n52584_ = \b[32]  & ~new_n52151_;
  assign new_n52585_ = ~new_n52145_ & new_n52584_;
  assign new_n52586_ = ~new_n52153_ & ~new_n52585_;
  assign new_n52587_ = ~new_n52583_ & new_n52586_;
  assign new_n52588_ = ~new_n52153_ & ~new_n52587_;
  assign new_n52589_ = \b[33]  & ~new_n52142_;
  assign new_n52590_ = ~new_n52136_ & new_n52589_;
  assign new_n52591_ = ~new_n52144_ & ~new_n52590_;
  assign new_n52592_ = ~new_n52588_ & new_n52591_;
  assign new_n52593_ = ~new_n52144_ & ~new_n52592_;
  assign new_n52594_ = \b[34]  & ~new_n52133_;
  assign new_n52595_ = ~new_n52127_ & new_n52594_;
  assign new_n52596_ = ~new_n52135_ & ~new_n52595_;
  assign new_n52597_ = ~new_n52593_ & new_n52596_;
  assign new_n52598_ = ~new_n52135_ & ~new_n52597_;
  assign new_n52599_ = \b[35]  & ~new_n52124_;
  assign new_n52600_ = ~new_n52118_ & new_n52599_;
  assign new_n52601_ = ~new_n52126_ & ~new_n52600_;
  assign new_n52602_ = ~new_n52598_ & new_n52601_;
  assign new_n52603_ = ~new_n52126_ & ~new_n52602_;
  assign new_n52604_ = \b[36]  & ~new_n52115_;
  assign new_n52605_ = ~new_n52109_ & new_n52604_;
  assign new_n52606_ = ~new_n52117_ & ~new_n52605_;
  assign new_n52607_ = ~new_n52603_ & new_n52606_;
  assign new_n52608_ = ~new_n52117_ & ~new_n52607_;
  assign new_n52609_ = \b[37]  & ~new_n52106_;
  assign new_n52610_ = ~new_n52100_ & new_n52609_;
  assign new_n52611_ = ~new_n52108_ & ~new_n52610_;
  assign new_n52612_ = ~new_n52608_ & new_n52611_;
  assign new_n52613_ = ~new_n52108_ & ~new_n52612_;
  assign new_n52614_ = \b[38]  & ~new_n52097_;
  assign new_n52615_ = ~new_n52091_ & new_n52614_;
  assign new_n52616_ = ~new_n52099_ & ~new_n52615_;
  assign new_n52617_ = ~new_n52613_ & new_n52616_;
  assign new_n52618_ = ~new_n52099_ & ~new_n52617_;
  assign new_n52619_ = \b[39]  & ~new_n52088_;
  assign new_n52620_ = ~new_n52082_ & new_n52619_;
  assign new_n52621_ = ~new_n52090_ & ~new_n52620_;
  assign new_n52622_ = ~new_n52618_ & new_n52621_;
  assign new_n52623_ = ~new_n52090_ & ~new_n52622_;
  assign new_n52624_ = \b[40]  & ~new_n52079_;
  assign new_n52625_ = ~new_n52073_ & new_n52624_;
  assign new_n52626_ = ~new_n52081_ & ~new_n52625_;
  assign new_n52627_ = ~new_n52623_ & new_n52626_;
  assign new_n52628_ = ~new_n52081_ & ~new_n52627_;
  assign new_n52629_ = \b[41]  & ~new_n52070_;
  assign new_n52630_ = ~new_n52064_ & new_n52629_;
  assign new_n52631_ = ~new_n52072_ & ~new_n52630_;
  assign new_n52632_ = ~new_n52628_ & new_n52631_;
  assign new_n52633_ = ~new_n52072_ & ~new_n52632_;
  assign new_n52634_ = \b[42]  & ~new_n52061_;
  assign new_n52635_ = ~new_n52055_ & new_n52634_;
  assign new_n52636_ = ~new_n52063_ & ~new_n52635_;
  assign new_n52637_ = ~new_n52633_ & new_n52636_;
  assign new_n52638_ = ~new_n52063_ & ~new_n52637_;
  assign new_n52639_ = \b[43]  & ~new_n52052_;
  assign new_n52640_ = ~new_n52046_ & new_n52639_;
  assign new_n52641_ = ~new_n52054_ & ~new_n52640_;
  assign new_n52642_ = ~new_n52638_ & new_n52641_;
  assign new_n52643_ = ~new_n52054_ & ~new_n52642_;
  assign new_n52644_ = \b[44]  & ~new_n52043_;
  assign new_n52645_ = ~new_n52037_ & new_n52644_;
  assign new_n52646_ = ~new_n52045_ & ~new_n52645_;
  assign new_n52647_ = ~new_n52643_ & new_n52646_;
  assign new_n52648_ = ~new_n52045_ & ~new_n52647_;
  assign new_n52649_ = \b[45]  & ~new_n52034_;
  assign new_n52650_ = ~new_n52028_ & new_n52649_;
  assign new_n52651_ = ~new_n52036_ & ~new_n52650_;
  assign new_n52652_ = ~new_n52648_ & new_n52651_;
  assign new_n52653_ = ~new_n52036_ & ~new_n52652_;
  assign new_n52654_ = \b[46]  & ~new_n52025_;
  assign new_n52655_ = ~new_n52019_ & new_n52654_;
  assign new_n52656_ = ~new_n52027_ & ~new_n52655_;
  assign new_n52657_ = ~new_n52653_ & new_n52656_;
  assign new_n52658_ = ~new_n52027_ & ~new_n52657_;
  assign new_n52659_ = \b[47]  & ~new_n52016_;
  assign new_n52660_ = ~new_n52010_ & new_n52659_;
  assign new_n52661_ = ~new_n52018_ & ~new_n52660_;
  assign new_n52662_ = ~new_n52658_ & new_n52661_;
  assign new_n52663_ = ~new_n52018_ & ~new_n52662_;
  assign new_n52664_ = \b[48]  & ~new_n52007_;
  assign new_n52665_ = ~new_n52001_ & new_n52664_;
  assign new_n52666_ = ~new_n52009_ & ~new_n52665_;
  assign new_n52667_ = ~new_n52663_ & new_n52666_;
  assign new_n52668_ = ~new_n52009_ & ~new_n52667_;
  assign new_n52669_ = \b[49]  & ~new_n51998_;
  assign new_n52670_ = ~new_n51992_ & new_n52669_;
  assign new_n52671_ = ~new_n52000_ & ~new_n52670_;
  assign new_n52672_ = ~new_n52668_ & new_n52671_;
  assign new_n52673_ = ~new_n52000_ & ~new_n52672_;
  assign new_n52674_ = \b[50]  & ~new_n51989_;
  assign new_n52675_ = ~new_n51983_ & new_n52674_;
  assign new_n52676_ = ~new_n51991_ & ~new_n52675_;
  assign new_n52677_ = ~new_n52673_ & new_n52676_;
  assign new_n52678_ = ~new_n51991_ & ~new_n52677_;
  assign new_n52679_ = \b[51]  & ~new_n51980_;
  assign new_n52680_ = ~new_n51974_ & new_n52679_;
  assign new_n52681_ = ~new_n51982_ & ~new_n52680_;
  assign new_n52682_ = ~new_n52678_ & new_n52681_;
  assign new_n52683_ = ~new_n51982_ & ~new_n52682_;
  assign new_n52684_ = \b[52]  & ~new_n51971_;
  assign new_n52685_ = ~new_n51965_ & new_n52684_;
  assign new_n52686_ = ~new_n51973_ & ~new_n52685_;
  assign new_n52687_ = ~new_n52683_ & new_n52686_;
  assign new_n52688_ = ~new_n51973_ & ~new_n52687_;
  assign new_n52689_ = \b[53]  & ~new_n51962_;
  assign new_n52690_ = ~new_n51956_ & new_n52689_;
  assign new_n52691_ = ~new_n51964_ & ~new_n52690_;
  assign new_n52692_ = ~new_n52688_ & new_n52691_;
  assign new_n52693_ = ~new_n51964_ & ~new_n52692_;
  assign new_n52694_ = \b[54]  & ~new_n51953_;
  assign new_n52695_ = ~new_n51947_ & new_n52694_;
  assign new_n52696_ = ~new_n51955_ & ~new_n52695_;
  assign new_n52697_ = ~new_n52693_ & new_n52696_;
  assign new_n52698_ = ~new_n51955_ & ~new_n52697_;
  assign new_n52699_ = \b[55]  & ~new_n51944_;
  assign new_n52700_ = ~new_n51938_ & new_n52699_;
  assign new_n52701_ = ~new_n51946_ & ~new_n52700_;
  assign new_n52702_ = ~new_n52698_ & new_n52701_;
  assign new_n52703_ = ~new_n51946_ & ~new_n52702_;
  assign new_n52704_ = \b[56]  & ~new_n51935_;
  assign new_n52705_ = ~new_n51929_ & new_n52704_;
  assign new_n52706_ = ~new_n51937_ & ~new_n52705_;
  assign new_n52707_ = ~new_n52703_ & new_n52706_;
  assign new_n52708_ = ~new_n51937_ & ~new_n52707_;
  assign new_n52709_ = \b[57]  & ~new_n51926_;
  assign new_n52710_ = ~new_n51920_ & new_n52709_;
  assign new_n52711_ = ~new_n51928_ & ~new_n52710_;
  assign new_n52712_ = ~new_n52708_ & new_n52711_;
  assign new_n52713_ = ~new_n51928_ & ~new_n52712_;
  assign new_n52714_ = ~new_n51140_ & ~new_n51919_;
  assign new_n52715_ = ~new_n51142_ & new_n51916_;
  assign new_n52716_ = ~new_n51912_ & new_n52715_;
  assign new_n52717_ = ~new_n51913_ & ~new_n51916_;
  assign new_n52718_ = ~new_n52716_ & ~new_n52717_;
  assign new_n52719_ = new_n51919_ & ~new_n52718_;
  assign new_n52720_ = ~new_n52714_ & ~new_n52719_;
  assign new_n52721_ = ~\b[58]  & ~new_n52720_;
  assign new_n52722_ = \b[58]  & ~new_n52714_;
  assign new_n52723_ = ~new_n52719_ & new_n52722_;
  assign new_n52724_ = new_n24707_ & ~new_n52723_;
  assign new_n52725_ = ~new_n52721_ & new_n52724_;
  assign new_n52726_ = ~new_n52713_ & new_n52725_;
  assign new_n52727_ = new_n23895_ & ~new_n52720_;
  assign new_n52728_ = ~new_n52726_ & ~new_n52727_;
  assign new_n52729_ = ~new_n51937_ & new_n52711_;
  assign new_n52730_ = ~new_n52707_ & new_n52729_;
  assign new_n52731_ = ~new_n52708_ & ~new_n52711_;
  assign new_n52732_ = ~new_n52730_ & ~new_n52731_;
  assign new_n52733_ = ~new_n52728_ & ~new_n52732_;
  assign new_n52734_ = ~new_n51927_ & ~new_n52727_;
  assign new_n52735_ = ~new_n52726_ & new_n52734_;
  assign new_n52736_ = ~new_n52733_ & ~new_n52735_;
  assign new_n52737_ = ~\b[58]  & ~new_n52736_;
  assign new_n52738_ = ~new_n51946_ & new_n52706_;
  assign new_n52739_ = ~new_n52702_ & new_n52738_;
  assign new_n52740_ = ~new_n52703_ & ~new_n52706_;
  assign new_n52741_ = ~new_n52739_ & ~new_n52740_;
  assign new_n52742_ = ~new_n52728_ & ~new_n52741_;
  assign new_n52743_ = ~new_n51936_ & ~new_n52727_;
  assign new_n52744_ = ~new_n52726_ & new_n52743_;
  assign new_n52745_ = ~new_n52742_ & ~new_n52744_;
  assign new_n52746_ = ~\b[57]  & ~new_n52745_;
  assign new_n52747_ = ~new_n51955_ & new_n52701_;
  assign new_n52748_ = ~new_n52697_ & new_n52747_;
  assign new_n52749_ = ~new_n52698_ & ~new_n52701_;
  assign new_n52750_ = ~new_n52748_ & ~new_n52749_;
  assign new_n52751_ = ~new_n52728_ & ~new_n52750_;
  assign new_n52752_ = ~new_n51945_ & ~new_n52727_;
  assign new_n52753_ = ~new_n52726_ & new_n52752_;
  assign new_n52754_ = ~new_n52751_ & ~new_n52753_;
  assign new_n52755_ = ~\b[56]  & ~new_n52754_;
  assign new_n52756_ = ~new_n51964_ & new_n52696_;
  assign new_n52757_ = ~new_n52692_ & new_n52756_;
  assign new_n52758_ = ~new_n52693_ & ~new_n52696_;
  assign new_n52759_ = ~new_n52757_ & ~new_n52758_;
  assign new_n52760_ = ~new_n52728_ & ~new_n52759_;
  assign new_n52761_ = ~new_n51954_ & ~new_n52727_;
  assign new_n52762_ = ~new_n52726_ & new_n52761_;
  assign new_n52763_ = ~new_n52760_ & ~new_n52762_;
  assign new_n52764_ = ~\b[55]  & ~new_n52763_;
  assign new_n52765_ = ~new_n51973_ & new_n52691_;
  assign new_n52766_ = ~new_n52687_ & new_n52765_;
  assign new_n52767_ = ~new_n52688_ & ~new_n52691_;
  assign new_n52768_ = ~new_n52766_ & ~new_n52767_;
  assign new_n52769_ = ~new_n52728_ & ~new_n52768_;
  assign new_n52770_ = ~new_n51963_ & ~new_n52727_;
  assign new_n52771_ = ~new_n52726_ & new_n52770_;
  assign new_n52772_ = ~new_n52769_ & ~new_n52771_;
  assign new_n52773_ = ~\b[54]  & ~new_n52772_;
  assign new_n52774_ = ~new_n51982_ & new_n52686_;
  assign new_n52775_ = ~new_n52682_ & new_n52774_;
  assign new_n52776_ = ~new_n52683_ & ~new_n52686_;
  assign new_n52777_ = ~new_n52775_ & ~new_n52776_;
  assign new_n52778_ = ~new_n52728_ & ~new_n52777_;
  assign new_n52779_ = ~new_n51972_ & ~new_n52727_;
  assign new_n52780_ = ~new_n52726_ & new_n52779_;
  assign new_n52781_ = ~new_n52778_ & ~new_n52780_;
  assign new_n52782_ = ~\b[53]  & ~new_n52781_;
  assign new_n52783_ = ~new_n51991_ & new_n52681_;
  assign new_n52784_ = ~new_n52677_ & new_n52783_;
  assign new_n52785_ = ~new_n52678_ & ~new_n52681_;
  assign new_n52786_ = ~new_n52784_ & ~new_n52785_;
  assign new_n52787_ = ~new_n52728_ & ~new_n52786_;
  assign new_n52788_ = ~new_n51981_ & ~new_n52727_;
  assign new_n52789_ = ~new_n52726_ & new_n52788_;
  assign new_n52790_ = ~new_n52787_ & ~new_n52789_;
  assign new_n52791_ = ~\b[52]  & ~new_n52790_;
  assign new_n52792_ = ~new_n52000_ & new_n52676_;
  assign new_n52793_ = ~new_n52672_ & new_n52792_;
  assign new_n52794_ = ~new_n52673_ & ~new_n52676_;
  assign new_n52795_ = ~new_n52793_ & ~new_n52794_;
  assign new_n52796_ = ~new_n52728_ & ~new_n52795_;
  assign new_n52797_ = ~new_n51990_ & ~new_n52727_;
  assign new_n52798_ = ~new_n52726_ & new_n52797_;
  assign new_n52799_ = ~new_n52796_ & ~new_n52798_;
  assign new_n52800_ = ~\b[51]  & ~new_n52799_;
  assign new_n52801_ = ~new_n52009_ & new_n52671_;
  assign new_n52802_ = ~new_n52667_ & new_n52801_;
  assign new_n52803_ = ~new_n52668_ & ~new_n52671_;
  assign new_n52804_ = ~new_n52802_ & ~new_n52803_;
  assign new_n52805_ = ~new_n52728_ & ~new_n52804_;
  assign new_n52806_ = ~new_n51999_ & ~new_n52727_;
  assign new_n52807_ = ~new_n52726_ & new_n52806_;
  assign new_n52808_ = ~new_n52805_ & ~new_n52807_;
  assign new_n52809_ = ~\b[50]  & ~new_n52808_;
  assign new_n52810_ = ~new_n52018_ & new_n52666_;
  assign new_n52811_ = ~new_n52662_ & new_n52810_;
  assign new_n52812_ = ~new_n52663_ & ~new_n52666_;
  assign new_n52813_ = ~new_n52811_ & ~new_n52812_;
  assign new_n52814_ = ~new_n52728_ & ~new_n52813_;
  assign new_n52815_ = ~new_n52008_ & ~new_n52727_;
  assign new_n52816_ = ~new_n52726_ & new_n52815_;
  assign new_n52817_ = ~new_n52814_ & ~new_n52816_;
  assign new_n52818_ = ~\b[49]  & ~new_n52817_;
  assign new_n52819_ = ~new_n52027_ & new_n52661_;
  assign new_n52820_ = ~new_n52657_ & new_n52819_;
  assign new_n52821_ = ~new_n52658_ & ~new_n52661_;
  assign new_n52822_ = ~new_n52820_ & ~new_n52821_;
  assign new_n52823_ = ~new_n52728_ & ~new_n52822_;
  assign new_n52824_ = ~new_n52017_ & ~new_n52727_;
  assign new_n52825_ = ~new_n52726_ & new_n52824_;
  assign new_n52826_ = ~new_n52823_ & ~new_n52825_;
  assign new_n52827_ = ~\b[48]  & ~new_n52826_;
  assign new_n52828_ = ~new_n52036_ & new_n52656_;
  assign new_n52829_ = ~new_n52652_ & new_n52828_;
  assign new_n52830_ = ~new_n52653_ & ~new_n52656_;
  assign new_n52831_ = ~new_n52829_ & ~new_n52830_;
  assign new_n52832_ = ~new_n52728_ & ~new_n52831_;
  assign new_n52833_ = ~new_n52026_ & ~new_n52727_;
  assign new_n52834_ = ~new_n52726_ & new_n52833_;
  assign new_n52835_ = ~new_n52832_ & ~new_n52834_;
  assign new_n52836_ = ~\b[47]  & ~new_n52835_;
  assign new_n52837_ = ~new_n52045_ & new_n52651_;
  assign new_n52838_ = ~new_n52647_ & new_n52837_;
  assign new_n52839_ = ~new_n52648_ & ~new_n52651_;
  assign new_n52840_ = ~new_n52838_ & ~new_n52839_;
  assign new_n52841_ = ~new_n52728_ & ~new_n52840_;
  assign new_n52842_ = ~new_n52035_ & ~new_n52727_;
  assign new_n52843_ = ~new_n52726_ & new_n52842_;
  assign new_n52844_ = ~new_n52841_ & ~new_n52843_;
  assign new_n52845_ = ~\b[46]  & ~new_n52844_;
  assign new_n52846_ = ~new_n52054_ & new_n52646_;
  assign new_n52847_ = ~new_n52642_ & new_n52846_;
  assign new_n52848_ = ~new_n52643_ & ~new_n52646_;
  assign new_n52849_ = ~new_n52847_ & ~new_n52848_;
  assign new_n52850_ = ~new_n52728_ & ~new_n52849_;
  assign new_n52851_ = ~new_n52044_ & ~new_n52727_;
  assign new_n52852_ = ~new_n52726_ & new_n52851_;
  assign new_n52853_ = ~new_n52850_ & ~new_n52852_;
  assign new_n52854_ = ~\b[45]  & ~new_n52853_;
  assign new_n52855_ = ~new_n52063_ & new_n52641_;
  assign new_n52856_ = ~new_n52637_ & new_n52855_;
  assign new_n52857_ = ~new_n52638_ & ~new_n52641_;
  assign new_n52858_ = ~new_n52856_ & ~new_n52857_;
  assign new_n52859_ = ~new_n52728_ & ~new_n52858_;
  assign new_n52860_ = ~new_n52053_ & ~new_n52727_;
  assign new_n52861_ = ~new_n52726_ & new_n52860_;
  assign new_n52862_ = ~new_n52859_ & ~new_n52861_;
  assign new_n52863_ = ~\b[44]  & ~new_n52862_;
  assign new_n52864_ = ~new_n52072_ & new_n52636_;
  assign new_n52865_ = ~new_n52632_ & new_n52864_;
  assign new_n52866_ = ~new_n52633_ & ~new_n52636_;
  assign new_n52867_ = ~new_n52865_ & ~new_n52866_;
  assign new_n52868_ = ~new_n52728_ & ~new_n52867_;
  assign new_n52869_ = ~new_n52062_ & ~new_n52727_;
  assign new_n52870_ = ~new_n52726_ & new_n52869_;
  assign new_n52871_ = ~new_n52868_ & ~new_n52870_;
  assign new_n52872_ = ~\b[43]  & ~new_n52871_;
  assign new_n52873_ = ~new_n52081_ & new_n52631_;
  assign new_n52874_ = ~new_n52627_ & new_n52873_;
  assign new_n52875_ = ~new_n52628_ & ~new_n52631_;
  assign new_n52876_ = ~new_n52874_ & ~new_n52875_;
  assign new_n52877_ = ~new_n52728_ & ~new_n52876_;
  assign new_n52878_ = ~new_n52071_ & ~new_n52727_;
  assign new_n52879_ = ~new_n52726_ & new_n52878_;
  assign new_n52880_ = ~new_n52877_ & ~new_n52879_;
  assign new_n52881_ = ~\b[42]  & ~new_n52880_;
  assign new_n52882_ = ~new_n52090_ & new_n52626_;
  assign new_n52883_ = ~new_n52622_ & new_n52882_;
  assign new_n52884_ = ~new_n52623_ & ~new_n52626_;
  assign new_n52885_ = ~new_n52883_ & ~new_n52884_;
  assign new_n52886_ = ~new_n52728_ & ~new_n52885_;
  assign new_n52887_ = ~new_n52080_ & ~new_n52727_;
  assign new_n52888_ = ~new_n52726_ & new_n52887_;
  assign new_n52889_ = ~new_n52886_ & ~new_n52888_;
  assign new_n52890_ = ~\b[41]  & ~new_n52889_;
  assign new_n52891_ = ~new_n52099_ & new_n52621_;
  assign new_n52892_ = ~new_n52617_ & new_n52891_;
  assign new_n52893_ = ~new_n52618_ & ~new_n52621_;
  assign new_n52894_ = ~new_n52892_ & ~new_n52893_;
  assign new_n52895_ = ~new_n52728_ & ~new_n52894_;
  assign new_n52896_ = ~new_n52089_ & ~new_n52727_;
  assign new_n52897_ = ~new_n52726_ & new_n52896_;
  assign new_n52898_ = ~new_n52895_ & ~new_n52897_;
  assign new_n52899_ = ~\b[40]  & ~new_n52898_;
  assign new_n52900_ = ~new_n52108_ & new_n52616_;
  assign new_n52901_ = ~new_n52612_ & new_n52900_;
  assign new_n52902_ = ~new_n52613_ & ~new_n52616_;
  assign new_n52903_ = ~new_n52901_ & ~new_n52902_;
  assign new_n52904_ = ~new_n52728_ & ~new_n52903_;
  assign new_n52905_ = ~new_n52098_ & ~new_n52727_;
  assign new_n52906_ = ~new_n52726_ & new_n52905_;
  assign new_n52907_ = ~new_n52904_ & ~new_n52906_;
  assign new_n52908_ = ~\b[39]  & ~new_n52907_;
  assign new_n52909_ = ~new_n52117_ & new_n52611_;
  assign new_n52910_ = ~new_n52607_ & new_n52909_;
  assign new_n52911_ = ~new_n52608_ & ~new_n52611_;
  assign new_n52912_ = ~new_n52910_ & ~new_n52911_;
  assign new_n52913_ = ~new_n52728_ & ~new_n52912_;
  assign new_n52914_ = ~new_n52107_ & ~new_n52727_;
  assign new_n52915_ = ~new_n52726_ & new_n52914_;
  assign new_n52916_ = ~new_n52913_ & ~new_n52915_;
  assign new_n52917_ = ~\b[38]  & ~new_n52916_;
  assign new_n52918_ = ~new_n52126_ & new_n52606_;
  assign new_n52919_ = ~new_n52602_ & new_n52918_;
  assign new_n52920_ = ~new_n52603_ & ~new_n52606_;
  assign new_n52921_ = ~new_n52919_ & ~new_n52920_;
  assign new_n52922_ = ~new_n52728_ & ~new_n52921_;
  assign new_n52923_ = ~new_n52116_ & ~new_n52727_;
  assign new_n52924_ = ~new_n52726_ & new_n52923_;
  assign new_n52925_ = ~new_n52922_ & ~new_n52924_;
  assign new_n52926_ = ~\b[37]  & ~new_n52925_;
  assign new_n52927_ = ~new_n52135_ & new_n52601_;
  assign new_n52928_ = ~new_n52597_ & new_n52927_;
  assign new_n52929_ = ~new_n52598_ & ~new_n52601_;
  assign new_n52930_ = ~new_n52928_ & ~new_n52929_;
  assign new_n52931_ = ~new_n52728_ & ~new_n52930_;
  assign new_n52932_ = ~new_n52125_ & ~new_n52727_;
  assign new_n52933_ = ~new_n52726_ & new_n52932_;
  assign new_n52934_ = ~new_n52931_ & ~new_n52933_;
  assign new_n52935_ = ~\b[36]  & ~new_n52934_;
  assign new_n52936_ = ~new_n52144_ & new_n52596_;
  assign new_n52937_ = ~new_n52592_ & new_n52936_;
  assign new_n52938_ = ~new_n52593_ & ~new_n52596_;
  assign new_n52939_ = ~new_n52937_ & ~new_n52938_;
  assign new_n52940_ = ~new_n52728_ & ~new_n52939_;
  assign new_n52941_ = ~new_n52134_ & ~new_n52727_;
  assign new_n52942_ = ~new_n52726_ & new_n52941_;
  assign new_n52943_ = ~new_n52940_ & ~new_n52942_;
  assign new_n52944_ = ~\b[35]  & ~new_n52943_;
  assign new_n52945_ = ~new_n52153_ & new_n52591_;
  assign new_n52946_ = ~new_n52587_ & new_n52945_;
  assign new_n52947_ = ~new_n52588_ & ~new_n52591_;
  assign new_n52948_ = ~new_n52946_ & ~new_n52947_;
  assign new_n52949_ = ~new_n52728_ & ~new_n52948_;
  assign new_n52950_ = ~new_n52143_ & ~new_n52727_;
  assign new_n52951_ = ~new_n52726_ & new_n52950_;
  assign new_n52952_ = ~new_n52949_ & ~new_n52951_;
  assign new_n52953_ = ~\b[34]  & ~new_n52952_;
  assign new_n52954_ = ~new_n52162_ & new_n52586_;
  assign new_n52955_ = ~new_n52582_ & new_n52954_;
  assign new_n52956_ = ~new_n52583_ & ~new_n52586_;
  assign new_n52957_ = ~new_n52955_ & ~new_n52956_;
  assign new_n52958_ = ~new_n52728_ & ~new_n52957_;
  assign new_n52959_ = ~new_n52152_ & ~new_n52727_;
  assign new_n52960_ = ~new_n52726_ & new_n52959_;
  assign new_n52961_ = ~new_n52958_ & ~new_n52960_;
  assign new_n52962_ = ~\b[33]  & ~new_n52961_;
  assign new_n52963_ = ~new_n52171_ & new_n52581_;
  assign new_n52964_ = ~new_n52577_ & new_n52963_;
  assign new_n52965_ = ~new_n52578_ & ~new_n52581_;
  assign new_n52966_ = ~new_n52964_ & ~new_n52965_;
  assign new_n52967_ = ~new_n52728_ & ~new_n52966_;
  assign new_n52968_ = ~new_n52161_ & ~new_n52727_;
  assign new_n52969_ = ~new_n52726_ & new_n52968_;
  assign new_n52970_ = ~new_n52967_ & ~new_n52969_;
  assign new_n52971_ = ~\b[32]  & ~new_n52970_;
  assign new_n52972_ = ~new_n52180_ & new_n52576_;
  assign new_n52973_ = ~new_n52572_ & new_n52972_;
  assign new_n52974_ = ~new_n52573_ & ~new_n52576_;
  assign new_n52975_ = ~new_n52973_ & ~new_n52974_;
  assign new_n52976_ = ~new_n52728_ & ~new_n52975_;
  assign new_n52977_ = ~new_n52170_ & ~new_n52727_;
  assign new_n52978_ = ~new_n52726_ & new_n52977_;
  assign new_n52979_ = ~new_n52976_ & ~new_n52978_;
  assign new_n52980_ = ~\b[31]  & ~new_n52979_;
  assign new_n52981_ = ~new_n52189_ & new_n52571_;
  assign new_n52982_ = ~new_n52567_ & new_n52981_;
  assign new_n52983_ = ~new_n52568_ & ~new_n52571_;
  assign new_n52984_ = ~new_n52982_ & ~new_n52983_;
  assign new_n52985_ = ~new_n52728_ & ~new_n52984_;
  assign new_n52986_ = ~new_n52179_ & ~new_n52727_;
  assign new_n52987_ = ~new_n52726_ & new_n52986_;
  assign new_n52988_ = ~new_n52985_ & ~new_n52987_;
  assign new_n52989_ = ~\b[30]  & ~new_n52988_;
  assign new_n52990_ = ~new_n52198_ & new_n52566_;
  assign new_n52991_ = ~new_n52562_ & new_n52990_;
  assign new_n52992_ = ~new_n52563_ & ~new_n52566_;
  assign new_n52993_ = ~new_n52991_ & ~new_n52992_;
  assign new_n52994_ = ~new_n52728_ & ~new_n52993_;
  assign new_n52995_ = ~new_n52188_ & ~new_n52727_;
  assign new_n52996_ = ~new_n52726_ & new_n52995_;
  assign new_n52997_ = ~new_n52994_ & ~new_n52996_;
  assign new_n52998_ = ~\b[29]  & ~new_n52997_;
  assign new_n52999_ = ~new_n52207_ & new_n52561_;
  assign new_n53000_ = ~new_n52557_ & new_n52999_;
  assign new_n53001_ = ~new_n52558_ & ~new_n52561_;
  assign new_n53002_ = ~new_n53000_ & ~new_n53001_;
  assign new_n53003_ = ~new_n52728_ & ~new_n53002_;
  assign new_n53004_ = ~new_n52197_ & ~new_n52727_;
  assign new_n53005_ = ~new_n52726_ & new_n53004_;
  assign new_n53006_ = ~new_n53003_ & ~new_n53005_;
  assign new_n53007_ = ~\b[28]  & ~new_n53006_;
  assign new_n53008_ = ~new_n52216_ & new_n52556_;
  assign new_n53009_ = ~new_n52552_ & new_n53008_;
  assign new_n53010_ = ~new_n52553_ & ~new_n52556_;
  assign new_n53011_ = ~new_n53009_ & ~new_n53010_;
  assign new_n53012_ = ~new_n52728_ & ~new_n53011_;
  assign new_n53013_ = ~new_n52206_ & ~new_n52727_;
  assign new_n53014_ = ~new_n52726_ & new_n53013_;
  assign new_n53015_ = ~new_n53012_ & ~new_n53014_;
  assign new_n53016_ = ~\b[27]  & ~new_n53015_;
  assign new_n53017_ = ~new_n52225_ & new_n52551_;
  assign new_n53018_ = ~new_n52547_ & new_n53017_;
  assign new_n53019_ = ~new_n52548_ & ~new_n52551_;
  assign new_n53020_ = ~new_n53018_ & ~new_n53019_;
  assign new_n53021_ = ~new_n52728_ & ~new_n53020_;
  assign new_n53022_ = ~new_n52215_ & ~new_n52727_;
  assign new_n53023_ = ~new_n52726_ & new_n53022_;
  assign new_n53024_ = ~new_n53021_ & ~new_n53023_;
  assign new_n53025_ = ~\b[26]  & ~new_n53024_;
  assign new_n53026_ = ~new_n52234_ & new_n52546_;
  assign new_n53027_ = ~new_n52542_ & new_n53026_;
  assign new_n53028_ = ~new_n52543_ & ~new_n52546_;
  assign new_n53029_ = ~new_n53027_ & ~new_n53028_;
  assign new_n53030_ = ~new_n52728_ & ~new_n53029_;
  assign new_n53031_ = ~new_n52224_ & ~new_n52727_;
  assign new_n53032_ = ~new_n52726_ & new_n53031_;
  assign new_n53033_ = ~new_n53030_ & ~new_n53032_;
  assign new_n53034_ = ~\b[25]  & ~new_n53033_;
  assign new_n53035_ = ~new_n52243_ & new_n52541_;
  assign new_n53036_ = ~new_n52537_ & new_n53035_;
  assign new_n53037_ = ~new_n52538_ & ~new_n52541_;
  assign new_n53038_ = ~new_n53036_ & ~new_n53037_;
  assign new_n53039_ = ~new_n52728_ & ~new_n53038_;
  assign new_n53040_ = ~new_n52233_ & ~new_n52727_;
  assign new_n53041_ = ~new_n52726_ & new_n53040_;
  assign new_n53042_ = ~new_n53039_ & ~new_n53041_;
  assign new_n53043_ = ~\b[24]  & ~new_n53042_;
  assign new_n53044_ = ~new_n52252_ & new_n52536_;
  assign new_n53045_ = ~new_n52532_ & new_n53044_;
  assign new_n53046_ = ~new_n52533_ & ~new_n52536_;
  assign new_n53047_ = ~new_n53045_ & ~new_n53046_;
  assign new_n53048_ = ~new_n52728_ & ~new_n53047_;
  assign new_n53049_ = ~new_n52242_ & ~new_n52727_;
  assign new_n53050_ = ~new_n52726_ & new_n53049_;
  assign new_n53051_ = ~new_n53048_ & ~new_n53050_;
  assign new_n53052_ = ~\b[23]  & ~new_n53051_;
  assign new_n53053_ = ~new_n52261_ & new_n52531_;
  assign new_n53054_ = ~new_n52527_ & new_n53053_;
  assign new_n53055_ = ~new_n52528_ & ~new_n52531_;
  assign new_n53056_ = ~new_n53054_ & ~new_n53055_;
  assign new_n53057_ = ~new_n52728_ & ~new_n53056_;
  assign new_n53058_ = ~new_n52251_ & ~new_n52727_;
  assign new_n53059_ = ~new_n52726_ & new_n53058_;
  assign new_n53060_ = ~new_n53057_ & ~new_n53059_;
  assign new_n53061_ = ~\b[22]  & ~new_n53060_;
  assign new_n53062_ = ~new_n52270_ & new_n52526_;
  assign new_n53063_ = ~new_n52522_ & new_n53062_;
  assign new_n53064_ = ~new_n52523_ & ~new_n52526_;
  assign new_n53065_ = ~new_n53063_ & ~new_n53064_;
  assign new_n53066_ = ~new_n52728_ & ~new_n53065_;
  assign new_n53067_ = ~new_n52260_ & ~new_n52727_;
  assign new_n53068_ = ~new_n52726_ & new_n53067_;
  assign new_n53069_ = ~new_n53066_ & ~new_n53068_;
  assign new_n53070_ = ~\b[21]  & ~new_n53069_;
  assign new_n53071_ = ~new_n52279_ & new_n52521_;
  assign new_n53072_ = ~new_n52517_ & new_n53071_;
  assign new_n53073_ = ~new_n52518_ & ~new_n52521_;
  assign new_n53074_ = ~new_n53072_ & ~new_n53073_;
  assign new_n53075_ = ~new_n52728_ & ~new_n53074_;
  assign new_n53076_ = ~new_n52269_ & ~new_n52727_;
  assign new_n53077_ = ~new_n52726_ & new_n53076_;
  assign new_n53078_ = ~new_n53075_ & ~new_n53077_;
  assign new_n53079_ = ~\b[20]  & ~new_n53078_;
  assign new_n53080_ = ~new_n52288_ & new_n52516_;
  assign new_n53081_ = ~new_n52512_ & new_n53080_;
  assign new_n53082_ = ~new_n52513_ & ~new_n52516_;
  assign new_n53083_ = ~new_n53081_ & ~new_n53082_;
  assign new_n53084_ = ~new_n52728_ & ~new_n53083_;
  assign new_n53085_ = ~new_n52278_ & ~new_n52727_;
  assign new_n53086_ = ~new_n52726_ & new_n53085_;
  assign new_n53087_ = ~new_n53084_ & ~new_n53086_;
  assign new_n53088_ = ~\b[19]  & ~new_n53087_;
  assign new_n53089_ = ~new_n52297_ & new_n52511_;
  assign new_n53090_ = ~new_n52507_ & new_n53089_;
  assign new_n53091_ = ~new_n52508_ & ~new_n52511_;
  assign new_n53092_ = ~new_n53090_ & ~new_n53091_;
  assign new_n53093_ = ~new_n52728_ & ~new_n53092_;
  assign new_n53094_ = ~new_n52287_ & ~new_n52727_;
  assign new_n53095_ = ~new_n52726_ & new_n53094_;
  assign new_n53096_ = ~new_n53093_ & ~new_n53095_;
  assign new_n53097_ = ~\b[18]  & ~new_n53096_;
  assign new_n53098_ = ~new_n52306_ & new_n52506_;
  assign new_n53099_ = ~new_n52502_ & new_n53098_;
  assign new_n53100_ = ~new_n52503_ & ~new_n52506_;
  assign new_n53101_ = ~new_n53099_ & ~new_n53100_;
  assign new_n53102_ = ~new_n52728_ & ~new_n53101_;
  assign new_n53103_ = ~new_n52296_ & ~new_n52727_;
  assign new_n53104_ = ~new_n52726_ & new_n53103_;
  assign new_n53105_ = ~new_n53102_ & ~new_n53104_;
  assign new_n53106_ = ~\b[17]  & ~new_n53105_;
  assign new_n53107_ = ~new_n52315_ & new_n52501_;
  assign new_n53108_ = ~new_n52497_ & new_n53107_;
  assign new_n53109_ = ~new_n52498_ & ~new_n52501_;
  assign new_n53110_ = ~new_n53108_ & ~new_n53109_;
  assign new_n53111_ = ~new_n52728_ & ~new_n53110_;
  assign new_n53112_ = ~new_n52305_ & ~new_n52727_;
  assign new_n53113_ = ~new_n52726_ & new_n53112_;
  assign new_n53114_ = ~new_n53111_ & ~new_n53113_;
  assign new_n53115_ = ~\b[16]  & ~new_n53114_;
  assign new_n53116_ = ~new_n52324_ & new_n52496_;
  assign new_n53117_ = ~new_n52492_ & new_n53116_;
  assign new_n53118_ = ~new_n52493_ & ~new_n52496_;
  assign new_n53119_ = ~new_n53117_ & ~new_n53118_;
  assign new_n53120_ = ~new_n52728_ & ~new_n53119_;
  assign new_n53121_ = ~new_n52314_ & ~new_n52727_;
  assign new_n53122_ = ~new_n52726_ & new_n53121_;
  assign new_n53123_ = ~new_n53120_ & ~new_n53122_;
  assign new_n53124_ = ~\b[15]  & ~new_n53123_;
  assign new_n53125_ = ~new_n52333_ & new_n52491_;
  assign new_n53126_ = ~new_n52487_ & new_n53125_;
  assign new_n53127_ = ~new_n52488_ & ~new_n52491_;
  assign new_n53128_ = ~new_n53126_ & ~new_n53127_;
  assign new_n53129_ = ~new_n52728_ & ~new_n53128_;
  assign new_n53130_ = ~new_n52323_ & ~new_n52727_;
  assign new_n53131_ = ~new_n52726_ & new_n53130_;
  assign new_n53132_ = ~new_n53129_ & ~new_n53131_;
  assign new_n53133_ = ~\b[14]  & ~new_n53132_;
  assign new_n53134_ = ~new_n52342_ & new_n52486_;
  assign new_n53135_ = ~new_n52482_ & new_n53134_;
  assign new_n53136_ = ~new_n52483_ & ~new_n52486_;
  assign new_n53137_ = ~new_n53135_ & ~new_n53136_;
  assign new_n53138_ = ~new_n52728_ & ~new_n53137_;
  assign new_n53139_ = ~new_n52332_ & ~new_n52727_;
  assign new_n53140_ = ~new_n52726_ & new_n53139_;
  assign new_n53141_ = ~new_n53138_ & ~new_n53140_;
  assign new_n53142_ = ~\b[13]  & ~new_n53141_;
  assign new_n53143_ = ~new_n52351_ & new_n52481_;
  assign new_n53144_ = ~new_n52477_ & new_n53143_;
  assign new_n53145_ = ~new_n52478_ & ~new_n52481_;
  assign new_n53146_ = ~new_n53144_ & ~new_n53145_;
  assign new_n53147_ = ~new_n52728_ & ~new_n53146_;
  assign new_n53148_ = ~new_n52341_ & ~new_n52727_;
  assign new_n53149_ = ~new_n52726_ & new_n53148_;
  assign new_n53150_ = ~new_n53147_ & ~new_n53149_;
  assign new_n53151_ = ~\b[12]  & ~new_n53150_;
  assign new_n53152_ = ~new_n52360_ & new_n52476_;
  assign new_n53153_ = ~new_n52472_ & new_n53152_;
  assign new_n53154_ = ~new_n52473_ & ~new_n52476_;
  assign new_n53155_ = ~new_n53153_ & ~new_n53154_;
  assign new_n53156_ = ~new_n52728_ & ~new_n53155_;
  assign new_n53157_ = ~new_n52350_ & ~new_n52727_;
  assign new_n53158_ = ~new_n52726_ & new_n53157_;
  assign new_n53159_ = ~new_n53156_ & ~new_n53158_;
  assign new_n53160_ = ~\b[11]  & ~new_n53159_;
  assign new_n53161_ = ~new_n52369_ & new_n52471_;
  assign new_n53162_ = ~new_n52467_ & new_n53161_;
  assign new_n53163_ = ~new_n52468_ & ~new_n52471_;
  assign new_n53164_ = ~new_n53162_ & ~new_n53163_;
  assign new_n53165_ = ~new_n52728_ & ~new_n53164_;
  assign new_n53166_ = ~new_n52359_ & ~new_n52727_;
  assign new_n53167_ = ~new_n52726_ & new_n53166_;
  assign new_n53168_ = ~new_n53165_ & ~new_n53167_;
  assign new_n53169_ = ~\b[10]  & ~new_n53168_;
  assign new_n53170_ = ~new_n52378_ & new_n52466_;
  assign new_n53171_ = ~new_n52462_ & new_n53170_;
  assign new_n53172_ = ~new_n52463_ & ~new_n52466_;
  assign new_n53173_ = ~new_n53171_ & ~new_n53172_;
  assign new_n53174_ = ~new_n52728_ & ~new_n53173_;
  assign new_n53175_ = ~new_n52368_ & ~new_n52727_;
  assign new_n53176_ = ~new_n52726_ & new_n53175_;
  assign new_n53177_ = ~new_n53174_ & ~new_n53176_;
  assign new_n53178_ = ~\b[9]  & ~new_n53177_;
  assign new_n53179_ = ~new_n52387_ & new_n52461_;
  assign new_n53180_ = ~new_n52457_ & new_n53179_;
  assign new_n53181_ = ~new_n52458_ & ~new_n52461_;
  assign new_n53182_ = ~new_n53180_ & ~new_n53181_;
  assign new_n53183_ = ~new_n52728_ & ~new_n53182_;
  assign new_n53184_ = ~new_n52377_ & ~new_n52727_;
  assign new_n53185_ = ~new_n52726_ & new_n53184_;
  assign new_n53186_ = ~new_n53183_ & ~new_n53185_;
  assign new_n53187_ = ~\b[8]  & ~new_n53186_;
  assign new_n53188_ = ~new_n52396_ & new_n52456_;
  assign new_n53189_ = ~new_n52452_ & new_n53188_;
  assign new_n53190_ = ~new_n52453_ & ~new_n52456_;
  assign new_n53191_ = ~new_n53189_ & ~new_n53190_;
  assign new_n53192_ = ~new_n52728_ & ~new_n53191_;
  assign new_n53193_ = ~new_n52386_ & ~new_n52727_;
  assign new_n53194_ = ~new_n52726_ & new_n53193_;
  assign new_n53195_ = ~new_n53192_ & ~new_n53194_;
  assign new_n53196_ = ~\b[7]  & ~new_n53195_;
  assign new_n53197_ = ~new_n52405_ & new_n52451_;
  assign new_n53198_ = ~new_n52447_ & new_n53197_;
  assign new_n53199_ = ~new_n52448_ & ~new_n52451_;
  assign new_n53200_ = ~new_n53198_ & ~new_n53199_;
  assign new_n53201_ = ~new_n52728_ & ~new_n53200_;
  assign new_n53202_ = ~new_n52395_ & ~new_n52727_;
  assign new_n53203_ = ~new_n52726_ & new_n53202_;
  assign new_n53204_ = ~new_n53201_ & ~new_n53203_;
  assign new_n53205_ = ~\b[6]  & ~new_n53204_;
  assign new_n53206_ = ~new_n52414_ & new_n52446_;
  assign new_n53207_ = ~new_n52442_ & new_n53206_;
  assign new_n53208_ = ~new_n52443_ & ~new_n52446_;
  assign new_n53209_ = ~new_n53207_ & ~new_n53208_;
  assign new_n53210_ = ~new_n52728_ & ~new_n53209_;
  assign new_n53211_ = ~new_n52404_ & ~new_n52727_;
  assign new_n53212_ = ~new_n52726_ & new_n53211_;
  assign new_n53213_ = ~new_n53210_ & ~new_n53212_;
  assign new_n53214_ = ~\b[5]  & ~new_n53213_;
  assign new_n53215_ = ~new_n52422_ & new_n52441_;
  assign new_n53216_ = ~new_n52437_ & new_n53215_;
  assign new_n53217_ = ~new_n52438_ & ~new_n52441_;
  assign new_n53218_ = ~new_n53216_ & ~new_n53217_;
  assign new_n53219_ = ~new_n52728_ & ~new_n53218_;
  assign new_n53220_ = ~new_n52413_ & ~new_n52727_;
  assign new_n53221_ = ~new_n52726_ & new_n53220_;
  assign new_n53222_ = ~new_n53219_ & ~new_n53221_;
  assign new_n53223_ = ~\b[4]  & ~new_n53222_;
  assign new_n53224_ = ~new_n52432_ & new_n52436_;
  assign new_n53225_ = ~new_n52431_ & new_n53224_;
  assign new_n53226_ = ~new_n52433_ & ~new_n52436_;
  assign new_n53227_ = ~new_n53225_ & ~new_n53226_;
  assign new_n53228_ = ~new_n52728_ & ~new_n53227_;
  assign new_n53229_ = ~new_n52421_ & ~new_n52727_;
  assign new_n53230_ = ~new_n52726_ & new_n53229_;
  assign new_n53231_ = ~new_n53228_ & ~new_n53230_;
  assign new_n53232_ = ~\b[3]  & ~new_n53231_;
  assign new_n53233_ = new_n24413_ & ~new_n52429_;
  assign new_n53234_ = ~new_n52427_ & new_n53233_;
  assign new_n53235_ = ~new_n52431_ & ~new_n53234_;
  assign new_n53236_ = ~new_n52728_ & new_n53235_;
  assign new_n53237_ = ~new_n52426_ & ~new_n52727_;
  assign new_n53238_ = ~new_n52726_ & new_n53237_;
  assign new_n53239_ = ~new_n53236_ & ~new_n53238_;
  assign new_n53240_ = ~\b[2]  & ~new_n53239_;
  assign new_n53241_ = \b[0]  & ~new_n52728_;
  assign new_n53242_ = \a[5]  & ~new_n53241_;
  assign new_n53243_ = new_n24413_ & ~new_n52728_;
  assign new_n53244_ = ~new_n53242_ & ~new_n53243_;
  assign new_n53245_ = \b[1]  & ~new_n53244_;
  assign new_n53246_ = ~\b[1]  & ~new_n53243_;
  assign new_n53247_ = ~new_n53242_ & new_n53246_;
  assign new_n53248_ = ~new_n53245_ & ~new_n53247_;
  assign new_n53249_ = ~new_n25233_ & ~new_n53248_;
  assign new_n53250_ = ~\b[1]  & ~new_n53244_;
  assign new_n53251_ = ~new_n53249_ & ~new_n53250_;
  assign new_n53252_ = \b[2]  & ~new_n53238_;
  assign new_n53253_ = ~new_n53236_ & new_n53252_;
  assign new_n53254_ = ~new_n53240_ & ~new_n53253_;
  assign new_n53255_ = ~new_n53251_ & new_n53254_;
  assign new_n53256_ = ~new_n53240_ & ~new_n53255_;
  assign new_n53257_ = \b[3]  & ~new_n53230_;
  assign new_n53258_ = ~new_n53228_ & new_n53257_;
  assign new_n53259_ = ~new_n53232_ & ~new_n53258_;
  assign new_n53260_ = ~new_n53256_ & new_n53259_;
  assign new_n53261_ = ~new_n53232_ & ~new_n53260_;
  assign new_n53262_ = \b[4]  & ~new_n53221_;
  assign new_n53263_ = ~new_n53219_ & new_n53262_;
  assign new_n53264_ = ~new_n53223_ & ~new_n53263_;
  assign new_n53265_ = ~new_n53261_ & new_n53264_;
  assign new_n53266_ = ~new_n53223_ & ~new_n53265_;
  assign new_n53267_ = \b[5]  & ~new_n53212_;
  assign new_n53268_ = ~new_n53210_ & new_n53267_;
  assign new_n53269_ = ~new_n53214_ & ~new_n53268_;
  assign new_n53270_ = ~new_n53266_ & new_n53269_;
  assign new_n53271_ = ~new_n53214_ & ~new_n53270_;
  assign new_n53272_ = \b[6]  & ~new_n53203_;
  assign new_n53273_ = ~new_n53201_ & new_n53272_;
  assign new_n53274_ = ~new_n53205_ & ~new_n53273_;
  assign new_n53275_ = ~new_n53271_ & new_n53274_;
  assign new_n53276_ = ~new_n53205_ & ~new_n53275_;
  assign new_n53277_ = \b[7]  & ~new_n53194_;
  assign new_n53278_ = ~new_n53192_ & new_n53277_;
  assign new_n53279_ = ~new_n53196_ & ~new_n53278_;
  assign new_n53280_ = ~new_n53276_ & new_n53279_;
  assign new_n53281_ = ~new_n53196_ & ~new_n53280_;
  assign new_n53282_ = \b[8]  & ~new_n53185_;
  assign new_n53283_ = ~new_n53183_ & new_n53282_;
  assign new_n53284_ = ~new_n53187_ & ~new_n53283_;
  assign new_n53285_ = ~new_n53281_ & new_n53284_;
  assign new_n53286_ = ~new_n53187_ & ~new_n53285_;
  assign new_n53287_ = \b[9]  & ~new_n53176_;
  assign new_n53288_ = ~new_n53174_ & new_n53287_;
  assign new_n53289_ = ~new_n53178_ & ~new_n53288_;
  assign new_n53290_ = ~new_n53286_ & new_n53289_;
  assign new_n53291_ = ~new_n53178_ & ~new_n53290_;
  assign new_n53292_ = \b[10]  & ~new_n53167_;
  assign new_n53293_ = ~new_n53165_ & new_n53292_;
  assign new_n53294_ = ~new_n53169_ & ~new_n53293_;
  assign new_n53295_ = ~new_n53291_ & new_n53294_;
  assign new_n53296_ = ~new_n53169_ & ~new_n53295_;
  assign new_n53297_ = \b[11]  & ~new_n53158_;
  assign new_n53298_ = ~new_n53156_ & new_n53297_;
  assign new_n53299_ = ~new_n53160_ & ~new_n53298_;
  assign new_n53300_ = ~new_n53296_ & new_n53299_;
  assign new_n53301_ = ~new_n53160_ & ~new_n53300_;
  assign new_n53302_ = \b[12]  & ~new_n53149_;
  assign new_n53303_ = ~new_n53147_ & new_n53302_;
  assign new_n53304_ = ~new_n53151_ & ~new_n53303_;
  assign new_n53305_ = ~new_n53301_ & new_n53304_;
  assign new_n53306_ = ~new_n53151_ & ~new_n53305_;
  assign new_n53307_ = \b[13]  & ~new_n53140_;
  assign new_n53308_ = ~new_n53138_ & new_n53307_;
  assign new_n53309_ = ~new_n53142_ & ~new_n53308_;
  assign new_n53310_ = ~new_n53306_ & new_n53309_;
  assign new_n53311_ = ~new_n53142_ & ~new_n53310_;
  assign new_n53312_ = \b[14]  & ~new_n53131_;
  assign new_n53313_ = ~new_n53129_ & new_n53312_;
  assign new_n53314_ = ~new_n53133_ & ~new_n53313_;
  assign new_n53315_ = ~new_n53311_ & new_n53314_;
  assign new_n53316_ = ~new_n53133_ & ~new_n53315_;
  assign new_n53317_ = \b[15]  & ~new_n53122_;
  assign new_n53318_ = ~new_n53120_ & new_n53317_;
  assign new_n53319_ = ~new_n53124_ & ~new_n53318_;
  assign new_n53320_ = ~new_n53316_ & new_n53319_;
  assign new_n53321_ = ~new_n53124_ & ~new_n53320_;
  assign new_n53322_ = \b[16]  & ~new_n53113_;
  assign new_n53323_ = ~new_n53111_ & new_n53322_;
  assign new_n53324_ = ~new_n53115_ & ~new_n53323_;
  assign new_n53325_ = ~new_n53321_ & new_n53324_;
  assign new_n53326_ = ~new_n53115_ & ~new_n53325_;
  assign new_n53327_ = \b[17]  & ~new_n53104_;
  assign new_n53328_ = ~new_n53102_ & new_n53327_;
  assign new_n53329_ = ~new_n53106_ & ~new_n53328_;
  assign new_n53330_ = ~new_n53326_ & new_n53329_;
  assign new_n53331_ = ~new_n53106_ & ~new_n53330_;
  assign new_n53332_ = \b[18]  & ~new_n53095_;
  assign new_n53333_ = ~new_n53093_ & new_n53332_;
  assign new_n53334_ = ~new_n53097_ & ~new_n53333_;
  assign new_n53335_ = ~new_n53331_ & new_n53334_;
  assign new_n53336_ = ~new_n53097_ & ~new_n53335_;
  assign new_n53337_ = \b[19]  & ~new_n53086_;
  assign new_n53338_ = ~new_n53084_ & new_n53337_;
  assign new_n53339_ = ~new_n53088_ & ~new_n53338_;
  assign new_n53340_ = ~new_n53336_ & new_n53339_;
  assign new_n53341_ = ~new_n53088_ & ~new_n53340_;
  assign new_n53342_ = \b[20]  & ~new_n53077_;
  assign new_n53343_ = ~new_n53075_ & new_n53342_;
  assign new_n53344_ = ~new_n53079_ & ~new_n53343_;
  assign new_n53345_ = ~new_n53341_ & new_n53344_;
  assign new_n53346_ = ~new_n53079_ & ~new_n53345_;
  assign new_n53347_ = \b[21]  & ~new_n53068_;
  assign new_n53348_ = ~new_n53066_ & new_n53347_;
  assign new_n53349_ = ~new_n53070_ & ~new_n53348_;
  assign new_n53350_ = ~new_n53346_ & new_n53349_;
  assign new_n53351_ = ~new_n53070_ & ~new_n53350_;
  assign new_n53352_ = \b[22]  & ~new_n53059_;
  assign new_n53353_ = ~new_n53057_ & new_n53352_;
  assign new_n53354_ = ~new_n53061_ & ~new_n53353_;
  assign new_n53355_ = ~new_n53351_ & new_n53354_;
  assign new_n53356_ = ~new_n53061_ & ~new_n53355_;
  assign new_n53357_ = \b[23]  & ~new_n53050_;
  assign new_n53358_ = ~new_n53048_ & new_n53357_;
  assign new_n53359_ = ~new_n53052_ & ~new_n53358_;
  assign new_n53360_ = ~new_n53356_ & new_n53359_;
  assign new_n53361_ = ~new_n53052_ & ~new_n53360_;
  assign new_n53362_ = \b[24]  & ~new_n53041_;
  assign new_n53363_ = ~new_n53039_ & new_n53362_;
  assign new_n53364_ = ~new_n53043_ & ~new_n53363_;
  assign new_n53365_ = ~new_n53361_ & new_n53364_;
  assign new_n53366_ = ~new_n53043_ & ~new_n53365_;
  assign new_n53367_ = \b[25]  & ~new_n53032_;
  assign new_n53368_ = ~new_n53030_ & new_n53367_;
  assign new_n53369_ = ~new_n53034_ & ~new_n53368_;
  assign new_n53370_ = ~new_n53366_ & new_n53369_;
  assign new_n53371_ = ~new_n53034_ & ~new_n53370_;
  assign new_n53372_ = \b[26]  & ~new_n53023_;
  assign new_n53373_ = ~new_n53021_ & new_n53372_;
  assign new_n53374_ = ~new_n53025_ & ~new_n53373_;
  assign new_n53375_ = ~new_n53371_ & new_n53374_;
  assign new_n53376_ = ~new_n53025_ & ~new_n53375_;
  assign new_n53377_ = \b[27]  & ~new_n53014_;
  assign new_n53378_ = ~new_n53012_ & new_n53377_;
  assign new_n53379_ = ~new_n53016_ & ~new_n53378_;
  assign new_n53380_ = ~new_n53376_ & new_n53379_;
  assign new_n53381_ = ~new_n53016_ & ~new_n53380_;
  assign new_n53382_ = \b[28]  & ~new_n53005_;
  assign new_n53383_ = ~new_n53003_ & new_n53382_;
  assign new_n53384_ = ~new_n53007_ & ~new_n53383_;
  assign new_n53385_ = ~new_n53381_ & new_n53384_;
  assign new_n53386_ = ~new_n53007_ & ~new_n53385_;
  assign new_n53387_ = \b[29]  & ~new_n52996_;
  assign new_n53388_ = ~new_n52994_ & new_n53387_;
  assign new_n53389_ = ~new_n52998_ & ~new_n53388_;
  assign new_n53390_ = ~new_n53386_ & new_n53389_;
  assign new_n53391_ = ~new_n52998_ & ~new_n53390_;
  assign new_n53392_ = \b[30]  & ~new_n52987_;
  assign new_n53393_ = ~new_n52985_ & new_n53392_;
  assign new_n53394_ = ~new_n52989_ & ~new_n53393_;
  assign new_n53395_ = ~new_n53391_ & new_n53394_;
  assign new_n53396_ = ~new_n52989_ & ~new_n53395_;
  assign new_n53397_ = \b[31]  & ~new_n52978_;
  assign new_n53398_ = ~new_n52976_ & new_n53397_;
  assign new_n53399_ = ~new_n52980_ & ~new_n53398_;
  assign new_n53400_ = ~new_n53396_ & new_n53399_;
  assign new_n53401_ = ~new_n52980_ & ~new_n53400_;
  assign new_n53402_ = \b[32]  & ~new_n52969_;
  assign new_n53403_ = ~new_n52967_ & new_n53402_;
  assign new_n53404_ = ~new_n52971_ & ~new_n53403_;
  assign new_n53405_ = ~new_n53401_ & new_n53404_;
  assign new_n53406_ = ~new_n52971_ & ~new_n53405_;
  assign new_n53407_ = \b[33]  & ~new_n52960_;
  assign new_n53408_ = ~new_n52958_ & new_n53407_;
  assign new_n53409_ = ~new_n52962_ & ~new_n53408_;
  assign new_n53410_ = ~new_n53406_ & new_n53409_;
  assign new_n53411_ = ~new_n52962_ & ~new_n53410_;
  assign new_n53412_ = \b[34]  & ~new_n52951_;
  assign new_n53413_ = ~new_n52949_ & new_n53412_;
  assign new_n53414_ = ~new_n52953_ & ~new_n53413_;
  assign new_n53415_ = ~new_n53411_ & new_n53414_;
  assign new_n53416_ = ~new_n52953_ & ~new_n53415_;
  assign new_n53417_ = \b[35]  & ~new_n52942_;
  assign new_n53418_ = ~new_n52940_ & new_n53417_;
  assign new_n53419_ = ~new_n52944_ & ~new_n53418_;
  assign new_n53420_ = ~new_n53416_ & new_n53419_;
  assign new_n53421_ = ~new_n52944_ & ~new_n53420_;
  assign new_n53422_ = \b[36]  & ~new_n52933_;
  assign new_n53423_ = ~new_n52931_ & new_n53422_;
  assign new_n53424_ = ~new_n52935_ & ~new_n53423_;
  assign new_n53425_ = ~new_n53421_ & new_n53424_;
  assign new_n53426_ = ~new_n52935_ & ~new_n53425_;
  assign new_n53427_ = \b[37]  & ~new_n52924_;
  assign new_n53428_ = ~new_n52922_ & new_n53427_;
  assign new_n53429_ = ~new_n52926_ & ~new_n53428_;
  assign new_n53430_ = ~new_n53426_ & new_n53429_;
  assign new_n53431_ = ~new_n52926_ & ~new_n53430_;
  assign new_n53432_ = \b[38]  & ~new_n52915_;
  assign new_n53433_ = ~new_n52913_ & new_n53432_;
  assign new_n53434_ = ~new_n52917_ & ~new_n53433_;
  assign new_n53435_ = ~new_n53431_ & new_n53434_;
  assign new_n53436_ = ~new_n52917_ & ~new_n53435_;
  assign new_n53437_ = \b[39]  & ~new_n52906_;
  assign new_n53438_ = ~new_n52904_ & new_n53437_;
  assign new_n53439_ = ~new_n52908_ & ~new_n53438_;
  assign new_n53440_ = ~new_n53436_ & new_n53439_;
  assign new_n53441_ = ~new_n52908_ & ~new_n53440_;
  assign new_n53442_ = \b[40]  & ~new_n52897_;
  assign new_n53443_ = ~new_n52895_ & new_n53442_;
  assign new_n53444_ = ~new_n52899_ & ~new_n53443_;
  assign new_n53445_ = ~new_n53441_ & new_n53444_;
  assign new_n53446_ = ~new_n52899_ & ~new_n53445_;
  assign new_n53447_ = \b[41]  & ~new_n52888_;
  assign new_n53448_ = ~new_n52886_ & new_n53447_;
  assign new_n53449_ = ~new_n52890_ & ~new_n53448_;
  assign new_n53450_ = ~new_n53446_ & new_n53449_;
  assign new_n53451_ = ~new_n52890_ & ~new_n53450_;
  assign new_n53452_ = \b[42]  & ~new_n52879_;
  assign new_n53453_ = ~new_n52877_ & new_n53452_;
  assign new_n53454_ = ~new_n52881_ & ~new_n53453_;
  assign new_n53455_ = ~new_n53451_ & new_n53454_;
  assign new_n53456_ = ~new_n52881_ & ~new_n53455_;
  assign new_n53457_ = \b[43]  & ~new_n52870_;
  assign new_n53458_ = ~new_n52868_ & new_n53457_;
  assign new_n53459_ = ~new_n52872_ & ~new_n53458_;
  assign new_n53460_ = ~new_n53456_ & new_n53459_;
  assign new_n53461_ = ~new_n52872_ & ~new_n53460_;
  assign new_n53462_ = \b[44]  & ~new_n52861_;
  assign new_n53463_ = ~new_n52859_ & new_n53462_;
  assign new_n53464_ = ~new_n52863_ & ~new_n53463_;
  assign new_n53465_ = ~new_n53461_ & new_n53464_;
  assign new_n53466_ = ~new_n52863_ & ~new_n53465_;
  assign new_n53467_ = \b[45]  & ~new_n52852_;
  assign new_n53468_ = ~new_n52850_ & new_n53467_;
  assign new_n53469_ = ~new_n52854_ & ~new_n53468_;
  assign new_n53470_ = ~new_n53466_ & new_n53469_;
  assign new_n53471_ = ~new_n52854_ & ~new_n53470_;
  assign new_n53472_ = \b[46]  & ~new_n52843_;
  assign new_n53473_ = ~new_n52841_ & new_n53472_;
  assign new_n53474_ = ~new_n52845_ & ~new_n53473_;
  assign new_n53475_ = ~new_n53471_ & new_n53474_;
  assign new_n53476_ = ~new_n52845_ & ~new_n53475_;
  assign new_n53477_ = \b[47]  & ~new_n52834_;
  assign new_n53478_ = ~new_n52832_ & new_n53477_;
  assign new_n53479_ = ~new_n52836_ & ~new_n53478_;
  assign new_n53480_ = ~new_n53476_ & new_n53479_;
  assign new_n53481_ = ~new_n52836_ & ~new_n53480_;
  assign new_n53482_ = \b[48]  & ~new_n52825_;
  assign new_n53483_ = ~new_n52823_ & new_n53482_;
  assign new_n53484_ = ~new_n52827_ & ~new_n53483_;
  assign new_n53485_ = ~new_n53481_ & new_n53484_;
  assign new_n53486_ = ~new_n52827_ & ~new_n53485_;
  assign new_n53487_ = \b[49]  & ~new_n52816_;
  assign new_n53488_ = ~new_n52814_ & new_n53487_;
  assign new_n53489_ = ~new_n52818_ & ~new_n53488_;
  assign new_n53490_ = ~new_n53486_ & new_n53489_;
  assign new_n53491_ = ~new_n52818_ & ~new_n53490_;
  assign new_n53492_ = \b[50]  & ~new_n52807_;
  assign new_n53493_ = ~new_n52805_ & new_n53492_;
  assign new_n53494_ = ~new_n52809_ & ~new_n53493_;
  assign new_n53495_ = ~new_n53491_ & new_n53494_;
  assign new_n53496_ = ~new_n52809_ & ~new_n53495_;
  assign new_n53497_ = \b[51]  & ~new_n52798_;
  assign new_n53498_ = ~new_n52796_ & new_n53497_;
  assign new_n53499_ = ~new_n52800_ & ~new_n53498_;
  assign new_n53500_ = ~new_n53496_ & new_n53499_;
  assign new_n53501_ = ~new_n52800_ & ~new_n53500_;
  assign new_n53502_ = \b[52]  & ~new_n52789_;
  assign new_n53503_ = ~new_n52787_ & new_n53502_;
  assign new_n53504_ = ~new_n52791_ & ~new_n53503_;
  assign new_n53505_ = ~new_n53501_ & new_n53504_;
  assign new_n53506_ = ~new_n52791_ & ~new_n53505_;
  assign new_n53507_ = \b[53]  & ~new_n52780_;
  assign new_n53508_ = ~new_n52778_ & new_n53507_;
  assign new_n53509_ = ~new_n52782_ & ~new_n53508_;
  assign new_n53510_ = ~new_n53506_ & new_n53509_;
  assign new_n53511_ = ~new_n52782_ & ~new_n53510_;
  assign new_n53512_ = \b[54]  & ~new_n52771_;
  assign new_n53513_ = ~new_n52769_ & new_n53512_;
  assign new_n53514_ = ~new_n52773_ & ~new_n53513_;
  assign new_n53515_ = ~new_n53511_ & new_n53514_;
  assign new_n53516_ = ~new_n52773_ & ~new_n53515_;
  assign new_n53517_ = \b[55]  & ~new_n52762_;
  assign new_n53518_ = ~new_n52760_ & new_n53517_;
  assign new_n53519_ = ~new_n52764_ & ~new_n53518_;
  assign new_n53520_ = ~new_n53516_ & new_n53519_;
  assign new_n53521_ = ~new_n52764_ & ~new_n53520_;
  assign new_n53522_ = \b[56]  & ~new_n52753_;
  assign new_n53523_ = ~new_n52751_ & new_n53522_;
  assign new_n53524_ = ~new_n52755_ & ~new_n53523_;
  assign new_n53525_ = ~new_n53521_ & new_n53524_;
  assign new_n53526_ = ~new_n52755_ & ~new_n53525_;
  assign new_n53527_ = \b[57]  & ~new_n52744_;
  assign new_n53528_ = ~new_n52742_ & new_n53527_;
  assign new_n53529_ = ~new_n52746_ & ~new_n53528_;
  assign new_n53530_ = ~new_n53526_ & new_n53529_;
  assign new_n53531_ = ~new_n52746_ & ~new_n53530_;
  assign new_n53532_ = \b[58]  & ~new_n52735_;
  assign new_n53533_ = ~new_n52733_ & new_n53532_;
  assign new_n53534_ = ~new_n52737_ & ~new_n53533_;
  assign new_n53535_ = ~new_n53531_ & new_n53534_;
  assign new_n53536_ = ~new_n52737_ & ~new_n53535_;
  assign new_n53537_ = ~new_n51928_ & ~new_n52723_;
  assign new_n53538_ = ~new_n52721_ & new_n53537_;
  assign new_n53539_ = ~new_n52712_ & new_n53538_;
  assign new_n53540_ = ~new_n52721_ & ~new_n52723_;
  assign new_n53541_ = ~new_n52713_ & ~new_n53540_;
  assign new_n53542_ = ~new_n53539_ & ~new_n53541_;
  assign new_n53543_ = ~new_n52728_ & ~new_n53542_;
  assign new_n53544_ = ~new_n52720_ & ~new_n52727_;
  assign new_n53545_ = ~new_n52726_ & new_n53544_;
  assign new_n53546_ = ~new_n53543_ & ~new_n53545_;
  assign new_n53547_ = ~\b[59]  & ~new_n53546_;
  assign new_n53548_ = \b[59]  & ~new_n53545_;
  assign new_n53549_ = ~new_n53543_ & new_n53548_;
  assign new_n53550_ = new_n280_ & ~new_n53549_;
  assign new_n53551_ = ~new_n53547_ & new_n53550_;
  assign new_n53552_ = ~new_n53536_ & new_n53551_;
  assign new_n53553_ = new_n24707_ & ~new_n53546_;
  assign new_n53554_ = ~new_n53552_ & ~new_n53553_;
  assign new_n53555_ = ~new_n52746_ & new_n53534_;
  assign new_n53556_ = ~new_n53530_ & new_n53555_;
  assign new_n53557_ = ~new_n53531_ & ~new_n53534_;
  assign new_n53558_ = ~new_n53556_ & ~new_n53557_;
  assign new_n53559_ = ~new_n53554_ & ~new_n53558_;
  assign new_n53560_ = ~new_n52736_ & ~new_n53553_;
  assign new_n53561_ = ~new_n53552_ & new_n53560_;
  assign new_n53562_ = ~new_n53559_ & ~new_n53561_;
  assign new_n53563_ = ~\b[59]  & ~new_n53562_;
  assign new_n53564_ = ~new_n52755_ & new_n53529_;
  assign new_n53565_ = ~new_n53525_ & new_n53564_;
  assign new_n53566_ = ~new_n53526_ & ~new_n53529_;
  assign new_n53567_ = ~new_n53565_ & ~new_n53566_;
  assign new_n53568_ = ~new_n53554_ & ~new_n53567_;
  assign new_n53569_ = ~new_n52745_ & ~new_n53553_;
  assign new_n53570_ = ~new_n53552_ & new_n53569_;
  assign new_n53571_ = ~new_n53568_ & ~new_n53570_;
  assign new_n53572_ = ~\b[58]  & ~new_n53571_;
  assign new_n53573_ = ~new_n52764_ & new_n53524_;
  assign new_n53574_ = ~new_n53520_ & new_n53573_;
  assign new_n53575_ = ~new_n53521_ & ~new_n53524_;
  assign new_n53576_ = ~new_n53574_ & ~new_n53575_;
  assign new_n53577_ = ~new_n53554_ & ~new_n53576_;
  assign new_n53578_ = ~new_n52754_ & ~new_n53553_;
  assign new_n53579_ = ~new_n53552_ & new_n53578_;
  assign new_n53580_ = ~new_n53577_ & ~new_n53579_;
  assign new_n53581_ = ~\b[57]  & ~new_n53580_;
  assign new_n53582_ = ~new_n52773_ & new_n53519_;
  assign new_n53583_ = ~new_n53515_ & new_n53582_;
  assign new_n53584_ = ~new_n53516_ & ~new_n53519_;
  assign new_n53585_ = ~new_n53583_ & ~new_n53584_;
  assign new_n53586_ = ~new_n53554_ & ~new_n53585_;
  assign new_n53587_ = ~new_n52763_ & ~new_n53553_;
  assign new_n53588_ = ~new_n53552_ & new_n53587_;
  assign new_n53589_ = ~new_n53586_ & ~new_n53588_;
  assign new_n53590_ = ~\b[56]  & ~new_n53589_;
  assign new_n53591_ = ~new_n52782_ & new_n53514_;
  assign new_n53592_ = ~new_n53510_ & new_n53591_;
  assign new_n53593_ = ~new_n53511_ & ~new_n53514_;
  assign new_n53594_ = ~new_n53592_ & ~new_n53593_;
  assign new_n53595_ = ~new_n53554_ & ~new_n53594_;
  assign new_n53596_ = ~new_n52772_ & ~new_n53553_;
  assign new_n53597_ = ~new_n53552_ & new_n53596_;
  assign new_n53598_ = ~new_n53595_ & ~new_n53597_;
  assign new_n53599_ = ~\b[55]  & ~new_n53598_;
  assign new_n53600_ = ~new_n52791_ & new_n53509_;
  assign new_n53601_ = ~new_n53505_ & new_n53600_;
  assign new_n53602_ = ~new_n53506_ & ~new_n53509_;
  assign new_n53603_ = ~new_n53601_ & ~new_n53602_;
  assign new_n53604_ = ~new_n53554_ & ~new_n53603_;
  assign new_n53605_ = ~new_n52781_ & ~new_n53553_;
  assign new_n53606_ = ~new_n53552_ & new_n53605_;
  assign new_n53607_ = ~new_n53604_ & ~new_n53606_;
  assign new_n53608_ = ~\b[54]  & ~new_n53607_;
  assign new_n53609_ = ~new_n52800_ & new_n53504_;
  assign new_n53610_ = ~new_n53500_ & new_n53609_;
  assign new_n53611_ = ~new_n53501_ & ~new_n53504_;
  assign new_n53612_ = ~new_n53610_ & ~new_n53611_;
  assign new_n53613_ = ~new_n53554_ & ~new_n53612_;
  assign new_n53614_ = ~new_n52790_ & ~new_n53553_;
  assign new_n53615_ = ~new_n53552_ & new_n53614_;
  assign new_n53616_ = ~new_n53613_ & ~new_n53615_;
  assign new_n53617_ = ~\b[53]  & ~new_n53616_;
  assign new_n53618_ = ~new_n52809_ & new_n53499_;
  assign new_n53619_ = ~new_n53495_ & new_n53618_;
  assign new_n53620_ = ~new_n53496_ & ~new_n53499_;
  assign new_n53621_ = ~new_n53619_ & ~new_n53620_;
  assign new_n53622_ = ~new_n53554_ & ~new_n53621_;
  assign new_n53623_ = ~new_n52799_ & ~new_n53553_;
  assign new_n53624_ = ~new_n53552_ & new_n53623_;
  assign new_n53625_ = ~new_n53622_ & ~new_n53624_;
  assign new_n53626_ = ~\b[52]  & ~new_n53625_;
  assign new_n53627_ = ~new_n52818_ & new_n53494_;
  assign new_n53628_ = ~new_n53490_ & new_n53627_;
  assign new_n53629_ = ~new_n53491_ & ~new_n53494_;
  assign new_n53630_ = ~new_n53628_ & ~new_n53629_;
  assign new_n53631_ = ~new_n53554_ & ~new_n53630_;
  assign new_n53632_ = ~new_n52808_ & ~new_n53553_;
  assign new_n53633_ = ~new_n53552_ & new_n53632_;
  assign new_n53634_ = ~new_n53631_ & ~new_n53633_;
  assign new_n53635_ = ~\b[51]  & ~new_n53634_;
  assign new_n53636_ = ~new_n52827_ & new_n53489_;
  assign new_n53637_ = ~new_n53485_ & new_n53636_;
  assign new_n53638_ = ~new_n53486_ & ~new_n53489_;
  assign new_n53639_ = ~new_n53637_ & ~new_n53638_;
  assign new_n53640_ = ~new_n53554_ & ~new_n53639_;
  assign new_n53641_ = ~new_n52817_ & ~new_n53553_;
  assign new_n53642_ = ~new_n53552_ & new_n53641_;
  assign new_n53643_ = ~new_n53640_ & ~new_n53642_;
  assign new_n53644_ = ~\b[50]  & ~new_n53643_;
  assign new_n53645_ = ~new_n52836_ & new_n53484_;
  assign new_n53646_ = ~new_n53480_ & new_n53645_;
  assign new_n53647_ = ~new_n53481_ & ~new_n53484_;
  assign new_n53648_ = ~new_n53646_ & ~new_n53647_;
  assign new_n53649_ = ~new_n53554_ & ~new_n53648_;
  assign new_n53650_ = ~new_n52826_ & ~new_n53553_;
  assign new_n53651_ = ~new_n53552_ & new_n53650_;
  assign new_n53652_ = ~new_n53649_ & ~new_n53651_;
  assign new_n53653_ = ~\b[49]  & ~new_n53652_;
  assign new_n53654_ = ~new_n52845_ & new_n53479_;
  assign new_n53655_ = ~new_n53475_ & new_n53654_;
  assign new_n53656_ = ~new_n53476_ & ~new_n53479_;
  assign new_n53657_ = ~new_n53655_ & ~new_n53656_;
  assign new_n53658_ = ~new_n53554_ & ~new_n53657_;
  assign new_n53659_ = ~new_n52835_ & ~new_n53553_;
  assign new_n53660_ = ~new_n53552_ & new_n53659_;
  assign new_n53661_ = ~new_n53658_ & ~new_n53660_;
  assign new_n53662_ = ~\b[48]  & ~new_n53661_;
  assign new_n53663_ = ~new_n52854_ & new_n53474_;
  assign new_n53664_ = ~new_n53470_ & new_n53663_;
  assign new_n53665_ = ~new_n53471_ & ~new_n53474_;
  assign new_n53666_ = ~new_n53664_ & ~new_n53665_;
  assign new_n53667_ = ~new_n53554_ & ~new_n53666_;
  assign new_n53668_ = ~new_n52844_ & ~new_n53553_;
  assign new_n53669_ = ~new_n53552_ & new_n53668_;
  assign new_n53670_ = ~new_n53667_ & ~new_n53669_;
  assign new_n53671_ = ~\b[47]  & ~new_n53670_;
  assign new_n53672_ = ~new_n52863_ & new_n53469_;
  assign new_n53673_ = ~new_n53465_ & new_n53672_;
  assign new_n53674_ = ~new_n53466_ & ~new_n53469_;
  assign new_n53675_ = ~new_n53673_ & ~new_n53674_;
  assign new_n53676_ = ~new_n53554_ & ~new_n53675_;
  assign new_n53677_ = ~new_n52853_ & ~new_n53553_;
  assign new_n53678_ = ~new_n53552_ & new_n53677_;
  assign new_n53679_ = ~new_n53676_ & ~new_n53678_;
  assign new_n53680_ = ~\b[46]  & ~new_n53679_;
  assign new_n53681_ = ~new_n52872_ & new_n53464_;
  assign new_n53682_ = ~new_n53460_ & new_n53681_;
  assign new_n53683_ = ~new_n53461_ & ~new_n53464_;
  assign new_n53684_ = ~new_n53682_ & ~new_n53683_;
  assign new_n53685_ = ~new_n53554_ & ~new_n53684_;
  assign new_n53686_ = ~new_n52862_ & ~new_n53553_;
  assign new_n53687_ = ~new_n53552_ & new_n53686_;
  assign new_n53688_ = ~new_n53685_ & ~new_n53687_;
  assign new_n53689_ = ~\b[45]  & ~new_n53688_;
  assign new_n53690_ = ~new_n52881_ & new_n53459_;
  assign new_n53691_ = ~new_n53455_ & new_n53690_;
  assign new_n53692_ = ~new_n53456_ & ~new_n53459_;
  assign new_n53693_ = ~new_n53691_ & ~new_n53692_;
  assign new_n53694_ = ~new_n53554_ & ~new_n53693_;
  assign new_n53695_ = ~new_n52871_ & ~new_n53553_;
  assign new_n53696_ = ~new_n53552_ & new_n53695_;
  assign new_n53697_ = ~new_n53694_ & ~new_n53696_;
  assign new_n53698_ = ~\b[44]  & ~new_n53697_;
  assign new_n53699_ = ~new_n52890_ & new_n53454_;
  assign new_n53700_ = ~new_n53450_ & new_n53699_;
  assign new_n53701_ = ~new_n53451_ & ~new_n53454_;
  assign new_n53702_ = ~new_n53700_ & ~new_n53701_;
  assign new_n53703_ = ~new_n53554_ & ~new_n53702_;
  assign new_n53704_ = ~new_n52880_ & ~new_n53553_;
  assign new_n53705_ = ~new_n53552_ & new_n53704_;
  assign new_n53706_ = ~new_n53703_ & ~new_n53705_;
  assign new_n53707_ = ~\b[43]  & ~new_n53706_;
  assign new_n53708_ = ~new_n52899_ & new_n53449_;
  assign new_n53709_ = ~new_n53445_ & new_n53708_;
  assign new_n53710_ = ~new_n53446_ & ~new_n53449_;
  assign new_n53711_ = ~new_n53709_ & ~new_n53710_;
  assign new_n53712_ = ~new_n53554_ & ~new_n53711_;
  assign new_n53713_ = ~new_n52889_ & ~new_n53553_;
  assign new_n53714_ = ~new_n53552_ & new_n53713_;
  assign new_n53715_ = ~new_n53712_ & ~new_n53714_;
  assign new_n53716_ = ~\b[42]  & ~new_n53715_;
  assign new_n53717_ = ~new_n52908_ & new_n53444_;
  assign new_n53718_ = ~new_n53440_ & new_n53717_;
  assign new_n53719_ = ~new_n53441_ & ~new_n53444_;
  assign new_n53720_ = ~new_n53718_ & ~new_n53719_;
  assign new_n53721_ = ~new_n53554_ & ~new_n53720_;
  assign new_n53722_ = ~new_n52898_ & ~new_n53553_;
  assign new_n53723_ = ~new_n53552_ & new_n53722_;
  assign new_n53724_ = ~new_n53721_ & ~new_n53723_;
  assign new_n53725_ = ~\b[41]  & ~new_n53724_;
  assign new_n53726_ = ~new_n52917_ & new_n53439_;
  assign new_n53727_ = ~new_n53435_ & new_n53726_;
  assign new_n53728_ = ~new_n53436_ & ~new_n53439_;
  assign new_n53729_ = ~new_n53727_ & ~new_n53728_;
  assign new_n53730_ = ~new_n53554_ & ~new_n53729_;
  assign new_n53731_ = ~new_n52907_ & ~new_n53553_;
  assign new_n53732_ = ~new_n53552_ & new_n53731_;
  assign new_n53733_ = ~new_n53730_ & ~new_n53732_;
  assign new_n53734_ = ~\b[40]  & ~new_n53733_;
  assign new_n53735_ = ~new_n52926_ & new_n53434_;
  assign new_n53736_ = ~new_n53430_ & new_n53735_;
  assign new_n53737_ = ~new_n53431_ & ~new_n53434_;
  assign new_n53738_ = ~new_n53736_ & ~new_n53737_;
  assign new_n53739_ = ~new_n53554_ & ~new_n53738_;
  assign new_n53740_ = ~new_n52916_ & ~new_n53553_;
  assign new_n53741_ = ~new_n53552_ & new_n53740_;
  assign new_n53742_ = ~new_n53739_ & ~new_n53741_;
  assign new_n53743_ = ~\b[39]  & ~new_n53742_;
  assign new_n53744_ = ~new_n52935_ & new_n53429_;
  assign new_n53745_ = ~new_n53425_ & new_n53744_;
  assign new_n53746_ = ~new_n53426_ & ~new_n53429_;
  assign new_n53747_ = ~new_n53745_ & ~new_n53746_;
  assign new_n53748_ = ~new_n53554_ & ~new_n53747_;
  assign new_n53749_ = ~new_n52925_ & ~new_n53553_;
  assign new_n53750_ = ~new_n53552_ & new_n53749_;
  assign new_n53751_ = ~new_n53748_ & ~new_n53750_;
  assign new_n53752_ = ~\b[38]  & ~new_n53751_;
  assign new_n53753_ = ~new_n52944_ & new_n53424_;
  assign new_n53754_ = ~new_n53420_ & new_n53753_;
  assign new_n53755_ = ~new_n53421_ & ~new_n53424_;
  assign new_n53756_ = ~new_n53754_ & ~new_n53755_;
  assign new_n53757_ = ~new_n53554_ & ~new_n53756_;
  assign new_n53758_ = ~new_n52934_ & ~new_n53553_;
  assign new_n53759_ = ~new_n53552_ & new_n53758_;
  assign new_n53760_ = ~new_n53757_ & ~new_n53759_;
  assign new_n53761_ = ~\b[37]  & ~new_n53760_;
  assign new_n53762_ = ~new_n52953_ & new_n53419_;
  assign new_n53763_ = ~new_n53415_ & new_n53762_;
  assign new_n53764_ = ~new_n53416_ & ~new_n53419_;
  assign new_n53765_ = ~new_n53763_ & ~new_n53764_;
  assign new_n53766_ = ~new_n53554_ & ~new_n53765_;
  assign new_n53767_ = ~new_n52943_ & ~new_n53553_;
  assign new_n53768_ = ~new_n53552_ & new_n53767_;
  assign new_n53769_ = ~new_n53766_ & ~new_n53768_;
  assign new_n53770_ = ~\b[36]  & ~new_n53769_;
  assign new_n53771_ = ~new_n52962_ & new_n53414_;
  assign new_n53772_ = ~new_n53410_ & new_n53771_;
  assign new_n53773_ = ~new_n53411_ & ~new_n53414_;
  assign new_n53774_ = ~new_n53772_ & ~new_n53773_;
  assign new_n53775_ = ~new_n53554_ & ~new_n53774_;
  assign new_n53776_ = ~new_n52952_ & ~new_n53553_;
  assign new_n53777_ = ~new_n53552_ & new_n53776_;
  assign new_n53778_ = ~new_n53775_ & ~new_n53777_;
  assign new_n53779_ = ~\b[35]  & ~new_n53778_;
  assign new_n53780_ = ~new_n52971_ & new_n53409_;
  assign new_n53781_ = ~new_n53405_ & new_n53780_;
  assign new_n53782_ = ~new_n53406_ & ~new_n53409_;
  assign new_n53783_ = ~new_n53781_ & ~new_n53782_;
  assign new_n53784_ = ~new_n53554_ & ~new_n53783_;
  assign new_n53785_ = ~new_n52961_ & ~new_n53553_;
  assign new_n53786_ = ~new_n53552_ & new_n53785_;
  assign new_n53787_ = ~new_n53784_ & ~new_n53786_;
  assign new_n53788_ = ~\b[34]  & ~new_n53787_;
  assign new_n53789_ = ~new_n52980_ & new_n53404_;
  assign new_n53790_ = ~new_n53400_ & new_n53789_;
  assign new_n53791_ = ~new_n53401_ & ~new_n53404_;
  assign new_n53792_ = ~new_n53790_ & ~new_n53791_;
  assign new_n53793_ = ~new_n53554_ & ~new_n53792_;
  assign new_n53794_ = ~new_n52970_ & ~new_n53553_;
  assign new_n53795_ = ~new_n53552_ & new_n53794_;
  assign new_n53796_ = ~new_n53793_ & ~new_n53795_;
  assign new_n53797_ = ~\b[33]  & ~new_n53796_;
  assign new_n53798_ = ~new_n52989_ & new_n53399_;
  assign new_n53799_ = ~new_n53395_ & new_n53798_;
  assign new_n53800_ = ~new_n53396_ & ~new_n53399_;
  assign new_n53801_ = ~new_n53799_ & ~new_n53800_;
  assign new_n53802_ = ~new_n53554_ & ~new_n53801_;
  assign new_n53803_ = ~new_n52979_ & ~new_n53553_;
  assign new_n53804_ = ~new_n53552_ & new_n53803_;
  assign new_n53805_ = ~new_n53802_ & ~new_n53804_;
  assign new_n53806_ = ~\b[32]  & ~new_n53805_;
  assign new_n53807_ = ~new_n52998_ & new_n53394_;
  assign new_n53808_ = ~new_n53390_ & new_n53807_;
  assign new_n53809_ = ~new_n53391_ & ~new_n53394_;
  assign new_n53810_ = ~new_n53808_ & ~new_n53809_;
  assign new_n53811_ = ~new_n53554_ & ~new_n53810_;
  assign new_n53812_ = ~new_n52988_ & ~new_n53553_;
  assign new_n53813_ = ~new_n53552_ & new_n53812_;
  assign new_n53814_ = ~new_n53811_ & ~new_n53813_;
  assign new_n53815_ = ~\b[31]  & ~new_n53814_;
  assign new_n53816_ = ~new_n53007_ & new_n53389_;
  assign new_n53817_ = ~new_n53385_ & new_n53816_;
  assign new_n53818_ = ~new_n53386_ & ~new_n53389_;
  assign new_n53819_ = ~new_n53817_ & ~new_n53818_;
  assign new_n53820_ = ~new_n53554_ & ~new_n53819_;
  assign new_n53821_ = ~new_n52997_ & ~new_n53553_;
  assign new_n53822_ = ~new_n53552_ & new_n53821_;
  assign new_n53823_ = ~new_n53820_ & ~new_n53822_;
  assign new_n53824_ = ~\b[30]  & ~new_n53823_;
  assign new_n53825_ = ~new_n53016_ & new_n53384_;
  assign new_n53826_ = ~new_n53380_ & new_n53825_;
  assign new_n53827_ = ~new_n53381_ & ~new_n53384_;
  assign new_n53828_ = ~new_n53826_ & ~new_n53827_;
  assign new_n53829_ = ~new_n53554_ & ~new_n53828_;
  assign new_n53830_ = ~new_n53006_ & ~new_n53553_;
  assign new_n53831_ = ~new_n53552_ & new_n53830_;
  assign new_n53832_ = ~new_n53829_ & ~new_n53831_;
  assign new_n53833_ = ~\b[29]  & ~new_n53832_;
  assign new_n53834_ = ~new_n53025_ & new_n53379_;
  assign new_n53835_ = ~new_n53375_ & new_n53834_;
  assign new_n53836_ = ~new_n53376_ & ~new_n53379_;
  assign new_n53837_ = ~new_n53835_ & ~new_n53836_;
  assign new_n53838_ = ~new_n53554_ & ~new_n53837_;
  assign new_n53839_ = ~new_n53015_ & ~new_n53553_;
  assign new_n53840_ = ~new_n53552_ & new_n53839_;
  assign new_n53841_ = ~new_n53838_ & ~new_n53840_;
  assign new_n53842_ = ~\b[28]  & ~new_n53841_;
  assign new_n53843_ = ~new_n53034_ & new_n53374_;
  assign new_n53844_ = ~new_n53370_ & new_n53843_;
  assign new_n53845_ = ~new_n53371_ & ~new_n53374_;
  assign new_n53846_ = ~new_n53844_ & ~new_n53845_;
  assign new_n53847_ = ~new_n53554_ & ~new_n53846_;
  assign new_n53848_ = ~new_n53024_ & ~new_n53553_;
  assign new_n53849_ = ~new_n53552_ & new_n53848_;
  assign new_n53850_ = ~new_n53847_ & ~new_n53849_;
  assign new_n53851_ = ~\b[27]  & ~new_n53850_;
  assign new_n53852_ = ~new_n53043_ & new_n53369_;
  assign new_n53853_ = ~new_n53365_ & new_n53852_;
  assign new_n53854_ = ~new_n53366_ & ~new_n53369_;
  assign new_n53855_ = ~new_n53853_ & ~new_n53854_;
  assign new_n53856_ = ~new_n53554_ & ~new_n53855_;
  assign new_n53857_ = ~new_n53033_ & ~new_n53553_;
  assign new_n53858_ = ~new_n53552_ & new_n53857_;
  assign new_n53859_ = ~new_n53856_ & ~new_n53858_;
  assign new_n53860_ = ~\b[26]  & ~new_n53859_;
  assign new_n53861_ = ~new_n53052_ & new_n53364_;
  assign new_n53862_ = ~new_n53360_ & new_n53861_;
  assign new_n53863_ = ~new_n53361_ & ~new_n53364_;
  assign new_n53864_ = ~new_n53862_ & ~new_n53863_;
  assign new_n53865_ = ~new_n53554_ & ~new_n53864_;
  assign new_n53866_ = ~new_n53042_ & ~new_n53553_;
  assign new_n53867_ = ~new_n53552_ & new_n53866_;
  assign new_n53868_ = ~new_n53865_ & ~new_n53867_;
  assign new_n53869_ = ~\b[25]  & ~new_n53868_;
  assign new_n53870_ = ~new_n53061_ & new_n53359_;
  assign new_n53871_ = ~new_n53355_ & new_n53870_;
  assign new_n53872_ = ~new_n53356_ & ~new_n53359_;
  assign new_n53873_ = ~new_n53871_ & ~new_n53872_;
  assign new_n53874_ = ~new_n53554_ & ~new_n53873_;
  assign new_n53875_ = ~new_n53051_ & ~new_n53553_;
  assign new_n53876_ = ~new_n53552_ & new_n53875_;
  assign new_n53877_ = ~new_n53874_ & ~new_n53876_;
  assign new_n53878_ = ~\b[24]  & ~new_n53877_;
  assign new_n53879_ = ~new_n53070_ & new_n53354_;
  assign new_n53880_ = ~new_n53350_ & new_n53879_;
  assign new_n53881_ = ~new_n53351_ & ~new_n53354_;
  assign new_n53882_ = ~new_n53880_ & ~new_n53881_;
  assign new_n53883_ = ~new_n53554_ & ~new_n53882_;
  assign new_n53884_ = ~new_n53060_ & ~new_n53553_;
  assign new_n53885_ = ~new_n53552_ & new_n53884_;
  assign new_n53886_ = ~new_n53883_ & ~new_n53885_;
  assign new_n53887_ = ~\b[23]  & ~new_n53886_;
  assign new_n53888_ = ~new_n53079_ & new_n53349_;
  assign new_n53889_ = ~new_n53345_ & new_n53888_;
  assign new_n53890_ = ~new_n53346_ & ~new_n53349_;
  assign new_n53891_ = ~new_n53889_ & ~new_n53890_;
  assign new_n53892_ = ~new_n53554_ & ~new_n53891_;
  assign new_n53893_ = ~new_n53069_ & ~new_n53553_;
  assign new_n53894_ = ~new_n53552_ & new_n53893_;
  assign new_n53895_ = ~new_n53892_ & ~new_n53894_;
  assign new_n53896_ = ~\b[22]  & ~new_n53895_;
  assign new_n53897_ = ~new_n53088_ & new_n53344_;
  assign new_n53898_ = ~new_n53340_ & new_n53897_;
  assign new_n53899_ = ~new_n53341_ & ~new_n53344_;
  assign new_n53900_ = ~new_n53898_ & ~new_n53899_;
  assign new_n53901_ = ~new_n53554_ & ~new_n53900_;
  assign new_n53902_ = ~new_n53078_ & ~new_n53553_;
  assign new_n53903_ = ~new_n53552_ & new_n53902_;
  assign new_n53904_ = ~new_n53901_ & ~new_n53903_;
  assign new_n53905_ = ~\b[21]  & ~new_n53904_;
  assign new_n53906_ = ~new_n53097_ & new_n53339_;
  assign new_n53907_ = ~new_n53335_ & new_n53906_;
  assign new_n53908_ = ~new_n53336_ & ~new_n53339_;
  assign new_n53909_ = ~new_n53907_ & ~new_n53908_;
  assign new_n53910_ = ~new_n53554_ & ~new_n53909_;
  assign new_n53911_ = ~new_n53087_ & ~new_n53553_;
  assign new_n53912_ = ~new_n53552_ & new_n53911_;
  assign new_n53913_ = ~new_n53910_ & ~new_n53912_;
  assign new_n53914_ = ~\b[20]  & ~new_n53913_;
  assign new_n53915_ = ~new_n53106_ & new_n53334_;
  assign new_n53916_ = ~new_n53330_ & new_n53915_;
  assign new_n53917_ = ~new_n53331_ & ~new_n53334_;
  assign new_n53918_ = ~new_n53916_ & ~new_n53917_;
  assign new_n53919_ = ~new_n53554_ & ~new_n53918_;
  assign new_n53920_ = ~new_n53096_ & ~new_n53553_;
  assign new_n53921_ = ~new_n53552_ & new_n53920_;
  assign new_n53922_ = ~new_n53919_ & ~new_n53921_;
  assign new_n53923_ = ~\b[19]  & ~new_n53922_;
  assign new_n53924_ = ~new_n53115_ & new_n53329_;
  assign new_n53925_ = ~new_n53325_ & new_n53924_;
  assign new_n53926_ = ~new_n53326_ & ~new_n53329_;
  assign new_n53927_ = ~new_n53925_ & ~new_n53926_;
  assign new_n53928_ = ~new_n53554_ & ~new_n53927_;
  assign new_n53929_ = ~new_n53105_ & ~new_n53553_;
  assign new_n53930_ = ~new_n53552_ & new_n53929_;
  assign new_n53931_ = ~new_n53928_ & ~new_n53930_;
  assign new_n53932_ = ~\b[18]  & ~new_n53931_;
  assign new_n53933_ = ~new_n53124_ & new_n53324_;
  assign new_n53934_ = ~new_n53320_ & new_n53933_;
  assign new_n53935_ = ~new_n53321_ & ~new_n53324_;
  assign new_n53936_ = ~new_n53934_ & ~new_n53935_;
  assign new_n53937_ = ~new_n53554_ & ~new_n53936_;
  assign new_n53938_ = ~new_n53114_ & ~new_n53553_;
  assign new_n53939_ = ~new_n53552_ & new_n53938_;
  assign new_n53940_ = ~new_n53937_ & ~new_n53939_;
  assign new_n53941_ = ~\b[17]  & ~new_n53940_;
  assign new_n53942_ = ~new_n53133_ & new_n53319_;
  assign new_n53943_ = ~new_n53315_ & new_n53942_;
  assign new_n53944_ = ~new_n53316_ & ~new_n53319_;
  assign new_n53945_ = ~new_n53943_ & ~new_n53944_;
  assign new_n53946_ = ~new_n53554_ & ~new_n53945_;
  assign new_n53947_ = ~new_n53123_ & ~new_n53553_;
  assign new_n53948_ = ~new_n53552_ & new_n53947_;
  assign new_n53949_ = ~new_n53946_ & ~new_n53948_;
  assign new_n53950_ = ~\b[16]  & ~new_n53949_;
  assign new_n53951_ = ~new_n53142_ & new_n53314_;
  assign new_n53952_ = ~new_n53310_ & new_n53951_;
  assign new_n53953_ = ~new_n53311_ & ~new_n53314_;
  assign new_n53954_ = ~new_n53952_ & ~new_n53953_;
  assign new_n53955_ = ~new_n53554_ & ~new_n53954_;
  assign new_n53956_ = ~new_n53132_ & ~new_n53553_;
  assign new_n53957_ = ~new_n53552_ & new_n53956_;
  assign new_n53958_ = ~new_n53955_ & ~new_n53957_;
  assign new_n53959_ = ~\b[15]  & ~new_n53958_;
  assign new_n53960_ = ~new_n53151_ & new_n53309_;
  assign new_n53961_ = ~new_n53305_ & new_n53960_;
  assign new_n53962_ = ~new_n53306_ & ~new_n53309_;
  assign new_n53963_ = ~new_n53961_ & ~new_n53962_;
  assign new_n53964_ = ~new_n53554_ & ~new_n53963_;
  assign new_n53965_ = ~new_n53141_ & ~new_n53553_;
  assign new_n53966_ = ~new_n53552_ & new_n53965_;
  assign new_n53967_ = ~new_n53964_ & ~new_n53966_;
  assign new_n53968_ = ~\b[14]  & ~new_n53967_;
  assign new_n53969_ = ~new_n53160_ & new_n53304_;
  assign new_n53970_ = ~new_n53300_ & new_n53969_;
  assign new_n53971_ = ~new_n53301_ & ~new_n53304_;
  assign new_n53972_ = ~new_n53970_ & ~new_n53971_;
  assign new_n53973_ = ~new_n53554_ & ~new_n53972_;
  assign new_n53974_ = ~new_n53150_ & ~new_n53553_;
  assign new_n53975_ = ~new_n53552_ & new_n53974_;
  assign new_n53976_ = ~new_n53973_ & ~new_n53975_;
  assign new_n53977_ = ~\b[13]  & ~new_n53976_;
  assign new_n53978_ = ~new_n53169_ & new_n53299_;
  assign new_n53979_ = ~new_n53295_ & new_n53978_;
  assign new_n53980_ = ~new_n53296_ & ~new_n53299_;
  assign new_n53981_ = ~new_n53979_ & ~new_n53980_;
  assign new_n53982_ = ~new_n53554_ & ~new_n53981_;
  assign new_n53983_ = ~new_n53159_ & ~new_n53553_;
  assign new_n53984_ = ~new_n53552_ & new_n53983_;
  assign new_n53985_ = ~new_n53982_ & ~new_n53984_;
  assign new_n53986_ = ~\b[12]  & ~new_n53985_;
  assign new_n53987_ = ~new_n53178_ & new_n53294_;
  assign new_n53988_ = ~new_n53290_ & new_n53987_;
  assign new_n53989_ = ~new_n53291_ & ~new_n53294_;
  assign new_n53990_ = ~new_n53988_ & ~new_n53989_;
  assign new_n53991_ = ~new_n53554_ & ~new_n53990_;
  assign new_n53992_ = ~new_n53168_ & ~new_n53553_;
  assign new_n53993_ = ~new_n53552_ & new_n53992_;
  assign new_n53994_ = ~new_n53991_ & ~new_n53993_;
  assign new_n53995_ = ~\b[11]  & ~new_n53994_;
  assign new_n53996_ = ~new_n53187_ & new_n53289_;
  assign new_n53997_ = ~new_n53285_ & new_n53996_;
  assign new_n53998_ = ~new_n53286_ & ~new_n53289_;
  assign new_n53999_ = ~new_n53997_ & ~new_n53998_;
  assign new_n54000_ = ~new_n53554_ & ~new_n53999_;
  assign new_n54001_ = ~new_n53177_ & ~new_n53553_;
  assign new_n54002_ = ~new_n53552_ & new_n54001_;
  assign new_n54003_ = ~new_n54000_ & ~new_n54002_;
  assign new_n54004_ = ~\b[10]  & ~new_n54003_;
  assign new_n54005_ = ~new_n53196_ & new_n53284_;
  assign new_n54006_ = ~new_n53280_ & new_n54005_;
  assign new_n54007_ = ~new_n53281_ & ~new_n53284_;
  assign new_n54008_ = ~new_n54006_ & ~new_n54007_;
  assign new_n54009_ = ~new_n53554_ & ~new_n54008_;
  assign new_n54010_ = ~new_n53186_ & ~new_n53553_;
  assign new_n54011_ = ~new_n53552_ & new_n54010_;
  assign new_n54012_ = ~new_n54009_ & ~new_n54011_;
  assign new_n54013_ = ~\b[9]  & ~new_n54012_;
  assign new_n54014_ = ~new_n53205_ & new_n53279_;
  assign new_n54015_ = ~new_n53275_ & new_n54014_;
  assign new_n54016_ = ~new_n53276_ & ~new_n53279_;
  assign new_n54017_ = ~new_n54015_ & ~new_n54016_;
  assign new_n54018_ = ~new_n53554_ & ~new_n54017_;
  assign new_n54019_ = ~new_n53195_ & ~new_n53553_;
  assign new_n54020_ = ~new_n53552_ & new_n54019_;
  assign new_n54021_ = ~new_n54018_ & ~new_n54020_;
  assign new_n54022_ = ~\b[8]  & ~new_n54021_;
  assign new_n54023_ = ~new_n53214_ & new_n53274_;
  assign new_n54024_ = ~new_n53270_ & new_n54023_;
  assign new_n54025_ = ~new_n53271_ & ~new_n53274_;
  assign new_n54026_ = ~new_n54024_ & ~new_n54025_;
  assign new_n54027_ = ~new_n53554_ & ~new_n54026_;
  assign new_n54028_ = ~new_n53204_ & ~new_n53553_;
  assign new_n54029_ = ~new_n53552_ & new_n54028_;
  assign new_n54030_ = ~new_n54027_ & ~new_n54029_;
  assign new_n54031_ = ~\b[7]  & ~new_n54030_;
  assign new_n54032_ = ~new_n53223_ & new_n53269_;
  assign new_n54033_ = ~new_n53265_ & new_n54032_;
  assign new_n54034_ = ~new_n53266_ & ~new_n53269_;
  assign new_n54035_ = ~new_n54033_ & ~new_n54034_;
  assign new_n54036_ = ~new_n53554_ & ~new_n54035_;
  assign new_n54037_ = ~new_n53213_ & ~new_n53553_;
  assign new_n54038_ = ~new_n53552_ & new_n54037_;
  assign new_n54039_ = ~new_n54036_ & ~new_n54038_;
  assign new_n54040_ = ~\b[6]  & ~new_n54039_;
  assign new_n54041_ = ~new_n53232_ & new_n53264_;
  assign new_n54042_ = ~new_n53260_ & new_n54041_;
  assign new_n54043_ = ~new_n53261_ & ~new_n53264_;
  assign new_n54044_ = ~new_n54042_ & ~new_n54043_;
  assign new_n54045_ = ~new_n53554_ & ~new_n54044_;
  assign new_n54046_ = ~new_n53222_ & ~new_n53553_;
  assign new_n54047_ = ~new_n53552_ & new_n54046_;
  assign new_n54048_ = ~new_n54045_ & ~new_n54047_;
  assign new_n54049_ = ~\b[5]  & ~new_n54048_;
  assign new_n54050_ = ~new_n53240_ & new_n53259_;
  assign new_n54051_ = ~new_n53255_ & new_n54050_;
  assign new_n54052_ = ~new_n53256_ & ~new_n53259_;
  assign new_n54053_ = ~new_n54051_ & ~new_n54052_;
  assign new_n54054_ = ~new_n53554_ & ~new_n54053_;
  assign new_n54055_ = ~new_n53231_ & ~new_n53553_;
  assign new_n54056_ = ~new_n53552_ & new_n54055_;
  assign new_n54057_ = ~new_n54054_ & ~new_n54056_;
  assign new_n54058_ = ~\b[4]  & ~new_n54057_;
  assign new_n54059_ = ~new_n53250_ & new_n53254_;
  assign new_n54060_ = ~new_n53249_ & new_n54059_;
  assign new_n54061_ = ~new_n53251_ & ~new_n53254_;
  assign new_n54062_ = ~new_n54060_ & ~new_n54061_;
  assign new_n54063_ = ~new_n53554_ & ~new_n54062_;
  assign new_n54064_ = ~new_n53239_ & ~new_n53553_;
  assign new_n54065_ = ~new_n53552_ & new_n54064_;
  assign new_n54066_ = ~new_n54063_ & ~new_n54065_;
  assign new_n54067_ = ~\b[3]  & ~new_n54066_;
  assign new_n54068_ = new_n25233_ & ~new_n53247_;
  assign new_n54069_ = ~new_n53245_ & new_n54068_;
  assign new_n54070_ = ~new_n53249_ & ~new_n54069_;
  assign new_n54071_ = ~new_n53554_ & new_n54070_;
  assign new_n54072_ = ~new_n53244_ & ~new_n53553_;
  assign new_n54073_ = ~new_n53552_ & new_n54072_;
  assign new_n54074_ = ~new_n54071_ & ~new_n54073_;
  assign new_n54075_ = ~\b[2]  & ~new_n54074_;
  assign new_n54076_ = \b[0]  & ~new_n53554_;
  assign new_n54077_ = \a[4]  & ~new_n54076_;
  assign new_n54078_ = new_n25233_ & ~new_n53554_;
  assign new_n54079_ = ~new_n54077_ & ~new_n54078_;
  assign new_n54080_ = \b[1]  & ~new_n54079_;
  assign new_n54081_ = ~\b[1]  & ~new_n54078_;
  assign new_n54082_ = ~new_n54077_ & new_n54081_;
  assign new_n54083_ = ~new_n54080_ & ~new_n54082_;
  assign new_n54084_ = ~new_n26069_ & ~new_n54083_;
  assign new_n54085_ = ~\b[1]  & ~new_n54079_;
  assign new_n54086_ = ~new_n54084_ & ~new_n54085_;
  assign new_n54087_ = \b[2]  & ~new_n54073_;
  assign new_n54088_ = ~new_n54071_ & new_n54087_;
  assign new_n54089_ = ~new_n54075_ & ~new_n54088_;
  assign new_n54090_ = ~new_n54086_ & new_n54089_;
  assign new_n54091_ = ~new_n54075_ & ~new_n54090_;
  assign new_n54092_ = \b[3]  & ~new_n54065_;
  assign new_n54093_ = ~new_n54063_ & new_n54092_;
  assign new_n54094_ = ~new_n54067_ & ~new_n54093_;
  assign new_n54095_ = ~new_n54091_ & new_n54094_;
  assign new_n54096_ = ~new_n54067_ & ~new_n54095_;
  assign new_n54097_ = \b[4]  & ~new_n54056_;
  assign new_n54098_ = ~new_n54054_ & new_n54097_;
  assign new_n54099_ = ~new_n54058_ & ~new_n54098_;
  assign new_n54100_ = ~new_n54096_ & new_n54099_;
  assign new_n54101_ = ~new_n54058_ & ~new_n54100_;
  assign new_n54102_ = \b[5]  & ~new_n54047_;
  assign new_n54103_ = ~new_n54045_ & new_n54102_;
  assign new_n54104_ = ~new_n54049_ & ~new_n54103_;
  assign new_n54105_ = ~new_n54101_ & new_n54104_;
  assign new_n54106_ = ~new_n54049_ & ~new_n54105_;
  assign new_n54107_ = \b[6]  & ~new_n54038_;
  assign new_n54108_ = ~new_n54036_ & new_n54107_;
  assign new_n54109_ = ~new_n54040_ & ~new_n54108_;
  assign new_n54110_ = ~new_n54106_ & new_n54109_;
  assign new_n54111_ = ~new_n54040_ & ~new_n54110_;
  assign new_n54112_ = \b[7]  & ~new_n54029_;
  assign new_n54113_ = ~new_n54027_ & new_n54112_;
  assign new_n54114_ = ~new_n54031_ & ~new_n54113_;
  assign new_n54115_ = ~new_n54111_ & new_n54114_;
  assign new_n54116_ = ~new_n54031_ & ~new_n54115_;
  assign new_n54117_ = \b[8]  & ~new_n54020_;
  assign new_n54118_ = ~new_n54018_ & new_n54117_;
  assign new_n54119_ = ~new_n54022_ & ~new_n54118_;
  assign new_n54120_ = ~new_n54116_ & new_n54119_;
  assign new_n54121_ = ~new_n54022_ & ~new_n54120_;
  assign new_n54122_ = \b[9]  & ~new_n54011_;
  assign new_n54123_ = ~new_n54009_ & new_n54122_;
  assign new_n54124_ = ~new_n54013_ & ~new_n54123_;
  assign new_n54125_ = ~new_n54121_ & new_n54124_;
  assign new_n54126_ = ~new_n54013_ & ~new_n54125_;
  assign new_n54127_ = \b[10]  & ~new_n54002_;
  assign new_n54128_ = ~new_n54000_ & new_n54127_;
  assign new_n54129_ = ~new_n54004_ & ~new_n54128_;
  assign new_n54130_ = ~new_n54126_ & new_n54129_;
  assign new_n54131_ = ~new_n54004_ & ~new_n54130_;
  assign new_n54132_ = \b[11]  & ~new_n53993_;
  assign new_n54133_ = ~new_n53991_ & new_n54132_;
  assign new_n54134_ = ~new_n53995_ & ~new_n54133_;
  assign new_n54135_ = ~new_n54131_ & new_n54134_;
  assign new_n54136_ = ~new_n53995_ & ~new_n54135_;
  assign new_n54137_ = \b[12]  & ~new_n53984_;
  assign new_n54138_ = ~new_n53982_ & new_n54137_;
  assign new_n54139_ = ~new_n53986_ & ~new_n54138_;
  assign new_n54140_ = ~new_n54136_ & new_n54139_;
  assign new_n54141_ = ~new_n53986_ & ~new_n54140_;
  assign new_n54142_ = \b[13]  & ~new_n53975_;
  assign new_n54143_ = ~new_n53973_ & new_n54142_;
  assign new_n54144_ = ~new_n53977_ & ~new_n54143_;
  assign new_n54145_ = ~new_n54141_ & new_n54144_;
  assign new_n54146_ = ~new_n53977_ & ~new_n54145_;
  assign new_n54147_ = \b[14]  & ~new_n53966_;
  assign new_n54148_ = ~new_n53964_ & new_n54147_;
  assign new_n54149_ = ~new_n53968_ & ~new_n54148_;
  assign new_n54150_ = ~new_n54146_ & new_n54149_;
  assign new_n54151_ = ~new_n53968_ & ~new_n54150_;
  assign new_n54152_ = \b[15]  & ~new_n53957_;
  assign new_n54153_ = ~new_n53955_ & new_n54152_;
  assign new_n54154_ = ~new_n53959_ & ~new_n54153_;
  assign new_n54155_ = ~new_n54151_ & new_n54154_;
  assign new_n54156_ = ~new_n53959_ & ~new_n54155_;
  assign new_n54157_ = \b[16]  & ~new_n53948_;
  assign new_n54158_ = ~new_n53946_ & new_n54157_;
  assign new_n54159_ = ~new_n53950_ & ~new_n54158_;
  assign new_n54160_ = ~new_n54156_ & new_n54159_;
  assign new_n54161_ = ~new_n53950_ & ~new_n54160_;
  assign new_n54162_ = \b[17]  & ~new_n53939_;
  assign new_n54163_ = ~new_n53937_ & new_n54162_;
  assign new_n54164_ = ~new_n53941_ & ~new_n54163_;
  assign new_n54165_ = ~new_n54161_ & new_n54164_;
  assign new_n54166_ = ~new_n53941_ & ~new_n54165_;
  assign new_n54167_ = \b[18]  & ~new_n53930_;
  assign new_n54168_ = ~new_n53928_ & new_n54167_;
  assign new_n54169_ = ~new_n53932_ & ~new_n54168_;
  assign new_n54170_ = ~new_n54166_ & new_n54169_;
  assign new_n54171_ = ~new_n53932_ & ~new_n54170_;
  assign new_n54172_ = \b[19]  & ~new_n53921_;
  assign new_n54173_ = ~new_n53919_ & new_n54172_;
  assign new_n54174_ = ~new_n53923_ & ~new_n54173_;
  assign new_n54175_ = ~new_n54171_ & new_n54174_;
  assign new_n54176_ = ~new_n53923_ & ~new_n54175_;
  assign new_n54177_ = \b[20]  & ~new_n53912_;
  assign new_n54178_ = ~new_n53910_ & new_n54177_;
  assign new_n54179_ = ~new_n53914_ & ~new_n54178_;
  assign new_n54180_ = ~new_n54176_ & new_n54179_;
  assign new_n54181_ = ~new_n53914_ & ~new_n54180_;
  assign new_n54182_ = \b[21]  & ~new_n53903_;
  assign new_n54183_ = ~new_n53901_ & new_n54182_;
  assign new_n54184_ = ~new_n53905_ & ~new_n54183_;
  assign new_n54185_ = ~new_n54181_ & new_n54184_;
  assign new_n54186_ = ~new_n53905_ & ~new_n54185_;
  assign new_n54187_ = \b[22]  & ~new_n53894_;
  assign new_n54188_ = ~new_n53892_ & new_n54187_;
  assign new_n54189_ = ~new_n53896_ & ~new_n54188_;
  assign new_n54190_ = ~new_n54186_ & new_n54189_;
  assign new_n54191_ = ~new_n53896_ & ~new_n54190_;
  assign new_n54192_ = \b[23]  & ~new_n53885_;
  assign new_n54193_ = ~new_n53883_ & new_n54192_;
  assign new_n54194_ = ~new_n53887_ & ~new_n54193_;
  assign new_n54195_ = ~new_n54191_ & new_n54194_;
  assign new_n54196_ = ~new_n53887_ & ~new_n54195_;
  assign new_n54197_ = \b[24]  & ~new_n53876_;
  assign new_n54198_ = ~new_n53874_ & new_n54197_;
  assign new_n54199_ = ~new_n53878_ & ~new_n54198_;
  assign new_n54200_ = ~new_n54196_ & new_n54199_;
  assign new_n54201_ = ~new_n53878_ & ~new_n54200_;
  assign new_n54202_ = \b[25]  & ~new_n53867_;
  assign new_n54203_ = ~new_n53865_ & new_n54202_;
  assign new_n54204_ = ~new_n53869_ & ~new_n54203_;
  assign new_n54205_ = ~new_n54201_ & new_n54204_;
  assign new_n54206_ = ~new_n53869_ & ~new_n54205_;
  assign new_n54207_ = \b[26]  & ~new_n53858_;
  assign new_n54208_ = ~new_n53856_ & new_n54207_;
  assign new_n54209_ = ~new_n53860_ & ~new_n54208_;
  assign new_n54210_ = ~new_n54206_ & new_n54209_;
  assign new_n54211_ = ~new_n53860_ & ~new_n54210_;
  assign new_n54212_ = \b[27]  & ~new_n53849_;
  assign new_n54213_ = ~new_n53847_ & new_n54212_;
  assign new_n54214_ = ~new_n53851_ & ~new_n54213_;
  assign new_n54215_ = ~new_n54211_ & new_n54214_;
  assign new_n54216_ = ~new_n53851_ & ~new_n54215_;
  assign new_n54217_ = \b[28]  & ~new_n53840_;
  assign new_n54218_ = ~new_n53838_ & new_n54217_;
  assign new_n54219_ = ~new_n53842_ & ~new_n54218_;
  assign new_n54220_ = ~new_n54216_ & new_n54219_;
  assign new_n54221_ = ~new_n53842_ & ~new_n54220_;
  assign new_n54222_ = \b[29]  & ~new_n53831_;
  assign new_n54223_ = ~new_n53829_ & new_n54222_;
  assign new_n54224_ = ~new_n53833_ & ~new_n54223_;
  assign new_n54225_ = ~new_n54221_ & new_n54224_;
  assign new_n54226_ = ~new_n53833_ & ~new_n54225_;
  assign new_n54227_ = \b[30]  & ~new_n53822_;
  assign new_n54228_ = ~new_n53820_ & new_n54227_;
  assign new_n54229_ = ~new_n53824_ & ~new_n54228_;
  assign new_n54230_ = ~new_n54226_ & new_n54229_;
  assign new_n54231_ = ~new_n53824_ & ~new_n54230_;
  assign new_n54232_ = \b[31]  & ~new_n53813_;
  assign new_n54233_ = ~new_n53811_ & new_n54232_;
  assign new_n54234_ = ~new_n53815_ & ~new_n54233_;
  assign new_n54235_ = ~new_n54231_ & new_n54234_;
  assign new_n54236_ = ~new_n53815_ & ~new_n54235_;
  assign new_n54237_ = \b[32]  & ~new_n53804_;
  assign new_n54238_ = ~new_n53802_ & new_n54237_;
  assign new_n54239_ = ~new_n53806_ & ~new_n54238_;
  assign new_n54240_ = ~new_n54236_ & new_n54239_;
  assign new_n54241_ = ~new_n53806_ & ~new_n54240_;
  assign new_n54242_ = \b[33]  & ~new_n53795_;
  assign new_n54243_ = ~new_n53793_ & new_n54242_;
  assign new_n54244_ = ~new_n53797_ & ~new_n54243_;
  assign new_n54245_ = ~new_n54241_ & new_n54244_;
  assign new_n54246_ = ~new_n53797_ & ~new_n54245_;
  assign new_n54247_ = \b[34]  & ~new_n53786_;
  assign new_n54248_ = ~new_n53784_ & new_n54247_;
  assign new_n54249_ = ~new_n53788_ & ~new_n54248_;
  assign new_n54250_ = ~new_n54246_ & new_n54249_;
  assign new_n54251_ = ~new_n53788_ & ~new_n54250_;
  assign new_n54252_ = \b[35]  & ~new_n53777_;
  assign new_n54253_ = ~new_n53775_ & new_n54252_;
  assign new_n54254_ = ~new_n53779_ & ~new_n54253_;
  assign new_n54255_ = ~new_n54251_ & new_n54254_;
  assign new_n54256_ = ~new_n53779_ & ~new_n54255_;
  assign new_n54257_ = \b[36]  & ~new_n53768_;
  assign new_n54258_ = ~new_n53766_ & new_n54257_;
  assign new_n54259_ = ~new_n53770_ & ~new_n54258_;
  assign new_n54260_ = ~new_n54256_ & new_n54259_;
  assign new_n54261_ = ~new_n53770_ & ~new_n54260_;
  assign new_n54262_ = \b[37]  & ~new_n53759_;
  assign new_n54263_ = ~new_n53757_ & new_n54262_;
  assign new_n54264_ = ~new_n53761_ & ~new_n54263_;
  assign new_n54265_ = ~new_n54261_ & new_n54264_;
  assign new_n54266_ = ~new_n53761_ & ~new_n54265_;
  assign new_n54267_ = \b[38]  & ~new_n53750_;
  assign new_n54268_ = ~new_n53748_ & new_n54267_;
  assign new_n54269_ = ~new_n53752_ & ~new_n54268_;
  assign new_n54270_ = ~new_n54266_ & new_n54269_;
  assign new_n54271_ = ~new_n53752_ & ~new_n54270_;
  assign new_n54272_ = \b[39]  & ~new_n53741_;
  assign new_n54273_ = ~new_n53739_ & new_n54272_;
  assign new_n54274_ = ~new_n53743_ & ~new_n54273_;
  assign new_n54275_ = ~new_n54271_ & new_n54274_;
  assign new_n54276_ = ~new_n53743_ & ~new_n54275_;
  assign new_n54277_ = \b[40]  & ~new_n53732_;
  assign new_n54278_ = ~new_n53730_ & new_n54277_;
  assign new_n54279_ = ~new_n53734_ & ~new_n54278_;
  assign new_n54280_ = ~new_n54276_ & new_n54279_;
  assign new_n54281_ = ~new_n53734_ & ~new_n54280_;
  assign new_n54282_ = \b[41]  & ~new_n53723_;
  assign new_n54283_ = ~new_n53721_ & new_n54282_;
  assign new_n54284_ = ~new_n53725_ & ~new_n54283_;
  assign new_n54285_ = ~new_n54281_ & new_n54284_;
  assign new_n54286_ = ~new_n53725_ & ~new_n54285_;
  assign new_n54287_ = \b[42]  & ~new_n53714_;
  assign new_n54288_ = ~new_n53712_ & new_n54287_;
  assign new_n54289_ = ~new_n53716_ & ~new_n54288_;
  assign new_n54290_ = ~new_n54286_ & new_n54289_;
  assign new_n54291_ = ~new_n53716_ & ~new_n54290_;
  assign new_n54292_ = \b[43]  & ~new_n53705_;
  assign new_n54293_ = ~new_n53703_ & new_n54292_;
  assign new_n54294_ = ~new_n53707_ & ~new_n54293_;
  assign new_n54295_ = ~new_n54291_ & new_n54294_;
  assign new_n54296_ = ~new_n53707_ & ~new_n54295_;
  assign new_n54297_ = \b[44]  & ~new_n53696_;
  assign new_n54298_ = ~new_n53694_ & new_n54297_;
  assign new_n54299_ = ~new_n53698_ & ~new_n54298_;
  assign new_n54300_ = ~new_n54296_ & new_n54299_;
  assign new_n54301_ = ~new_n53698_ & ~new_n54300_;
  assign new_n54302_ = \b[45]  & ~new_n53687_;
  assign new_n54303_ = ~new_n53685_ & new_n54302_;
  assign new_n54304_ = ~new_n53689_ & ~new_n54303_;
  assign new_n54305_ = ~new_n54301_ & new_n54304_;
  assign new_n54306_ = ~new_n53689_ & ~new_n54305_;
  assign new_n54307_ = \b[46]  & ~new_n53678_;
  assign new_n54308_ = ~new_n53676_ & new_n54307_;
  assign new_n54309_ = ~new_n53680_ & ~new_n54308_;
  assign new_n54310_ = ~new_n54306_ & new_n54309_;
  assign new_n54311_ = ~new_n53680_ & ~new_n54310_;
  assign new_n54312_ = \b[47]  & ~new_n53669_;
  assign new_n54313_ = ~new_n53667_ & new_n54312_;
  assign new_n54314_ = ~new_n53671_ & ~new_n54313_;
  assign new_n54315_ = ~new_n54311_ & new_n54314_;
  assign new_n54316_ = ~new_n53671_ & ~new_n54315_;
  assign new_n54317_ = \b[48]  & ~new_n53660_;
  assign new_n54318_ = ~new_n53658_ & new_n54317_;
  assign new_n54319_ = ~new_n53662_ & ~new_n54318_;
  assign new_n54320_ = ~new_n54316_ & new_n54319_;
  assign new_n54321_ = ~new_n53662_ & ~new_n54320_;
  assign new_n54322_ = \b[49]  & ~new_n53651_;
  assign new_n54323_ = ~new_n53649_ & new_n54322_;
  assign new_n54324_ = ~new_n53653_ & ~new_n54323_;
  assign new_n54325_ = ~new_n54321_ & new_n54324_;
  assign new_n54326_ = ~new_n53653_ & ~new_n54325_;
  assign new_n54327_ = \b[50]  & ~new_n53642_;
  assign new_n54328_ = ~new_n53640_ & new_n54327_;
  assign new_n54329_ = ~new_n53644_ & ~new_n54328_;
  assign new_n54330_ = ~new_n54326_ & new_n54329_;
  assign new_n54331_ = ~new_n53644_ & ~new_n54330_;
  assign new_n54332_ = \b[51]  & ~new_n53633_;
  assign new_n54333_ = ~new_n53631_ & new_n54332_;
  assign new_n54334_ = ~new_n53635_ & ~new_n54333_;
  assign new_n54335_ = ~new_n54331_ & new_n54334_;
  assign new_n54336_ = ~new_n53635_ & ~new_n54335_;
  assign new_n54337_ = \b[52]  & ~new_n53624_;
  assign new_n54338_ = ~new_n53622_ & new_n54337_;
  assign new_n54339_ = ~new_n53626_ & ~new_n54338_;
  assign new_n54340_ = ~new_n54336_ & new_n54339_;
  assign new_n54341_ = ~new_n53626_ & ~new_n54340_;
  assign new_n54342_ = \b[53]  & ~new_n53615_;
  assign new_n54343_ = ~new_n53613_ & new_n54342_;
  assign new_n54344_ = ~new_n53617_ & ~new_n54343_;
  assign new_n54345_ = ~new_n54341_ & new_n54344_;
  assign new_n54346_ = ~new_n53617_ & ~new_n54345_;
  assign new_n54347_ = \b[54]  & ~new_n53606_;
  assign new_n54348_ = ~new_n53604_ & new_n54347_;
  assign new_n54349_ = ~new_n53608_ & ~new_n54348_;
  assign new_n54350_ = ~new_n54346_ & new_n54349_;
  assign new_n54351_ = ~new_n53608_ & ~new_n54350_;
  assign new_n54352_ = \b[55]  & ~new_n53597_;
  assign new_n54353_ = ~new_n53595_ & new_n54352_;
  assign new_n54354_ = ~new_n53599_ & ~new_n54353_;
  assign new_n54355_ = ~new_n54351_ & new_n54354_;
  assign new_n54356_ = ~new_n53599_ & ~new_n54355_;
  assign new_n54357_ = \b[56]  & ~new_n53588_;
  assign new_n54358_ = ~new_n53586_ & new_n54357_;
  assign new_n54359_ = ~new_n53590_ & ~new_n54358_;
  assign new_n54360_ = ~new_n54356_ & new_n54359_;
  assign new_n54361_ = ~new_n53590_ & ~new_n54360_;
  assign new_n54362_ = \b[57]  & ~new_n53579_;
  assign new_n54363_ = ~new_n53577_ & new_n54362_;
  assign new_n54364_ = ~new_n53581_ & ~new_n54363_;
  assign new_n54365_ = ~new_n54361_ & new_n54364_;
  assign new_n54366_ = ~new_n53581_ & ~new_n54365_;
  assign new_n54367_ = \b[58]  & ~new_n53570_;
  assign new_n54368_ = ~new_n53568_ & new_n54367_;
  assign new_n54369_ = ~new_n53572_ & ~new_n54368_;
  assign new_n54370_ = ~new_n54366_ & new_n54369_;
  assign new_n54371_ = ~new_n53572_ & ~new_n54370_;
  assign new_n54372_ = \b[59]  & ~new_n53561_;
  assign new_n54373_ = ~new_n53559_ & new_n54372_;
  assign new_n54374_ = ~new_n53563_ & ~new_n54373_;
  assign new_n54375_ = ~new_n54371_ & new_n54374_;
  assign new_n54376_ = ~new_n53563_ & ~new_n54375_;
  assign new_n54377_ = ~new_n52737_ & ~new_n53549_;
  assign new_n54378_ = ~new_n53547_ & new_n54377_;
  assign new_n54379_ = ~new_n53535_ & new_n54378_;
  assign new_n54380_ = ~new_n53547_ & ~new_n53549_;
  assign new_n54381_ = ~new_n53536_ & ~new_n54380_;
  assign new_n54382_ = ~new_n54379_ & ~new_n54381_;
  assign new_n54383_ = ~new_n53554_ & ~new_n54382_;
  assign new_n54384_ = ~new_n53546_ & ~new_n53553_;
  assign new_n54385_ = ~new_n53552_ & new_n54384_;
  assign new_n54386_ = ~new_n54383_ & ~new_n54385_;
  assign new_n54387_ = ~\b[60]  & ~new_n54386_;
  assign new_n54388_ = \b[60]  & ~new_n54385_;
  assign new_n54389_ = ~new_n54383_ & new_n54388_;
  assign new_n54390_ = new_n403_ & ~new_n54389_;
  assign new_n54391_ = ~new_n54387_ & new_n54390_;
  assign new_n54392_ = ~new_n54376_ & new_n54391_;
  assign new_n54393_ = new_n280_ & ~new_n54386_;
  assign new_n54394_ = ~new_n54392_ & ~new_n54393_;
  assign new_n54395_ = ~new_n53572_ & new_n54374_;
  assign new_n54396_ = ~new_n54370_ & new_n54395_;
  assign new_n54397_ = ~new_n54371_ & ~new_n54374_;
  assign new_n54398_ = ~new_n54396_ & ~new_n54397_;
  assign new_n54399_ = ~new_n54394_ & ~new_n54398_;
  assign new_n54400_ = ~new_n53562_ & ~new_n54393_;
  assign new_n54401_ = ~new_n54392_ & new_n54400_;
  assign new_n54402_ = ~new_n54399_ & ~new_n54401_;
  assign new_n54403_ = ~\b[60]  & ~new_n54402_;
  assign new_n54404_ = ~new_n53581_ & new_n54369_;
  assign new_n54405_ = ~new_n54365_ & new_n54404_;
  assign new_n54406_ = ~new_n54366_ & ~new_n54369_;
  assign new_n54407_ = ~new_n54405_ & ~new_n54406_;
  assign new_n54408_ = ~new_n54394_ & ~new_n54407_;
  assign new_n54409_ = ~new_n53571_ & ~new_n54393_;
  assign new_n54410_ = ~new_n54392_ & new_n54409_;
  assign new_n54411_ = ~new_n54408_ & ~new_n54410_;
  assign new_n54412_ = ~\b[59]  & ~new_n54411_;
  assign new_n54413_ = ~new_n53590_ & new_n54364_;
  assign new_n54414_ = ~new_n54360_ & new_n54413_;
  assign new_n54415_ = ~new_n54361_ & ~new_n54364_;
  assign new_n54416_ = ~new_n54414_ & ~new_n54415_;
  assign new_n54417_ = ~new_n54394_ & ~new_n54416_;
  assign new_n54418_ = ~new_n53580_ & ~new_n54393_;
  assign new_n54419_ = ~new_n54392_ & new_n54418_;
  assign new_n54420_ = ~new_n54417_ & ~new_n54419_;
  assign new_n54421_ = ~\b[58]  & ~new_n54420_;
  assign new_n54422_ = ~new_n53599_ & new_n54359_;
  assign new_n54423_ = ~new_n54355_ & new_n54422_;
  assign new_n54424_ = ~new_n54356_ & ~new_n54359_;
  assign new_n54425_ = ~new_n54423_ & ~new_n54424_;
  assign new_n54426_ = ~new_n54394_ & ~new_n54425_;
  assign new_n54427_ = ~new_n53589_ & ~new_n54393_;
  assign new_n54428_ = ~new_n54392_ & new_n54427_;
  assign new_n54429_ = ~new_n54426_ & ~new_n54428_;
  assign new_n54430_ = ~\b[57]  & ~new_n54429_;
  assign new_n54431_ = ~new_n53608_ & new_n54354_;
  assign new_n54432_ = ~new_n54350_ & new_n54431_;
  assign new_n54433_ = ~new_n54351_ & ~new_n54354_;
  assign new_n54434_ = ~new_n54432_ & ~new_n54433_;
  assign new_n54435_ = ~new_n54394_ & ~new_n54434_;
  assign new_n54436_ = ~new_n53598_ & ~new_n54393_;
  assign new_n54437_ = ~new_n54392_ & new_n54436_;
  assign new_n54438_ = ~new_n54435_ & ~new_n54437_;
  assign new_n54439_ = ~\b[56]  & ~new_n54438_;
  assign new_n54440_ = ~new_n53617_ & new_n54349_;
  assign new_n54441_ = ~new_n54345_ & new_n54440_;
  assign new_n54442_ = ~new_n54346_ & ~new_n54349_;
  assign new_n54443_ = ~new_n54441_ & ~new_n54442_;
  assign new_n54444_ = ~new_n54394_ & ~new_n54443_;
  assign new_n54445_ = ~new_n53607_ & ~new_n54393_;
  assign new_n54446_ = ~new_n54392_ & new_n54445_;
  assign new_n54447_ = ~new_n54444_ & ~new_n54446_;
  assign new_n54448_ = ~\b[55]  & ~new_n54447_;
  assign new_n54449_ = ~new_n53626_ & new_n54344_;
  assign new_n54450_ = ~new_n54340_ & new_n54449_;
  assign new_n54451_ = ~new_n54341_ & ~new_n54344_;
  assign new_n54452_ = ~new_n54450_ & ~new_n54451_;
  assign new_n54453_ = ~new_n54394_ & ~new_n54452_;
  assign new_n54454_ = ~new_n53616_ & ~new_n54393_;
  assign new_n54455_ = ~new_n54392_ & new_n54454_;
  assign new_n54456_ = ~new_n54453_ & ~new_n54455_;
  assign new_n54457_ = ~\b[54]  & ~new_n54456_;
  assign new_n54458_ = ~new_n53635_ & new_n54339_;
  assign new_n54459_ = ~new_n54335_ & new_n54458_;
  assign new_n54460_ = ~new_n54336_ & ~new_n54339_;
  assign new_n54461_ = ~new_n54459_ & ~new_n54460_;
  assign new_n54462_ = ~new_n54394_ & ~new_n54461_;
  assign new_n54463_ = ~new_n53625_ & ~new_n54393_;
  assign new_n54464_ = ~new_n54392_ & new_n54463_;
  assign new_n54465_ = ~new_n54462_ & ~new_n54464_;
  assign new_n54466_ = ~\b[53]  & ~new_n54465_;
  assign new_n54467_ = ~new_n53644_ & new_n54334_;
  assign new_n54468_ = ~new_n54330_ & new_n54467_;
  assign new_n54469_ = ~new_n54331_ & ~new_n54334_;
  assign new_n54470_ = ~new_n54468_ & ~new_n54469_;
  assign new_n54471_ = ~new_n54394_ & ~new_n54470_;
  assign new_n54472_ = ~new_n53634_ & ~new_n54393_;
  assign new_n54473_ = ~new_n54392_ & new_n54472_;
  assign new_n54474_ = ~new_n54471_ & ~new_n54473_;
  assign new_n54475_ = ~\b[52]  & ~new_n54474_;
  assign new_n54476_ = ~new_n53653_ & new_n54329_;
  assign new_n54477_ = ~new_n54325_ & new_n54476_;
  assign new_n54478_ = ~new_n54326_ & ~new_n54329_;
  assign new_n54479_ = ~new_n54477_ & ~new_n54478_;
  assign new_n54480_ = ~new_n54394_ & ~new_n54479_;
  assign new_n54481_ = ~new_n53643_ & ~new_n54393_;
  assign new_n54482_ = ~new_n54392_ & new_n54481_;
  assign new_n54483_ = ~new_n54480_ & ~new_n54482_;
  assign new_n54484_ = ~\b[51]  & ~new_n54483_;
  assign new_n54485_ = ~new_n53662_ & new_n54324_;
  assign new_n54486_ = ~new_n54320_ & new_n54485_;
  assign new_n54487_ = ~new_n54321_ & ~new_n54324_;
  assign new_n54488_ = ~new_n54486_ & ~new_n54487_;
  assign new_n54489_ = ~new_n54394_ & ~new_n54488_;
  assign new_n54490_ = ~new_n53652_ & ~new_n54393_;
  assign new_n54491_ = ~new_n54392_ & new_n54490_;
  assign new_n54492_ = ~new_n54489_ & ~new_n54491_;
  assign new_n54493_ = ~\b[50]  & ~new_n54492_;
  assign new_n54494_ = ~new_n53671_ & new_n54319_;
  assign new_n54495_ = ~new_n54315_ & new_n54494_;
  assign new_n54496_ = ~new_n54316_ & ~new_n54319_;
  assign new_n54497_ = ~new_n54495_ & ~new_n54496_;
  assign new_n54498_ = ~new_n54394_ & ~new_n54497_;
  assign new_n54499_ = ~new_n53661_ & ~new_n54393_;
  assign new_n54500_ = ~new_n54392_ & new_n54499_;
  assign new_n54501_ = ~new_n54498_ & ~new_n54500_;
  assign new_n54502_ = ~\b[49]  & ~new_n54501_;
  assign new_n54503_ = ~new_n53680_ & new_n54314_;
  assign new_n54504_ = ~new_n54310_ & new_n54503_;
  assign new_n54505_ = ~new_n54311_ & ~new_n54314_;
  assign new_n54506_ = ~new_n54504_ & ~new_n54505_;
  assign new_n54507_ = ~new_n54394_ & ~new_n54506_;
  assign new_n54508_ = ~new_n53670_ & ~new_n54393_;
  assign new_n54509_ = ~new_n54392_ & new_n54508_;
  assign new_n54510_ = ~new_n54507_ & ~new_n54509_;
  assign new_n54511_ = ~\b[48]  & ~new_n54510_;
  assign new_n54512_ = ~new_n53689_ & new_n54309_;
  assign new_n54513_ = ~new_n54305_ & new_n54512_;
  assign new_n54514_ = ~new_n54306_ & ~new_n54309_;
  assign new_n54515_ = ~new_n54513_ & ~new_n54514_;
  assign new_n54516_ = ~new_n54394_ & ~new_n54515_;
  assign new_n54517_ = ~new_n53679_ & ~new_n54393_;
  assign new_n54518_ = ~new_n54392_ & new_n54517_;
  assign new_n54519_ = ~new_n54516_ & ~new_n54518_;
  assign new_n54520_ = ~\b[47]  & ~new_n54519_;
  assign new_n54521_ = ~new_n53698_ & new_n54304_;
  assign new_n54522_ = ~new_n54300_ & new_n54521_;
  assign new_n54523_ = ~new_n54301_ & ~new_n54304_;
  assign new_n54524_ = ~new_n54522_ & ~new_n54523_;
  assign new_n54525_ = ~new_n54394_ & ~new_n54524_;
  assign new_n54526_ = ~new_n53688_ & ~new_n54393_;
  assign new_n54527_ = ~new_n54392_ & new_n54526_;
  assign new_n54528_ = ~new_n54525_ & ~new_n54527_;
  assign new_n54529_ = ~\b[46]  & ~new_n54528_;
  assign new_n54530_ = ~new_n53707_ & new_n54299_;
  assign new_n54531_ = ~new_n54295_ & new_n54530_;
  assign new_n54532_ = ~new_n54296_ & ~new_n54299_;
  assign new_n54533_ = ~new_n54531_ & ~new_n54532_;
  assign new_n54534_ = ~new_n54394_ & ~new_n54533_;
  assign new_n54535_ = ~new_n53697_ & ~new_n54393_;
  assign new_n54536_ = ~new_n54392_ & new_n54535_;
  assign new_n54537_ = ~new_n54534_ & ~new_n54536_;
  assign new_n54538_ = ~\b[45]  & ~new_n54537_;
  assign new_n54539_ = ~new_n53716_ & new_n54294_;
  assign new_n54540_ = ~new_n54290_ & new_n54539_;
  assign new_n54541_ = ~new_n54291_ & ~new_n54294_;
  assign new_n54542_ = ~new_n54540_ & ~new_n54541_;
  assign new_n54543_ = ~new_n54394_ & ~new_n54542_;
  assign new_n54544_ = ~new_n53706_ & ~new_n54393_;
  assign new_n54545_ = ~new_n54392_ & new_n54544_;
  assign new_n54546_ = ~new_n54543_ & ~new_n54545_;
  assign new_n54547_ = ~\b[44]  & ~new_n54546_;
  assign new_n54548_ = ~new_n53725_ & new_n54289_;
  assign new_n54549_ = ~new_n54285_ & new_n54548_;
  assign new_n54550_ = ~new_n54286_ & ~new_n54289_;
  assign new_n54551_ = ~new_n54549_ & ~new_n54550_;
  assign new_n54552_ = ~new_n54394_ & ~new_n54551_;
  assign new_n54553_ = ~new_n53715_ & ~new_n54393_;
  assign new_n54554_ = ~new_n54392_ & new_n54553_;
  assign new_n54555_ = ~new_n54552_ & ~new_n54554_;
  assign new_n54556_ = ~\b[43]  & ~new_n54555_;
  assign new_n54557_ = ~new_n53734_ & new_n54284_;
  assign new_n54558_ = ~new_n54280_ & new_n54557_;
  assign new_n54559_ = ~new_n54281_ & ~new_n54284_;
  assign new_n54560_ = ~new_n54558_ & ~new_n54559_;
  assign new_n54561_ = ~new_n54394_ & ~new_n54560_;
  assign new_n54562_ = ~new_n53724_ & ~new_n54393_;
  assign new_n54563_ = ~new_n54392_ & new_n54562_;
  assign new_n54564_ = ~new_n54561_ & ~new_n54563_;
  assign new_n54565_ = ~\b[42]  & ~new_n54564_;
  assign new_n54566_ = ~new_n53743_ & new_n54279_;
  assign new_n54567_ = ~new_n54275_ & new_n54566_;
  assign new_n54568_ = ~new_n54276_ & ~new_n54279_;
  assign new_n54569_ = ~new_n54567_ & ~new_n54568_;
  assign new_n54570_ = ~new_n54394_ & ~new_n54569_;
  assign new_n54571_ = ~new_n53733_ & ~new_n54393_;
  assign new_n54572_ = ~new_n54392_ & new_n54571_;
  assign new_n54573_ = ~new_n54570_ & ~new_n54572_;
  assign new_n54574_ = ~\b[41]  & ~new_n54573_;
  assign new_n54575_ = ~new_n53752_ & new_n54274_;
  assign new_n54576_ = ~new_n54270_ & new_n54575_;
  assign new_n54577_ = ~new_n54271_ & ~new_n54274_;
  assign new_n54578_ = ~new_n54576_ & ~new_n54577_;
  assign new_n54579_ = ~new_n54394_ & ~new_n54578_;
  assign new_n54580_ = ~new_n53742_ & ~new_n54393_;
  assign new_n54581_ = ~new_n54392_ & new_n54580_;
  assign new_n54582_ = ~new_n54579_ & ~new_n54581_;
  assign new_n54583_ = ~\b[40]  & ~new_n54582_;
  assign new_n54584_ = ~new_n53761_ & new_n54269_;
  assign new_n54585_ = ~new_n54265_ & new_n54584_;
  assign new_n54586_ = ~new_n54266_ & ~new_n54269_;
  assign new_n54587_ = ~new_n54585_ & ~new_n54586_;
  assign new_n54588_ = ~new_n54394_ & ~new_n54587_;
  assign new_n54589_ = ~new_n53751_ & ~new_n54393_;
  assign new_n54590_ = ~new_n54392_ & new_n54589_;
  assign new_n54591_ = ~new_n54588_ & ~new_n54590_;
  assign new_n54592_ = ~\b[39]  & ~new_n54591_;
  assign new_n54593_ = ~new_n53770_ & new_n54264_;
  assign new_n54594_ = ~new_n54260_ & new_n54593_;
  assign new_n54595_ = ~new_n54261_ & ~new_n54264_;
  assign new_n54596_ = ~new_n54594_ & ~new_n54595_;
  assign new_n54597_ = ~new_n54394_ & ~new_n54596_;
  assign new_n54598_ = ~new_n53760_ & ~new_n54393_;
  assign new_n54599_ = ~new_n54392_ & new_n54598_;
  assign new_n54600_ = ~new_n54597_ & ~new_n54599_;
  assign new_n54601_ = ~\b[38]  & ~new_n54600_;
  assign new_n54602_ = ~new_n53779_ & new_n54259_;
  assign new_n54603_ = ~new_n54255_ & new_n54602_;
  assign new_n54604_ = ~new_n54256_ & ~new_n54259_;
  assign new_n54605_ = ~new_n54603_ & ~new_n54604_;
  assign new_n54606_ = ~new_n54394_ & ~new_n54605_;
  assign new_n54607_ = ~new_n53769_ & ~new_n54393_;
  assign new_n54608_ = ~new_n54392_ & new_n54607_;
  assign new_n54609_ = ~new_n54606_ & ~new_n54608_;
  assign new_n54610_ = ~\b[37]  & ~new_n54609_;
  assign new_n54611_ = ~new_n53788_ & new_n54254_;
  assign new_n54612_ = ~new_n54250_ & new_n54611_;
  assign new_n54613_ = ~new_n54251_ & ~new_n54254_;
  assign new_n54614_ = ~new_n54612_ & ~new_n54613_;
  assign new_n54615_ = ~new_n54394_ & ~new_n54614_;
  assign new_n54616_ = ~new_n53778_ & ~new_n54393_;
  assign new_n54617_ = ~new_n54392_ & new_n54616_;
  assign new_n54618_ = ~new_n54615_ & ~new_n54617_;
  assign new_n54619_ = ~\b[36]  & ~new_n54618_;
  assign new_n54620_ = ~new_n53797_ & new_n54249_;
  assign new_n54621_ = ~new_n54245_ & new_n54620_;
  assign new_n54622_ = ~new_n54246_ & ~new_n54249_;
  assign new_n54623_ = ~new_n54621_ & ~new_n54622_;
  assign new_n54624_ = ~new_n54394_ & ~new_n54623_;
  assign new_n54625_ = ~new_n53787_ & ~new_n54393_;
  assign new_n54626_ = ~new_n54392_ & new_n54625_;
  assign new_n54627_ = ~new_n54624_ & ~new_n54626_;
  assign new_n54628_ = ~\b[35]  & ~new_n54627_;
  assign new_n54629_ = ~new_n53806_ & new_n54244_;
  assign new_n54630_ = ~new_n54240_ & new_n54629_;
  assign new_n54631_ = ~new_n54241_ & ~new_n54244_;
  assign new_n54632_ = ~new_n54630_ & ~new_n54631_;
  assign new_n54633_ = ~new_n54394_ & ~new_n54632_;
  assign new_n54634_ = ~new_n53796_ & ~new_n54393_;
  assign new_n54635_ = ~new_n54392_ & new_n54634_;
  assign new_n54636_ = ~new_n54633_ & ~new_n54635_;
  assign new_n54637_ = ~\b[34]  & ~new_n54636_;
  assign new_n54638_ = ~new_n53815_ & new_n54239_;
  assign new_n54639_ = ~new_n54235_ & new_n54638_;
  assign new_n54640_ = ~new_n54236_ & ~new_n54239_;
  assign new_n54641_ = ~new_n54639_ & ~new_n54640_;
  assign new_n54642_ = ~new_n54394_ & ~new_n54641_;
  assign new_n54643_ = ~new_n53805_ & ~new_n54393_;
  assign new_n54644_ = ~new_n54392_ & new_n54643_;
  assign new_n54645_ = ~new_n54642_ & ~new_n54644_;
  assign new_n54646_ = ~\b[33]  & ~new_n54645_;
  assign new_n54647_ = ~new_n53824_ & new_n54234_;
  assign new_n54648_ = ~new_n54230_ & new_n54647_;
  assign new_n54649_ = ~new_n54231_ & ~new_n54234_;
  assign new_n54650_ = ~new_n54648_ & ~new_n54649_;
  assign new_n54651_ = ~new_n54394_ & ~new_n54650_;
  assign new_n54652_ = ~new_n53814_ & ~new_n54393_;
  assign new_n54653_ = ~new_n54392_ & new_n54652_;
  assign new_n54654_ = ~new_n54651_ & ~new_n54653_;
  assign new_n54655_ = ~\b[32]  & ~new_n54654_;
  assign new_n54656_ = ~new_n53833_ & new_n54229_;
  assign new_n54657_ = ~new_n54225_ & new_n54656_;
  assign new_n54658_ = ~new_n54226_ & ~new_n54229_;
  assign new_n54659_ = ~new_n54657_ & ~new_n54658_;
  assign new_n54660_ = ~new_n54394_ & ~new_n54659_;
  assign new_n54661_ = ~new_n53823_ & ~new_n54393_;
  assign new_n54662_ = ~new_n54392_ & new_n54661_;
  assign new_n54663_ = ~new_n54660_ & ~new_n54662_;
  assign new_n54664_ = ~\b[31]  & ~new_n54663_;
  assign new_n54665_ = ~new_n53842_ & new_n54224_;
  assign new_n54666_ = ~new_n54220_ & new_n54665_;
  assign new_n54667_ = ~new_n54221_ & ~new_n54224_;
  assign new_n54668_ = ~new_n54666_ & ~new_n54667_;
  assign new_n54669_ = ~new_n54394_ & ~new_n54668_;
  assign new_n54670_ = ~new_n53832_ & ~new_n54393_;
  assign new_n54671_ = ~new_n54392_ & new_n54670_;
  assign new_n54672_ = ~new_n54669_ & ~new_n54671_;
  assign new_n54673_ = ~\b[30]  & ~new_n54672_;
  assign new_n54674_ = ~new_n53851_ & new_n54219_;
  assign new_n54675_ = ~new_n54215_ & new_n54674_;
  assign new_n54676_ = ~new_n54216_ & ~new_n54219_;
  assign new_n54677_ = ~new_n54675_ & ~new_n54676_;
  assign new_n54678_ = ~new_n54394_ & ~new_n54677_;
  assign new_n54679_ = ~new_n53841_ & ~new_n54393_;
  assign new_n54680_ = ~new_n54392_ & new_n54679_;
  assign new_n54681_ = ~new_n54678_ & ~new_n54680_;
  assign new_n54682_ = ~\b[29]  & ~new_n54681_;
  assign new_n54683_ = ~new_n53860_ & new_n54214_;
  assign new_n54684_ = ~new_n54210_ & new_n54683_;
  assign new_n54685_ = ~new_n54211_ & ~new_n54214_;
  assign new_n54686_ = ~new_n54684_ & ~new_n54685_;
  assign new_n54687_ = ~new_n54394_ & ~new_n54686_;
  assign new_n54688_ = ~new_n53850_ & ~new_n54393_;
  assign new_n54689_ = ~new_n54392_ & new_n54688_;
  assign new_n54690_ = ~new_n54687_ & ~new_n54689_;
  assign new_n54691_ = ~\b[28]  & ~new_n54690_;
  assign new_n54692_ = ~new_n53869_ & new_n54209_;
  assign new_n54693_ = ~new_n54205_ & new_n54692_;
  assign new_n54694_ = ~new_n54206_ & ~new_n54209_;
  assign new_n54695_ = ~new_n54693_ & ~new_n54694_;
  assign new_n54696_ = ~new_n54394_ & ~new_n54695_;
  assign new_n54697_ = ~new_n53859_ & ~new_n54393_;
  assign new_n54698_ = ~new_n54392_ & new_n54697_;
  assign new_n54699_ = ~new_n54696_ & ~new_n54698_;
  assign new_n54700_ = ~\b[27]  & ~new_n54699_;
  assign new_n54701_ = ~new_n53878_ & new_n54204_;
  assign new_n54702_ = ~new_n54200_ & new_n54701_;
  assign new_n54703_ = ~new_n54201_ & ~new_n54204_;
  assign new_n54704_ = ~new_n54702_ & ~new_n54703_;
  assign new_n54705_ = ~new_n54394_ & ~new_n54704_;
  assign new_n54706_ = ~new_n53868_ & ~new_n54393_;
  assign new_n54707_ = ~new_n54392_ & new_n54706_;
  assign new_n54708_ = ~new_n54705_ & ~new_n54707_;
  assign new_n54709_ = ~\b[26]  & ~new_n54708_;
  assign new_n54710_ = ~new_n53887_ & new_n54199_;
  assign new_n54711_ = ~new_n54195_ & new_n54710_;
  assign new_n54712_ = ~new_n54196_ & ~new_n54199_;
  assign new_n54713_ = ~new_n54711_ & ~new_n54712_;
  assign new_n54714_ = ~new_n54394_ & ~new_n54713_;
  assign new_n54715_ = ~new_n53877_ & ~new_n54393_;
  assign new_n54716_ = ~new_n54392_ & new_n54715_;
  assign new_n54717_ = ~new_n54714_ & ~new_n54716_;
  assign new_n54718_ = ~\b[25]  & ~new_n54717_;
  assign new_n54719_ = ~new_n53896_ & new_n54194_;
  assign new_n54720_ = ~new_n54190_ & new_n54719_;
  assign new_n54721_ = ~new_n54191_ & ~new_n54194_;
  assign new_n54722_ = ~new_n54720_ & ~new_n54721_;
  assign new_n54723_ = ~new_n54394_ & ~new_n54722_;
  assign new_n54724_ = ~new_n53886_ & ~new_n54393_;
  assign new_n54725_ = ~new_n54392_ & new_n54724_;
  assign new_n54726_ = ~new_n54723_ & ~new_n54725_;
  assign new_n54727_ = ~\b[24]  & ~new_n54726_;
  assign new_n54728_ = ~new_n53905_ & new_n54189_;
  assign new_n54729_ = ~new_n54185_ & new_n54728_;
  assign new_n54730_ = ~new_n54186_ & ~new_n54189_;
  assign new_n54731_ = ~new_n54729_ & ~new_n54730_;
  assign new_n54732_ = ~new_n54394_ & ~new_n54731_;
  assign new_n54733_ = ~new_n53895_ & ~new_n54393_;
  assign new_n54734_ = ~new_n54392_ & new_n54733_;
  assign new_n54735_ = ~new_n54732_ & ~new_n54734_;
  assign new_n54736_ = ~\b[23]  & ~new_n54735_;
  assign new_n54737_ = ~new_n53914_ & new_n54184_;
  assign new_n54738_ = ~new_n54180_ & new_n54737_;
  assign new_n54739_ = ~new_n54181_ & ~new_n54184_;
  assign new_n54740_ = ~new_n54738_ & ~new_n54739_;
  assign new_n54741_ = ~new_n54394_ & ~new_n54740_;
  assign new_n54742_ = ~new_n53904_ & ~new_n54393_;
  assign new_n54743_ = ~new_n54392_ & new_n54742_;
  assign new_n54744_ = ~new_n54741_ & ~new_n54743_;
  assign new_n54745_ = ~\b[22]  & ~new_n54744_;
  assign new_n54746_ = ~new_n53923_ & new_n54179_;
  assign new_n54747_ = ~new_n54175_ & new_n54746_;
  assign new_n54748_ = ~new_n54176_ & ~new_n54179_;
  assign new_n54749_ = ~new_n54747_ & ~new_n54748_;
  assign new_n54750_ = ~new_n54394_ & ~new_n54749_;
  assign new_n54751_ = ~new_n53913_ & ~new_n54393_;
  assign new_n54752_ = ~new_n54392_ & new_n54751_;
  assign new_n54753_ = ~new_n54750_ & ~new_n54752_;
  assign new_n54754_ = ~\b[21]  & ~new_n54753_;
  assign new_n54755_ = ~new_n53932_ & new_n54174_;
  assign new_n54756_ = ~new_n54170_ & new_n54755_;
  assign new_n54757_ = ~new_n54171_ & ~new_n54174_;
  assign new_n54758_ = ~new_n54756_ & ~new_n54757_;
  assign new_n54759_ = ~new_n54394_ & ~new_n54758_;
  assign new_n54760_ = ~new_n53922_ & ~new_n54393_;
  assign new_n54761_ = ~new_n54392_ & new_n54760_;
  assign new_n54762_ = ~new_n54759_ & ~new_n54761_;
  assign new_n54763_ = ~\b[20]  & ~new_n54762_;
  assign new_n54764_ = ~new_n53941_ & new_n54169_;
  assign new_n54765_ = ~new_n54165_ & new_n54764_;
  assign new_n54766_ = ~new_n54166_ & ~new_n54169_;
  assign new_n54767_ = ~new_n54765_ & ~new_n54766_;
  assign new_n54768_ = ~new_n54394_ & ~new_n54767_;
  assign new_n54769_ = ~new_n53931_ & ~new_n54393_;
  assign new_n54770_ = ~new_n54392_ & new_n54769_;
  assign new_n54771_ = ~new_n54768_ & ~new_n54770_;
  assign new_n54772_ = ~\b[19]  & ~new_n54771_;
  assign new_n54773_ = ~new_n53950_ & new_n54164_;
  assign new_n54774_ = ~new_n54160_ & new_n54773_;
  assign new_n54775_ = ~new_n54161_ & ~new_n54164_;
  assign new_n54776_ = ~new_n54774_ & ~new_n54775_;
  assign new_n54777_ = ~new_n54394_ & ~new_n54776_;
  assign new_n54778_ = ~new_n53940_ & ~new_n54393_;
  assign new_n54779_ = ~new_n54392_ & new_n54778_;
  assign new_n54780_ = ~new_n54777_ & ~new_n54779_;
  assign new_n54781_ = ~\b[18]  & ~new_n54780_;
  assign new_n54782_ = ~new_n53959_ & new_n54159_;
  assign new_n54783_ = ~new_n54155_ & new_n54782_;
  assign new_n54784_ = ~new_n54156_ & ~new_n54159_;
  assign new_n54785_ = ~new_n54783_ & ~new_n54784_;
  assign new_n54786_ = ~new_n54394_ & ~new_n54785_;
  assign new_n54787_ = ~new_n53949_ & ~new_n54393_;
  assign new_n54788_ = ~new_n54392_ & new_n54787_;
  assign new_n54789_ = ~new_n54786_ & ~new_n54788_;
  assign new_n54790_ = ~\b[17]  & ~new_n54789_;
  assign new_n54791_ = ~new_n53968_ & new_n54154_;
  assign new_n54792_ = ~new_n54150_ & new_n54791_;
  assign new_n54793_ = ~new_n54151_ & ~new_n54154_;
  assign new_n54794_ = ~new_n54792_ & ~new_n54793_;
  assign new_n54795_ = ~new_n54394_ & ~new_n54794_;
  assign new_n54796_ = ~new_n53958_ & ~new_n54393_;
  assign new_n54797_ = ~new_n54392_ & new_n54796_;
  assign new_n54798_ = ~new_n54795_ & ~new_n54797_;
  assign new_n54799_ = ~\b[16]  & ~new_n54798_;
  assign new_n54800_ = ~new_n53977_ & new_n54149_;
  assign new_n54801_ = ~new_n54145_ & new_n54800_;
  assign new_n54802_ = ~new_n54146_ & ~new_n54149_;
  assign new_n54803_ = ~new_n54801_ & ~new_n54802_;
  assign new_n54804_ = ~new_n54394_ & ~new_n54803_;
  assign new_n54805_ = ~new_n53967_ & ~new_n54393_;
  assign new_n54806_ = ~new_n54392_ & new_n54805_;
  assign new_n54807_ = ~new_n54804_ & ~new_n54806_;
  assign new_n54808_ = ~\b[15]  & ~new_n54807_;
  assign new_n54809_ = ~new_n53986_ & new_n54144_;
  assign new_n54810_ = ~new_n54140_ & new_n54809_;
  assign new_n54811_ = ~new_n54141_ & ~new_n54144_;
  assign new_n54812_ = ~new_n54810_ & ~new_n54811_;
  assign new_n54813_ = ~new_n54394_ & ~new_n54812_;
  assign new_n54814_ = ~new_n53976_ & ~new_n54393_;
  assign new_n54815_ = ~new_n54392_ & new_n54814_;
  assign new_n54816_ = ~new_n54813_ & ~new_n54815_;
  assign new_n54817_ = ~\b[14]  & ~new_n54816_;
  assign new_n54818_ = ~new_n53995_ & new_n54139_;
  assign new_n54819_ = ~new_n54135_ & new_n54818_;
  assign new_n54820_ = ~new_n54136_ & ~new_n54139_;
  assign new_n54821_ = ~new_n54819_ & ~new_n54820_;
  assign new_n54822_ = ~new_n54394_ & ~new_n54821_;
  assign new_n54823_ = ~new_n53985_ & ~new_n54393_;
  assign new_n54824_ = ~new_n54392_ & new_n54823_;
  assign new_n54825_ = ~new_n54822_ & ~new_n54824_;
  assign new_n54826_ = ~\b[13]  & ~new_n54825_;
  assign new_n54827_ = ~new_n54004_ & new_n54134_;
  assign new_n54828_ = ~new_n54130_ & new_n54827_;
  assign new_n54829_ = ~new_n54131_ & ~new_n54134_;
  assign new_n54830_ = ~new_n54828_ & ~new_n54829_;
  assign new_n54831_ = ~new_n54394_ & ~new_n54830_;
  assign new_n54832_ = ~new_n53994_ & ~new_n54393_;
  assign new_n54833_ = ~new_n54392_ & new_n54832_;
  assign new_n54834_ = ~new_n54831_ & ~new_n54833_;
  assign new_n54835_ = ~\b[12]  & ~new_n54834_;
  assign new_n54836_ = ~new_n54013_ & new_n54129_;
  assign new_n54837_ = ~new_n54125_ & new_n54836_;
  assign new_n54838_ = ~new_n54126_ & ~new_n54129_;
  assign new_n54839_ = ~new_n54837_ & ~new_n54838_;
  assign new_n54840_ = ~new_n54394_ & ~new_n54839_;
  assign new_n54841_ = ~new_n54003_ & ~new_n54393_;
  assign new_n54842_ = ~new_n54392_ & new_n54841_;
  assign new_n54843_ = ~new_n54840_ & ~new_n54842_;
  assign new_n54844_ = ~\b[11]  & ~new_n54843_;
  assign new_n54845_ = ~new_n54022_ & new_n54124_;
  assign new_n54846_ = ~new_n54120_ & new_n54845_;
  assign new_n54847_ = ~new_n54121_ & ~new_n54124_;
  assign new_n54848_ = ~new_n54846_ & ~new_n54847_;
  assign new_n54849_ = ~new_n54394_ & ~new_n54848_;
  assign new_n54850_ = ~new_n54012_ & ~new_n54393_;
  assign new_n54851_ = ~new_n54392_ & new_n54850_;
  assign new_n54852_ = ~new_n54849_ & ~new_n54851_;
  assign new_n54853_ = ~\b[10]  & ~new_n54852_;
  assign new_n54854_ = ~new_n54031_ & new_n54119_;
  assign new_n54855_ = ~new_n54115_ & new_n54854_;
  assign new_n54856_ = ~new_n54116_ & ~new_n54119_;
  assign new_n54857_ = ~new_n54855_ & ~new_n54856_;
  assign new_n54858_ = ~new_n54394_ & ~new_n54857_;
  assign new_n54859_ = ~new_n54021_ & ~new_n54393_;
  assign new_n54860_ = ~new_n54392_ & new_n54859_;
  assign new_n54861_ = ~new_n54858_ & ~new_n54860_;
  assign new_n54862_ = ~\b[9]  & ~new_n54861_;
  assign new_n54863_ = ~new_n54040_ & new_n54114_;
  assign new_n54864_ = ~new_n54110_ & new_n54863_;
  assign new_n54865_ = ~new_n54111_ & ~new_n54114_;
  assign new_n54866_ = ~new_n54864_ & ~new_n54865_;
  assign new_n54867_ = ~new_n54394_ & ~new_n54866_;
  assign new_n54868_ = ~new_n54030_ & ~new_n54393_;
  assign new_n54869_ = ~new_n54392_ & new_n54868_;
  assign new_n54870_ = ~new_n54867_ & ~new_n54869_;
  assign new_n54871_ = ~\b[8]  & ~new_n54870_;
  assign new_n54872_ = ~new_n54049_ & new_n54109_;
  assign new_n54873_ = ~new_n54105_ & new_n54872_;
  assign new_n54874_ = ~new_n54106_ & ~new_n54109_;
  assign new_n54875_ = ~new_n54873_ & ~new_n54874_;
  assign new_n54876_ = ~new_n54394_ & ~new_n54875_;
  assign new_n54877_ = ~new_n54039_ & ~new_n54393_;
  assign new_n54878_ = ~new_n54392_ & new_n54877_;
  assign new_n54879_ = ~new_n54876_ & ~new_n54878_;
  assign new_n54880_ = ~\b[7]  & ~new_n54879_;
  assign new_n54881_ = ~new_n54058_ & new_n54104_;
  assign new_n54882_ = ~new_n54100_ & new_n54881_;
  assign new_n54883_ = ~new_n54101_ & ~new_n54104_;
  assign new_n54884_ = ~new_n54882_ & ~new_n54883_;
  assign new_n54885_ = ~new_n54394_ & ~new_n54884_;
  assign new_n54886_ = ~new_n54048_ & ~new_n54393_;
  assign new_n54887_ = ~new_n54392_ & new_n54886_;
  assign new_n54888_ = ~new_n54885_ & ~new_n54887_;
  assign new_n54889_ = ~\b[6]  & ~new_n54888_;
  assign new_n54890_ = ~new_n54067_ & new_n54099_;
  assign new_n54891_ = ~new_n54095_ & new_n54890_;
  assign new_n54892_ = ~new_n54096_ & ~new_n54099_;
  assign new_n54893_ = ~new_n54891_ & ~new_n54892_;
  assign new_n54894_ = ~new_n54394_ & ~new_n54893_;
  assign new_n54895_ = ~new_n54057_ & ~new_n54393_;
  assign new_n54896_ = ~new_n54392_ & new_n54895_;
  assign new_n54897_ = ~new_n54894_ & ~new_n54896_;
  assign new_n54898_ = ~\b[5]  & ~new_n54897_;
  assign new_n54899_ = ~new_n54075_ & new_n54094_;
  assign new_n54900_ = ~new_n54090_ & new_n54899_;
  assign new_n54901_ = ~new_n54091_ & ~new_n54094_;
  assign new_n54902_ = ~new_n54900_ & ~new_n54901_;
  assign new_n54903_ = ~new_n54394_ & ~new_n54902_;
  assign new_n54904_ = ~new_n54066_ & ~new_n54393_;
  assign new_n54905_ = ~new_n54392_ & new_n54904_;
  assign new_n54906_ = ~new_n54903_ & ~new_n54905_;
  assign new_n54907_ = ~\b[4]  & ~new_n54906_;
  assign new_n54908_ = ~new_n54085_ & new_n54089_;
  assign new_n54909_ = ~new_n54084_ & new_n54908_;
  assign new_n54910_ = ~new_n54086_ & ~new_n54089_;
  assign new_n54911_ = ~new_n54909_ & ~new_n54910_;
  assign new_n54912_ = ~new_n54394_ & ~new_n54911_;
  assign new_n54913_ = ~new_n54074_ & ~new_n54393_;
  assign new_n54914_ = ~new_n54392_ & new_n54913_;
  assign new_n54915_ = ~new_n54912_ & ~new_n54914_;
  assign new_n54916_ = ~\b[3]  & ~new_n54915_;
  assign new_n54917_ = new_n26069_ & ~new_n54082_;
  assign new_n54918_ = ~new_n54080_ & new_n54917_;
  assign new_n54919_ = ~new_n54084_ & ~new_n54918_;
  assign new_n54920_ = ~new_n54394_ & new_n54919_;
  assign new_n54921_ = ~new_n54079_ & ~new_n54393_;
  assign new_n54922_ = ~new_n54392_ & new_n54921_;
  assign new_n54923_ = ~new_n54920_ & ~new_n54922_;
  assign new_n54924_ = ~\b[2]  & ~new_n54923_;
  assign new_n54925_ = \b[0]  & ~new_n54394_;
  assign new_n54926_ = \a[3]  & ~new_n54925_;
  assign new_n54927_ = new_n26069_ & ~new_n54394_;
  assign new_n54928_ = ~new_n54926_ & ~new_n54927_;
  assign new_n54929_ = \b[1]  & ~new_n54928_;
  assign new_n54930_ = ~\b[1]  & ~new_n54927_;
  assign new_n54931_ = ~new_n54926_ & new_n54930_;
  assign new_n54932_ = ~new_n54929_ & ~new_n54931_;
  assign new_n54933_ = ~new_n26919_ & ~new_n54932_;
  assign new_n54934_ = ~\b[1]  & ~new_n54928_;
  assign new_n54935_ = ~new_n54933_ & ~new_n54934_;
  assign new_n54936_ = \b[2]  & ~new_n54922_;
  assign new_n54937_ = ~new_n54920_ & new_n54936_;
  assign new_n54938_ = ~new_n54924_ & ~new_n54937_;
  assign new_n54939_ = ~new_n54935_ & new_n54938_;
  assign new_n54940_ = ~new_n54924_ & ~new_n54939_;
  assign new_n54941_ = \b[3]  & ~new_n54914_;
  assign new_n54942_ = ~new_n54912_ & new_n54941_;
  assign new_n54943_ = ~new_n54916_ & ~new_n54942_;
  assign new_n54944_ = ~new_n54940_ & new_n54943_;
  assign new_n54945_ = ~new_n54916_ & ~new_n54944_;
  assign new_n54946_ = \b[4]  & ~new_n54905_;
  assign new_n54947_ = ~new_n54903_ & new_n54946_;
  assign new_n54948_ = ~new_n54907_ & ~new_n54947_;
  assign new_n54949_ = ~new_n54945_ & new_n54948_;
  assign new_n54950_ = ~new_n54907_ & ~new_n54949_;
  assign new_n54951_ = \b[5]  & ~new_n54896_;
  assign new_n54952_ = ~new_n54894_ & new_n54951_;
  assign new_n54953_ = ~new_n54898_ & ~new_n54952_;
  assign new_n54954_ = ~new_n54950_ & new_n54953_;
  assign new_n54955_ = ~new_n54898_ & ~new_n54954_;
  assign new_n54956_ = \b[6]  & ~new_n54887_;
  assign new_n54957_ = ~new_n54885_ & new_n54956_;
  assign new_n54958_ = ~new_n54889_ & ~new_n54957_;
  assign new_n54959_ = ~new_n54955_ & new_n54958_;
  assign new_n54960_ = ~new_n54889_ & ~new_n54959_;
  assign new_n54961_ = \b[7]  & ~new_n54878_;
  assign new_n54962_ = ~new_n54876_ & new_n54961_;
  assign new_n54963_ = ~new_n54880_ & ~new_n54962_;
  assign new_n54964_ = ~new_n54960_ & new_n54963_;
  assign new_n54965_ = ~new_n54880_ & ~new_n54964_;
  assign new_n54966_ = \b[8]  & ~new_n54869_;
  assign new_n54967_ = ~new_n54867_ & new_n54966_;
  assign new_n54968_ = ~new_n54871_ & ~new_n54967_;
  assign new_n54969_ = ~new_n54965_ & new_n54968_;
  assign new_n54970_ = ~new_n54871_ & ~new_n54969_;
  assign new_n54971_ = \b[9]  & ~new_n54860_;
  assign new_n54972_ = ~new_n54858_ & new_n54971_;
  assign new_n54973_ = ~new_n54862_ & ~new_n54972_;
  assign new_n54974_ = ~new_n54970_ & new_n54973_;
  assign new_n54975_ = ~new_n54862_ & ~new_n54974_;
  assign new_n54976_ = \b[10]  & ~new_n54851_;
  assign new_n54977_ = ~new_n54849_ & new_n54976_;
  assign new_n54978_ = ~new_n54853_ & ~new_n54977_;
  assign new_n54979_ = ~new_n54975_ & new_n54978_;
  assign new_n54980_ = ~new_n54853_ & ~new_n54979_;
  assign new_n54981_ = \b[11]  & ~new_n54842_;
  assign new_n54982_ = ~new_n54840_ & new_n54981_;
  assign new_n54983_ = ~new_n54844_ & ~new_n54982_;
  assign new_n54984_ = ~new_n54980_ & new_n54983_;
  assign new_n54985_ = ~new_n54844_ & ~new_n54984_;
  assign new_n54986_ = \b[12]  & ~new_n54833_;
  assign new_n54987_ = ~new_n54831_ & new_n54986_;
  assign new_n54988_ = ~new_n54835_ & ~new_n54987_;
  assign new_n54989_ = ~new_n54985_ & new_n54988_;
  assign new_n54990_ = ~new_n54835_ & ~new_n54989_;
  assign new_n54991_ = \b[13]  & ~new_n54824_;
  assign new_n54992_ = ~new_n54822_ & new_n54991_;
  assign new_n54993_ = ~new_n54826_ & ~new_n54992_;
  assign new_n54994_ = ~new_n54990_ & new_n54993_;
  assign new_n54995_ = ~new_n54826_ & ~new_n54994_;
  assign new_n54996_ = \b[14]  & ~new_n54815_;
  assign new_n54997_ = ~new_n54813_ & new_n54996_;
  assign new_n54998_ = ~new_n54817_ & ~new_n54997_;
  assign new_n54999_ = ~new_n54995_ & new_n54998_;
  assign new_n55000_ = ~new_n54817_ & ~new_n54999_;
  assign new_n55001_ = \b[15]  & ~new_n54806_;
  assign new_n55002_ = ~new_n54804_ & new_n55001_;
  assign new_n55003_ = ~new_n54808_ & ~new_n55002_;
  assign new_n55004_ = ~new_n55000_ & new_n55003_;
  assign new_n55005_ = ~new_n54808_ & ~new_n55004_;
  assign new_n55006_ = \b[16]  & ~new_n54797_;
  assign new_n55007_ = ~new_n54795_ & new_n55006_;
  assign new_n55008_ = ~new_n54799_ & ~new_n55007_;
  assign new_n55009_ = ~new_n55005_ & new_n55008_;
  assign new_n55010_ = ~new_n54799_ & ~new_n55009_;
  assign new_n55011_ = \b[17]  & ~new_n54788_;
  assign new_n55012_ = ~new_n54786_ & new_n55011_;
  assign new_n55013_ = ~new_n54790_ & ~new_n55012_;
  assign new_n55014_ = ~new_n55010_ & new_n55013_;
  assign new_n55015_ = ~new_n54790_ & ~new_n55014_;
  assign new_n55016_ = \b[18]  & ~new_n54779_;
  assign new_n55017_ = ~new_n54777_ & new_n55016_;
  assign new_n55018_ = ~new_n54781_ & ~new_n55017_;
  assign new_n55019_ = ~new_n55015_ & new_n55018_;
  assign new_n55020_ = ~new_n54781_ & ~new_n55019_;
  assign new_n55021_ = \b[19]  & ~new_n54770_;
  assign new_n55022_ = ~new_n54768_ & new_n55021_;
  assign new_n55023_ = ~new_n54772_ & ~new_n55022_;
  assign new_n55024_ = ~new_n55020_ & new_n55023_;
  assign new_n55025_ = ~new_n54772_ & ~new_n55024_;
  assign new_n55026_ = \b[20]  & ~new_n54761_;
  assign new_n55027_ = ~new_n54759_ & new_n55026_;
  assign new_n55028_ = ~new_n54763_ & ~new_n55027_;
  assign new_n55029_ = ~new_n55025_ & new_n55028_;
  assign new_n55030_ = ~new_n54763_ & ~new_n55029_;
  assign new_n55031_ = \b[21]  & ~new_n54752_;
  assign new_n55032_ = ~new_n54750_ & new_n55031_;
  assign new_n55033_ = ~new_n54754_ & ~new_n55032_;
  assign new_n55034_ = ~new_n55030_ & new_n55033_;
  assign new_n55035_ = ~new_n54754_ & ~new_n55034_;
  assign new_n55036_ = \b[22]  & ~new_n54743_;
  assign new_n55037_ = ~new_n54741_ & new_n55036_;
  assign new_n55038_ = ~new_n54745_ & ~new_n55037_;
  assign new_n55039_ = ~new_n55035_ & new_n55038_;
  assign new_n55040_ = ~new_n54745_ & ~new_n55039_;
  assign new_n55041_ = \b[23]  & ~new_n54734_;
  assign new_n55042_ = ~new_n54732_ & new_n55041_;
  assign new_n55043_ = ~new_n54736_ & ~new_n55042_;
  assign new_n55044_ = ~new_n55040_ & new_n55043_;
  assign new_n55045_ = ~new_n54736_ & ~new_n55044_;
  assign new_n55046_ = \b[24]  & ~new_n54725_;
  assign new_n55047_ = ~new_n54723_ & new_n55046_;
  assign new_n55048_ = ~new_n54727_ & ~new_n55047_;
  assign new_n55049_ = ~new_n55045_ & new_n55048_;
  assign new_n55050_ = ~new_n54727_ & ~new_n55049_;
  assign new_n55051_ = \b[25]  & ~new_n54716_;
  assign new_n55052_ = ~new_n54714_ & new_n55051_;
  assign new_n55053_ = ~new_n54718_ & ~new_n55052_;
  assign new_n55054_ = ~new_n55050_ & new_n55053_;
  assign new_n55055_ = ~new_n54718_ & ~new_n55054_;
  assign new_n55056_ = \b[26]  & ~new_n54707_;
  assign new_n55057_ = ~new_n54705_ & new_n55056_;
  assign new_n55058_ = ~new_n54709_ & ~new_n55057_;
  assign new_n55059_ = ~new_n55055_ & new_n55058_;
  assign new_n55060_ = ~new_n54709_ & ~new_n55059_;
  assign new_n55061_ = \b[27]  & ~new_n54698_;
  assign new_n55062_ = ~new_n54696_ & new_n55061_;
  assign new_n55063_ = ~new_n54700_ & ~new_n55062_;
  assign new_n55064_ = ~new_n55060_ & new_n55063_;
  assign new_n55065_ = ~new_n54700_ & ~new_n55064_;
  assign new_n55066_ = \b[28]  & ~new_n54689_;
  assign new_n55067_ = ~new_n54687_ & new_n55066_;
  assign new_n55068_ = ~new_n54691_ & ~new_n55067_;
  assign new_n55069_ = ~new_n55065_ & new_n55068_;
  assign new_n55070_ = ~new_n54691_ & ~new_n55069_;
  assign new_n55071_ = \b[29]  & ~new_n54680_;
  assign new_n55072_ = ~new_n54678_ & new_n55071_;
  assign new_n55073_ = ~new_n54682_ & ~new_n55072_;
  assign new_n55074_ = ~new_n55070_ & new_n55073_;
  assign new_n55075_ = ~new_n54682_ & ~new_n55074_;
  assign new_n55076_ = \b[30]  & ~new_n54671_;
  assign new_n55077_ = ~new_n54669_ & new_n55076_;
  assign new_n55078_ = ~new_n54673_ & ~new_n55077_;
  assign new_n55079_ = ~new_n55075_ & new_n55078_;
  assign new_n55080_ = ~new_n54673_ & ~new_n55079_;
  assign new_n55081_ = \b[31]  & ~new_n54662_;
  assign new_n55082_ = ~new_n54660_ & new_n55081_;
  assign new_n55083_ = ~new_n54664_ & ~new_n55082_;
  assign new_n55084_ = ~new_n55080_ & new_n55083_;
  assign new_n55085_ = ~new_n54664_ & ~new_n55084_;
  assign new_n55086_ = \b[32]  & ~new_n54653_;
  assign new_n55087_ = ~new_n54651_ & new_n55086_;
  assign new_n55088_ = ~new_n54655_ & ~new_n55087_;
  assign new_n55089_ = ~new_n55085_ & new_n55088_;
  assign new_n55090_ = ~new_n54655_ & ~new_n55089_;
  assign new_n55091_ = \b[33]  & ~new_n54644_;
  assign new_n55092_ = ~new_n54642_ & new_n55091_;
  assign new_n55093_ = ~new_n54646_ & ~new_n55092_;
  assign new_n55094_ = ~new_n55090_ & new_n55093_;
  assign new_n55095_ = ~new_n54646_ & ~new_n55094_;
  assign new_n55096_ = \b[34]  & ~new_n54635_;
  assign new_n55097_ = ~new_n54633_ & new_n55096_;
  assign new_n55098_ = ~new_n54637_ & ~new_n55097_;
  assign new_n55099_ = ~new_n55095_ & new_n55098_;
  assign new_n55100_ = ~new_n54637_ & ~new_n55099_;
  assign new_n55101_ = \b[35]  & ~new_n54626_;
  assign new_n55102_ = ~new_n54624_ & new_n55101_;
  assign new_n55103_ = ~new_n54628_ & ~new_n55102_;
  assign new_n55104_ = ~new_n55100_ & new_n55103_;
  assign new_n55105_ = ~new_n54628_ & ~new_n55104_;
  assign new_n55106_ = \b[36]  & ~new_n54617_;
  assign new_n55107_ = ~new_n54615_ & new_n55106_;
  assign new_n55108_ = ~new_n54619_ & ~new_n55107_;
  assign new_n55109_ = ~new_n55105_ & new_n55108_;
  assign new_n55110_ = ~new_n54619_ & ~new_n55109_;
  assign new_n55111_ = \b[37]  & ~new_n54608_;
  assign new_n55112_ = ~new_n54606_ & new_n55111_;
  assign new_n55113_ = ~new_n54610_ & ~new_n55112_;
  assign new_n55114_ = ~new_n55110_ & new_n55113_;
  assign new_n55115_ = ~new_n54610_ & ~new_n55114_;
  assign new_n55116_ = \b[38]  & ~new_n54599_;
  assign new_n55117_ = ~new_n54597_ & new_n55116_;
  assign new_n55118_ = ~new_n54601_ & ~new_n55117_;
  assign new_n55119_ = ~new_n55115_ & new_n55118_;
  assign new_n55120_ = ~new_n54601_ & ~new_n55119_;
  assign new_n55121_ = \b[39]  & ~new_n54590_;
  assign new_n55122_ = ~new_n54588_ & new_n55121_;
  assign new_n55123_ = ~new_n54592_ & ~new_n55122_;
  assign new_n55124_ = ~new_n55120_ & new_n55123_;
  assign new_n55125_ = ~new_n54592_ & ~new_n55124_;
  assign new_n55126_ = \b[40]  & ~new_n54581_;
  assign new_n55127_ = ~new_n54579_ & new_n55126_;
  assign new_n55128_ = ~new_n54583_ & ~new_n55127_;
  assign new_n55129_ = ~new_n55125_ & new_n55128_;
  assign new_n55130_ = ~new_n54583_ & ~new_n55129_;
  assign new_n55131_ = \b[41]  & ~new_n54572_;
  assign new_n55132_ = ~new_n54570_ & new_n55131_;
  assign new_n55133_ = ~new_n54574_ & ~new_n55132_;
  assign new_n55134_ = ~new_n55130_ & new_n55133_;
  assign new_n55135_ = ~new_n54574_ & ~new_n55134_;
  assign new_n55136_ = \b[42]  & ~new_n54563_;
  assign new_n55137_ = ~new_n54561_ & new_n55136_;
  assign new_n55138_ = ~new_n54565_ & ~new_n55137_;
  assign new_n55139_ = ~new_n55135_ & new_n55138_;
  assign new_n55140_ = ~new_n54565_ & ~new_n55139_;
  assign new_n55141_ = \b[43]  & ~new_n54554_;
  assign new_n55142_ = ~new_n54552_ & new_n55141_;
  assign new_n55143_ = ~new_n54556_ & ~new_n55142_;
  assign new_n55144_ = ~new_n55140_ & new_n55143_;
  assign new_n55145_ = ~new_n54556_ & ~new_n55144_;
  assign new_n55146_ = \b[44]  & ~new_n54545_;
  assign new_n55147_ = ~new_n54543_ & new_n55146_;
  assign new_n55148_ = ~new_n54547_ & ~new_n55147_;
  assign new_n55149_ = ~new_n55145_ & new_n55148_;
  assign new_n55150_ = ~new_n54547_ & ~new_n55149_;
  assign new_n55151_ = \b[45]  & ~new_n54536_;
  assign new_n55152_ = ~new_n54534_ & new_n55151_;
  assign new_n55153_ = ~new_n54538_ & ~new_n55152_;
  assign new_n55154_ = ~new_n55150_ & new_n55153_;
  assign new_n55155_ = ~new_n54538_ & ~new_n55154_;
  assign new_n55156_ = \b[46]  & ~new_n54527_;
  assign new_n55157_ = ~new_n54525_ & new_n55156_;
  assign new_n55158_ = ~new_n54529_ & ~new_n55157_;
  assign new_n55159_ = ~new_n55155_ & new_n55158_;
  assign new_n55160_ = ~new_n54529_ & ~new_n55159_;
  assign new_n55161_ = \b[47]  & ~new_n54518_;
  assign new_n55162_ = ~new_n54516_ & new_n55161_;
  assign new_n55163_ = ~new_n54520_ & ~new_n55162_;
  assign new_n55164_ = ~new_n55160_ & new_n55163_;
  assign new_n55165_ = ~new_n54520_ & ~new_n55164_;
  assign new_n55166_ = \b[48]  & ~new_n54509_;
  assign new_n55167_ = ~new_n54507_ & new_n55166_;
  assign new_n55168_ = ~new_n54511_ & ~new_n55167_;
  assign new_n55169_ = ~new_n55165_ & new_n55168_;
  assign new_n55170_ = ~new_n54511_ & ~new_n55169_;
  assign new_n55171_ = \b[49]  & ~new_n54500_;
  assign new_n55172_ = ~new_n54498_ & new_n55171_;
  assign new_n55173_ = ~new_n54502_ & ~new_n55172_;
  assign new_n55174_ = ~new_n55170_ & new_n55173_;
  assign new_n55175_ = ~new_n54502_ & ~new_n55174_;
  assign new_n55176_ = \b[50]  & ~new_n54491_;
  assign new_n55177_ = ~new_n54489_ & new_n55176_;
  assign new_n55178_ = ~new_n54493_ & ~new_n55177_;
  assign new_n55179_ = ~new_n55175_ & new_n55178_;
  assign new_n55180_ = ~new_n54493_ & ~new_n55179_;
  assign new_n55181_ = \b[51]  & ~new_n54482_;
  assign new_n55182_ = ~new_n54480_ & new_n55181_;
  assign new_n55183_ = ~new_n54484_ & ~new_n55182_;
  assign new_n55184_ = ~new_n55180_ & new_n55183_;
  assign new_n55185_ = ~new_n54484_ & ~new_n55184_;
  assign new_n55186_ = \b[52]  & ~new_n54473_;
  assign new_n55187_ = ~new_n54471_ & new_n55186_;
  assign new_n55188_ = ~new_n54475_ & ~new_n55187_;
  assign new_n55189_ = ~new_n55185_ & new_n55188_;
  assign new_n55190_ = ~new_n54475_ & ~new_n55189_;
  assign new_n55191_ = \b[53]  & ~new_n54464_;
  assign new_n55192_ = ~new_n54462_ & new_n55191_;
  assign new_n55193_ = ~new_n54466_ & ~new_n55192_;
  assign new_n55194_ = ~new_n55190_ & new_n55193_;
  assign new_n55195_ = ~new_n54466_ & ~new_n55194_;
  assign new_n55196_ = \b[54]  & ~new_n54455_;
  assign new_n55197_ = ~new_n54453_ & new_n55196_;
  assign new_n55198_ = ~new_n54457_ & ~new_n55197_;
  assign new_n55199_ = ~new_n55195_ & new_n55198_;
  assign new_n55200_ = ~new_n54457_ & ~new_n55199_;
  assign new_n55201_ = \b[55]  & ~new_n54446_;
  assign new_n55202_ = ~new_n54444_ & new_n55201_;
  assign new_n55203_ = ~new_n54448_ & ~new_n55202_;
  assign new_n55204_ = ~new_n55200_ & new_n55203_;
  assign new_n55205_ = ~new_n54448_ & ~new_n55204_;
  assign new_n55206_ = \b[56]  & ~new_n54437_;
  assign new_n55207_ = ~new_n54435_ & new_n55206_;
  assign new_n55208_ = ~new_n54439_ & ~new_n55207_;
  assign new_n55209_ = ~new_n55205_ & new_n55208_;
  assign new_n55210_ = ~new_n54439_ & ~new_n55209_;
  assign new_n55211_ = \b[57]  & ~new_n54428_;
  assign new_n55212_ = ~new_n54426_ & new_n55211_;
  assign new_n55213_ = ~new_n54430_ & ~new_n55212_;
  assign new_n55214_ = ~new_n55210_ & new_n55213_;
  assign new_n55215_ = ~new_n54430_ & ~new_n55214_;
  assign new_n55216_ = \b[58]  & ~new_n54419_;
  assign new_n55217_ = ~new_n54417_ & new_n55216_;
  assign new_n55218_ = ~new_n54421_ & ~new_n55217_;
  assign new_n55219_ = ~new_n55215_ & new_n55218_;
  assign new_n55220_ = ~new_n54421_ & ~new_n55219_;
  assign new_n55221_ = \b[59]  & ~new_n54410_;
  assign new_n55222_ = ~new_n54408_ & new_n55221_;
  assign new_n55223_ = ~new_n54412_ & ~new_n55222_;
  assign new_n55224_ = ~new_n55220_ & new_n55223_;
  assign new_n55225_ = ~new_n54412_ & ~new_n55224_;
  assign new_n55226_ = \b[60]  & ~new_n54401_;
  assign new_n55227_ = ~new_n54399_ & new_n55226_;
  assign new_n55228_ = ~new_n54403_ & ~new_n55227_;
  assign new_n55229_ = ~new_n55225_ & new_n55228_;
  assign new_n55230_ = ~new_n54403_ & ~new_n55229_;
  assign new_n55231_ = ~new_n53563_ & ~new_n54389_;
  assign new_n55232_ = ~new_n54387_ & new_n55231_;
  assign new_n55233_ = ~new_n54375_ & new_n55232_;
  assign new_n55234_ = ~new_n54387_ & ~new_n54389_;
  assign new_n55235_ = ~new_n54376_ & ~new_n55234_;
  assign new_n55236_ = ~new_n55233_ & ~new_n55235_;
  assign new_n55237_ = ~new_n54394_ & ~new_n55236_;
  assign new_n55238_ = ~new_n54386_ & ~new_n54393_;
  assign new_n55239_ = ~new_n54392_ & new_n55238_;
  assign new_n55240_ = ~new_n55237_ & ~new_n55239_;
  assign new_n55241_ = ~\b[61]  & ~new_n55240_;
  assign new_n55242_ = \b[61]  & ~new_n55239_;
  assign new_n55243_ = ~new_n55237_ & new_n55242_;
  assign new_n55244_ = new_n279_ & ~new_n55243_;
  assign new_n55245_ = ~new_n55241_ & new_n55244_;
  assign new_n55246_ = ~new_n55230_ & new_n55245_;
  assign new_n55247_ = new_n403_ & ~new_n55240_;
  assign new_n55248_ = ~new_n55246_ & ~new_n55247_;
  assign new_n55249_ = ~new_n54412_ & new_n55228_;
  assign new_n55250_ = ~new_n55224_ & new_n55249_;
  assign new_n55251_ = ~new_n55225_ & ~new_n55228_;
  assign new_n55252_ = ~new_n55250_ & ~new_n55251_;
  assign new_n55253_ = ~new_n55248_ & ~new_n55252_;
  assign new_n55254_ = ~new_n54402_ & ~new_n55247_;
  assign new_n55255_ = ~new_n55246_ & new_n55254_;
  assign new_n55256_ = ~new_n55253_ & ~new_n55255_;
  assign new_n55257_ = ~\b[61]  & ~new_n55256_;
  assign new_n55258_ = ~new_n54421_ & new_n55223_;
  assign new_n55259_ = ~new_n55219_ & new_n55258_;
  assign new_n55260_ = ~new_n55220_ & ~new_n55223_;
  assign new_n55261_ = ~new_n55259_ & ~new_n55260_;
  assign new_n55262_ = ~new_n55248_ & ~new_n55261_;
  assign new_n55263_ = ~new_n54411_ & ~new_n55247_;
  assign new_n55264_ = ~new_n55246_ & new_n55263_;
  assign new_n55265_ = ~new_n55262_ & ~new_n55264_;
  assign new_n55266_ = ~\b[60]  & ~new_n55265_;
  assign new_n55267_ = ~new_n54430_ & new_n55218_;
  assign new_n55268_ = ~new_n55214_ & new_n55267_;
  assign new_n55269_ = ~new_n55215_ & ~new_n55218_;
  assign new_n55270_ = ~new_n55268_ & ~new_n55269_;
  assign new_n55271_ = ~new_n55248_ & ~new_n55270_;
  assign new_n55272_ = ~new_n54420_ & ~new_n55247_;
  assign new_n55273_ = ~new_n55246_ & new_n55272_;
  assign new_n55274_ = ~new_n55271_ & ~new_n55273_;
  assign new_n55275_ = ~\b[59]  & ~new_n55274_;
  assign new_n55276_ = ~new_n54439_ & new_n55213_;
  assign new_n55277_ = ~new_n55209_ & new_n55276_;
  assign new_n55278_ = ~new_n55210_ & ~new_n55213_;
  assign new_n55279_ = ~new_n55277_ & ~new_n55278_;
  assign new_n55280_ = ~new_n55248_ & ~new_n55279_;
  assign new_n55281_ = ~new_n54429_ & ~new_n55247_;
  assign new_n55282_ = ~new_n55246_ & new_n55281_;
  assign new_n55283_ = ~new_n55280_ & ~new_n55282_;
  assign new_n55284_ = ~\b[58]  & ~new_n55283_;
  assign new_n55285_ = ~new_n54448_ & new_n55208_;
  assign new_n55286_ = ~new_n55204_ & new_n55285_;
  assign new_n55287_ = ~new_n55205_ & ~new_n55208_;
  assign new_n55288_ = ~new_n55286_ & ~new_n55287_;
  assign new_n55289_ = ~new_n55248_ & ~new_n55288_;
  assign new_n55290_ = ~new_n54438_ & ~new_n55247_;
  assign new_n55291_ = ~new_n55246_ & new_n55290_;
  assign new_n55292_ = ~new_n55289_ & ~new_n55291_;
  assign new_n55293_ = ~\b[57]  & ~new_n55292_;
  assign new_n55294_ = ~new_n54457_ & new_n55203_;
  assign new_n55295_ = ~new_n55199_ & new_n55294_;
  assign new_n55296_ = ~new_n55200_ & ~new_n55203_;
  assign new_n55297_ = ~new_n55295_ & ~new_n55296_;
  assign new_n55298_ = ~new_n55248_ & ~new_n55297_;
  assign new_n55299_ = ~new_n54447_ & ~new_n55247_;
  assign new_n55300_ = ~new_n55246_ & new_n55299_;
  assign new_n55301_ = ~new_n55298_ & ~new_n55300_;
  assign new_n55302_ = ~\b[56]  & ~new_n55301_;
  assign new_n55303_ = ~new_n54466_ & new_n55198_;
  assign new_n55304_ = ~new_n55194_ & new_n55303_;
  assign new_n55305_ = ~new_n55195_ & ~new_n55198_;
  assign new_n55306_ = ~new_n55304_ & ~new_n55305_;
  assign new_n55307_ = ~new_n55248_ & ~new_n55306_;
  assign new_n55308_ = ~new_n54456_ & ~new_n55247_;
  assign new_n55309_ = ~new_n55246_ & new_n55308_;
  assign new_n55310_ = ~new_n55307_ & ~new_n55309_;
  assign new_n55311_ = ~\b[55]  & ~new_n55310_;
  assign new_n55312_ = ~new_n54475_ & new_n55193_;
  assign new_n55313_ = ~new_n55189_ & new_n55312_;
  assign new_n55314_ = ~new_n55190_ & ~new_n55193_;
  assign new_n55315_ = ~new_n55313_ & ~new_n55314_;
  assign new_n55316_ = ~new_n55248_ & ~new_n55315_;
  assign new_n55317_ = ~new_n54465_ & ~new_n55247_;
  assign new_n55318_ = ~new_n55246_ & new_n55317_;
  assign new_n55319_ = ~new_n55316_ & ~new_n55318_;
  assign new_n55320_ = ~\b[54]  & ~new_n55319_;
  assign new_n55321_ = ~new_n54484_ & new_n55188_;
  assign new_n55322_ = ~new_n55184_ & new_n55321_;
  assign new_n55323_ = ~new_n55185_ & ~new_n55188_;
  assign new_n55324_ = ~new_n55322_ & ~new_n55323_;
  assign new_n55325_ = ~new_n55248_ & ~new_n55324_;
  assign new_n55326_ = ~new_n54474_ & ~new_n55247_;
  assign new_n55327_ = ~new_n55246_ & new_n55326_;
  assign new_n55328_ = ~new_n55325_ & ~new_n55327_;
  assign new_n55329_ = ~\b[53]  & ~new_n55328_;
  assign new_n55330_ = ~new_n54493_ & new_n55183_;
  assign new_n55331_ = ~new_n55179_ & new_n55330_;
  assign new_n55332_ = ~new_n55180_ & ~new_n55183_;
  assign new_n55333_ = ~new_n55331_ & ~new_n55332_;
  assign new_n55334_ = ~new_n55248_ & ~new_n55333_;
  assign new_n55335_ = ~new_n54483_ & ~new_n55247_;
  assign new_n55336_ = ~new_n55246_ & new_n55335_;
  assign new_n55337_ = ~new_n55334_ & ~new_n55336_;
  assign new_n55338_ = ~\b[52]  & ~new_n55337_;
  assign new_n55339_ = ~new_n54502_ & new_n55178_;
  assign new_n55340_ = ~new_n55174_ & new_n55339_;
  assign new_n55341_ = ~new_n55175_ & ~new_n55178_;
  assign new_n55342_ = ~new_n55340_ & ~new_n55341_;
  assign new_n55343_ = ~new_n55248_ & ~new_n55342_;
  assign new_n55344_ = ~new_n54492_ & ~new_n55247_;
  assign new_n55345_ = ~new_n55246_ & new_n55344_;
  assign new_n55346_ = ~new_n55343_ & ~new_n55345_;
  assign new_n55347_ = ~\b[51]  & ~new_n55346_;
  assign new_n55348_ = ~new_n54511_ & new_n55173_;
  assign new_n55349_ = ~new_n55169_ & new_n55348_;
  assign new_n55350_ = ~new_n55170_ & ~new_n55173_;
  assign new_n55351_ = ~new_n55349_ & ~new_n55350_;
  assign new_n55352_ = ~new_n55248_ & ~new_n55351_;
  assign new_n55353_ = ~new_n54501_ & ~new_n55247_;
  assign new_n55354_ = ~new_n55246_ & new_n55353_;
  assign new_n55355_ = ~new_n55352_ & ~new_n55354_;
  assign new_n55356_ = ~\b[50]  & ~new_n55355_;
  assign new_n55357_ = ~new_n54520_ & new_n55168_;
  assign new_n55358_ = ~new_n55164_ & new_n55357_;
  assign new_n55359_ = ~new_n55165_ & ~new_n55168_;
  assign new_n55360_ = ~new_n55358_ & ~new_n55359_;
  assign new_n55361_ = ~new_n55248_ & ~new_n55360_;
  assign new_n55362_ = ~new_n54510_ & ~new_n55247_;
  assign new_n55363_ = ~new_n55246_ & new_n55362_;
  assign new_n55364_ = ~new_n55361_ & ~new_n55363_;
  assign new_n55365_ = ~\b[49]  & ~new_n55364_;
  assign new_n55366_ = ~new_n54529_ & new_n55163_;
  assign new_n55367_ = ~new_n55159_ & new_n55366_;
  assign new_n55368_ = ~new_n55160_ & ~new_n55163_;
  assign new_n55369_ = ~new_n55367_ & ~new_n55368_;
  assign new_n55370_ = ~new_n55248_ & ~new_n55369_;
  assign new_n55371_ = ~new_n54519_ & ~new_n55247_;
  assign new_n55372_ = ~new_n55246_ & new_n55371_;
  assign new_n55373_ = ~new_n55370_ & ~new_n55372_;
  assign new_n55374_ = ~\b[48]  & ~new_n55373_;
  assign new_n55375_ = ~new_n54538_ & new_n55158_;
  assign new_n55376_ = ~new_n55154_ & new_n55375_;
  assign new_n55377_ = ~new_n55155_ & ~new_n55158_;
  assign new_n55378_ = ~new_n55376_ & ~new_n55377_;
  assign new_n55379_ = ~new_n55248_ & ~new_n55378_;
  assign new_n55380_ = ~new_n54528_ & ~new_n55247_;
  assign new_n55381_ = ~new_n55246_ & new_n55380_;
  assign new_n55382_ = ~new_n55379_ & ~new_n55381_;
  assign new_n55383_ = ~\b[47]  & ~new_n55382_;
  assign new_n55384_ = ~new_n54547_ & new_n55153_;
  assign new_n55385_ = ~new_n55149_ & new_n55384_;
  assign new_n55386_ = ~new_n55150_ & ~new_n55153_;
  assign new_n55387_ = ~new_n55385_ & ~new_n55386_;
  assign new_n55388_ = ~new_n55248_ & ~new_n55387_;
  assign new_n55389_ = ~new_n54537_ & ~new_n55247_;
  assign new_n55390_ = ~new_n55246_ & new_n55389_;
  assign new_n55391_ = ~new_n55388_ & ~new_n55390_;
  assign new_n55392_ = ~\b[46]  & ~new_n55391_;
  assign new_n55393_ = ~new_n54556_ & new_n55148_;
  assign new_n55394_ = ~new_n55144_ & new_n55393_;
  assign new_n55395_ = ~new_n55145_ & ~new_n55148_;
  assign new_n55396_ = ~new_n55394_ & ~new_n55395_;
  assign new_n55397_ = ~new_n55248_ & ~new_n55396_;
  assign new_n55398_ = ~new_n54546_ & ~new_n55247_;
  assign new_n55399_ = ~new_n55246_ & new_n55398_;
  assign new_n55400_ = ~new_n55397_ & ~new_n55399_;
  assign new_n55401_ = ~\b[45]  & ~new_n55400_;
  assign new_n55402_ = ~new_n54565_ & new_n55143_;
  assign new_n55403_ = ~new_n55139_ & new_n55402_;
  assign new_n55404_ = ~new_n55140_ & ~new_n55143_;
  assign new_n55405_ = ~new_n55403_ & ~new_n55404_;
  assign new_n55406_ = ~new_n55248_ & ~new_n55405_;
  assign new_n55407_ = ~new_n54555_ & ~new_n55247_;
  assign new_n55408_ = ~new_n55246_ & new_n55407_;
  assign new_n55409_ = ~new_n55406_ & ~new_n55408_;
  assign new_n55410_ = ~\b[44]  & ~new_n55409_;
  assign new_n55411_ = ~new_n54574_ & new_n55138_;
  assign new_n55412_ = ~new_n55134_ & new_n55411_;
  assign new_n55413_ = ~new_n55135_ & ~new_n55138_;
  assign new_n55414_ = ~new_n55412_ & ~new_n55413_;
  assign new_n55415_ = ~new_n55248_ & ~new_n55414_;
  assign new_n55416_ = ~new_n54564_ & ~new_n55247_;
  assign new_n55417_ = ~new_n55246_ & new_n55416_;
  assign new_n55418_ = ~new_n55415_ & ~new_n55417_;
  assign new_n55419_ = ~\b[43]  & ~new_n55418_;
  assign new_n55420_ = ~new_n54583_ & new_n55133_;
  assign new_n55421_ = ~new_n55129_ & new_n55420_;
  assign new_n55422_ = ~new_n55130_ & ~new_n55133_;
  assign new_n55423_ = ~new_n55421_ & ~new_n55422_;
  assign new_n55424_ = ~new_n55248_ & ~new_n55423_;
  assign new_n55425_ = ~new_n54573_ & ~new_n55247_;
  assign new_n55426_ = ~new_n55246_ & new_n55425_;
  assign new_n55427_ = ~new_n55424_ & ~new_n55426_;
  assign new_n55428_ = ~\b[42]  & ~new_n55427_;
  assign new_n55429_ = ~new_n54592_ & new_n55128_;
  assign new_n55430_ = ~new_n55124_ & new_n55429_;
  assign new_n55431_ = ~new_n55125_ & ~new_n55128_;
  assign new_n55432_ = ~new_n55430_ & ~new_n55431_;
  assign new_n55433_ = ~new_n55248_ & ~new_n55432_;
  assign new_n55434_ = ~new_n54582_ & ~new_n55247_;
  assign new_n55435_ = ~new_n55246_ & new_n55434_;
  assign new_n55436_ = ~new_n55433_ & ~new_n55435_;
  assign new_n55437_ = ~\b[41]  & ~new_n55436_;
  assign new_n55438_ = ~new_n54601_ & new_n55123_;
  assign new_n55439_ = ~new_n55119_ & new_n55438_;
  assign new_n55440_ = ~new_n55120_ & ~new_n55123_;
  assign new_n55441_ = ~new_n55439_ & ~new_n55440_;
  assign new_n55442_ = ~new_n55248_ & ~new_n55441_;
  assign new_n55443_ = ~new_n54591_ & ~new_n55247_;
  assign new_n55444_ = ~new_n55246_ & new_n55443_;
  assign new_n55445_ = ~new_n55442_ & ~new_n55444_;
  assign new_n55446_ = ~\b[40]  & ~new_n55445_;
  assign new_n55447_ = ~new_n54610_ & new_n55118_;
  assign new_n55448_ = ~new_n55114_ & new_n55447_;
  assign new_n55449_ = ~new_n55115_ & ~new_n55118_;
  assign new_n55450_ = ~new_n55448_ & ~new_n55449_;
  assign new_n55451_ = ~new_n55248_ & ~new_n55450_;
  assign new_n55452_ = ~new_n54600_ & ~new_n55247_;
  assign new_n55453_ = ~new_n55246_ & new_n55452_;
  assign new_n55454_ = ~new_n55451_ & ~new_n55453_;
  assign new_n55455_ = ~\b[39]  & ~new_n55454_;
  assign new_n55456_ = ~new_n54619_ & new_n55113_;
  assign new_n55457_ = ~new_n55109_ & new_n55456_;
  assign new_n55458_ = ~new_n55110_ & ~new_n55113_;
  assign new_n55459_ = ~new_n55457_ & ~new_n55458_;
  assign new_n55460_ = ~new_n55248_ & ~new_n55459_;
  assign new_n55461_ = ~new_n54609_ & ~new_n55247_;
  assign new_n55462_ = ~new_n55246_ & new_n55461_;
  assign new_n55463_ = ~new_n55460_ & ~new_n55462_;
  assign new_n55464_ = ~\b[38]  & ~new_n55463_;
  assign new_n55465_ = ~new_n54628_ & new_n55108_;
  assign new_n55466_ = ~new_n55104_ & new_n55465_;
  assign new_n55467_ = ~new_n55105_ & ~new_n55108_;
  assign new_n55468_ = ~new_n55466_ & ~new_n55467_;
  assign new_n55469_ = ~new_n55248_ & ~new_n55468_;
  assign new_n55470_ = ~new_n54618_ & ~new_n55247_;
  assign new_n55471_ = ~new_n55246_ & new_n55470_;
  assign new_n55472_ = ~new_n55469_ & ~new_n55471_;
  assign new_n55473_ = ~\b[37]  & ~new_n55472_;
  assign new_n55474_ = ~new_n54637_ & new_n55103_;
  assign new_n55475_ = ~new_n55099_ & new_n55474_;
  assign new_n55476_ = ~new_n55100_ & ~new_n55103_;
  assign new_n55477_ = ~new_n55475_ & ~new_n55476_;
  assign new_n55478_ = ~new_n55248_ & ~new_n55477_;
  assign new_n55479_ = ~new_n54627_ & ~new_n55247_;
  assign new_n55480_ = ~new_n55246_ & new_n55479_;
  assign new_n55481_ = ~new_n55478_ & ~new_n55480_;
  assign new_n55482_ = ~\b[36]  & ~new_n55481_;
  assign new_n55483_ = ~new_n54646_ & new_n55098_;
  assign new_n55484_ = ~new_n55094_ & new_n55483_;
  assign new_n55485_ = ~new_n55095_ & ~new_n55098_;
  assign new_n55486_ = ~new_n55484_ & ~new_n55485_;
  assign new_n55487_ = ~new_n55248_ & ~new_n55486_;
  assign new_n55488_ = ~new_n54636_ & ~new_n55247_;
  assign new_n55489_ = ~new_n55246_ & new_n55488_;
  assign new_n55490_ = ~new_n55487_ & ~new_n55489_;
  assign new_n55491_ = ~\b[35]  & ~new_n55490_;
  assign new_n55492_ = ~new_n54655_ & new_n55093_;
  assign new_n55493_ = ~new_n55089_ & new_n55492_;
  assign new_n55494_ = ~new_n55090_ & ~new_n55093_;
  assign new_n55495_ = ~new_n55493_ & ~new_n55494_;
  assign new_n55496_ = ~new_n55248_ & ~new_n55495_;
  assign new_n55497_ = ~new_n54645_ & ~new_n55247_;
  assign new_n55498_ = ~new_n55246_ & new_n55497_;
  assign new_n55499_ = ~new_n55496_ & ~new_n55498_;
  assign new_n55500_ = ~\b[34]  & ~new_n55499_;
  assign new_n55501_ = ~new_n54664_ & new_n55088_;
  assign new_n55502_ = ~new_n55084_ & new_n55501_;
  assign new_n55503_ = ~new_n55085_ & ~new_n55088_;
  assign new_n55504_ = ~new_n55502_ & ~new_n55503_;
  assign new_n55505_ = ~new_n55248_ & ~new_n55504_;
  assign new_n55506_ = ~new_n54654_ & ~new_n55247_;
  assign new_n55507_ = ~new_n55246_ & new_n55506_;
  assign new_n55508_ = ~new_n55505_ & ~new_n55507_;
  assign new_n55509_ = ~\b[33]  & ~new_n55508_;
  assign new_n55510_ = ~new_n54673_ & new_n55083_;
  assign new_n55511_ = ~new_n55079_ & new_n55510_;
  assign new_n55512_ = ~new_n55080_ & ~new_n55083_;
  assign new_n55513_ = ~new_n55511_ & ~new_n55512_;
  assign new_n55514_ = ~new_n55248_ & ~new_n55513_;
  assign new_n55515_ = ~new_n54663_ & ~new_n55247_;
  assign new_n55516_ = ~new_n55246_ & new_n55515_;
  assign new_n55517_ = ~new_n55514_ & ~new_n55516_;
  assign new_n55518_ = ~\b[32]  & ~new_n55517_;
  assign new_n55519_ = ~new_n54682_ & new_n55078_;
  assign new_n55520_ = ~new_n55074_ & new_n55519_;
  assign new_n55521_ = ~new_n55075_ & ~new_n55078_;
  assign new_n55522_ = ~new_n55520_ & ~new_n55521_;
  assign new_n55523_ = ~new_n55248_ & ~new_n55522_;
  assign new_n55524_ = ~new_n54672_ & ~new_n55247_;
  assign new_n55525_ = ~new_n55246_ & new_n55524_;
  assign new_n55526_ = ~new_n55523_ & ~new_n55525_;
  assign new_n55527_ = ~\b[31]  & ~new_n55526_;
  assign new_n55528_ = ~new_n54691_ & new_n55073_;
  assign new_n55529_ = ~new_n55069_ & new_n55528_;
  assign new_n55530_ = ~new_n55070_ & ~new_n55073_;
  assign new_n55531_ = ~new_n55529_ & ~new_n55530_;
  assign new_n55532_ = ~new_n55248_ & ~new_n55531_;
  assign new_n55533_ = ~new_n54681_ & ~new_n55247_;
  assign new_n55534_ = ~new_n55246_ & new_n55533_;
  assign new_n55535_ = ~new_n55532_ & ~new_n55534_;
  assign new_n55536_ = ~\b[30]  & ~new_n55535_;
  assign new_n55537_ = ~new_n54700_ & new_n55068_;
  assign new_n55538_ = ~new_n55064_ & new_n55537_;
  assign new_n55539_ = ~new_n55065_ & ~new_n55068_;
  assign new_n55540_ = ~new_n55538_ & ~new_n55539_;
  assign new_n55541_ = ~new_n55248_ & ~new_n55540_;
  assign new_n55542_ = ~new_n54690_ & ~new_n55247_;
  assign new_n55543_ = ~new_n55246_ & new_n55542_;
  assign new_n55544_ = ~new_n55541_ & ~new_n55543_;
  assign new_n55545_ = ~\b[29]  & ~new_n55544_;
  assign new_n55546_ = ~new_n54709_ & new_n55063_;
  assign new_n55547_ = ~new_n55059_ & new_n55546_;
  assign new_n55548_ = ~new_n55060_ & ~new_n55063_;
  assign new_n55549_ = ~new_n55547_ & ~new_n55548_;
  assign new_n55550_ = ~new_n55248_ & ~new_n55549_;
  assign new_n55551_ = ~new_n54699_ & ~new_n55247_;
  assign new_n55552_ = ~new_n55246_ & new_n55551_;
  assign new_n55553_ = ~new_n55550_ & ~new_n55552_;
  assign new_n55554_ = ~\b[28]  & ~new_n55553_;
  assign new_n55555_ = ~new_n54718_ & new_n55058_;
  assign new_n55556_ = ~new_n55054_ & new_n55555_;
  assign new_n55557_ = ~new_n55055_ & ~new_n55058_;
  assign new_n55558_ = ~new_n55556_ & ~new_n55557_;
  assign new_n55559_ = ~new_n55248_ & ~new_n55558_;
  assign new_n55560_ = ~new_n54708_ & ~new_n55247_;
  assign new_n55561_ = ~new_n55246_ & new_n55560_;
  assign new_n55562_ = ~new_n55559_ & ~new_n55561_;
  assign new_n55563_ = ~\b[27]  & ~new_n55562_;
  assign new_n55564_ = ~new_n54727_ & new_n55053_;
  assign new_n55565_ = ~new_n55049_ & new_n55564_;
  assign new_n55566_ = ~new_n55050_ & ~new_n55053_;
  assign new_n55567_ = ~new_n55565_ & ~new_n55566_;
  assign new_n55568_ = ~new_n55248_ & ~new_n55567_;
  assign new_n55569_ = ~new_n54717_ & ~new_n55247_;
  assign new_n55570_ = ~new_n55246_ & new_n55569_;
  assign new_n55571_ = ~new_n55568_ & ~new_n55570_;
  assign new_n55572_ = ~\b[26]  & ~new_n55571_;
  assign new_n55573_ = ~new_n54736_ & new_n55048_;
  assign new_n55574_ = ~new_n55044_ & new_n55573_;
  assign new_n55575_ = ~new_n55045_ & ~new_n55048_;
  assign new_n55576_ = ~new_n55574_ & ~new_n55575_;
  assign new_n55577_ = ~new_n55248_ & ~new_n55576_;
  assign new_n55578_ = ~new_n54726_ & ~new_n55247_;
  assign new_n55579_ = ~new_n55246_ & new_n55578_;
  assign new_n55580_ = ~new_n55577_ & ~new_n55579_;
  assign new_n55581_ = ~\b[25]  & ~new_n55580_;
  assign new_n55582_ = ~new_n54745_ & new_n55043_;
  assign new_n55583_ = ~new_n55039_ & new_n55582_;
  assign new_n55584_ = ~new_n55040_ & ~new_n55043_;
  assign new_n55585_ = ~new_n55583_ & ~new_n55584_;
  assign new_n55586_ = ~new_n55248_ & ~new_n55585_;
  assign new_n55587_ = ~new_n54735_ & ~new_n55247_;
  assign new_n55588_ = ~new_n55246_ & new_n55587_;
  assign new_n55589_ = ~new_n55586_ & ~new_n55588_;
  assign new_n55590_ = ~\b[24]  & ~new_n55589_;
  assign new_n55591_ = ~new_n54754_ & new_n55038_;
  assign new_n55592_ = ~new_n55034_ & new_n55591_;
  assign new_n55593_ = ~new_n55035_ & ~new_n55038_;
  assign new_n55594_ = ~new_n55592_ & ~new_n55593_;
  assign new_n55595_ = ~new_n55248_ & ~new_n55594_;
  assign new_n55596_ = ~new_n54744_ & ~new_n55247_;
  assign new_n55597_ = ~new_n55246_ & new_n55596_;
  assign new_n55598_ = ~new_n55595_ & ~new_n55597_;
  assign new_n55599_ = ~\b[23]  & ~new_n55598_;
  assign new_n55600_ = ~new_n54763_ & new_n55033_;
  assign new_n55601_ = ~new_n55029_ & new_n55600_;
  assign new_n55602_ = ~new_n55030_ & ~new_n55033_;
  assign new_n55603_ = ~new_n55601_ & ~new_n55602_;
  assign new_n55604_ = ~new_n55248_ & ~new_n55603_;
  assign new_n55605_ = ~new_n54753_ & ~new_n55247_;
  assign new_n55606_ = ~new_n55246_ & new_n55605_;
  assign new_n55607_ = ~new_n55604_ & ~new_n55606_;
  assign new_n55608_ = ~\b[22]  & ~new_n55607_;
  assign new_n55609_ = ~new_n54772_ & new_n55028_;
  assign new_n55610_ = ~new_n55024_ & new_n55609_;
  assign new_n55611_ = ~new_n55025_ & ~new_n55028_;
  assign new_n55612_ = ~new_n55610_ & ~new_n55611_;
  assign new_n55613_ = ~new_n55248_ & ~new_n55612_;
  assign new_n55614_ = ~new_n54762_ & ~new_n55247_;
  assign new_n55615_ = ~new_n55246_ & new_n55614_;
  assign new_n55616_ = ~new_n55613_ & ~new_n55615_;
  assign new_n55617_ = ~\b[21]  & ~new_n55616_;
  assign new_n55618_ = ~new_n54781_ & new_n55023_;
  assign new_n55619_ = ~new_n55019_ & new_n55618_;
  assign new_n55620_ = ~new_n55020_ & ~new_n55023_;
  assign new_n55621_ = ~new_n55619_ & ~new_n55620_;
  assign new_n55622_ = ~new_n55248_ & ~new_n55621_;
  assign new_n55623_ = ~new_n54771_ & ~new_n55247_;
  assign new_n55624_ = ~new_n55246_ & new_n55623_;
  assign new_n55625_ = ~new_n55622_ & ~new_n55624_;
  assign new_n55626_ = ~\b[20]  & ~new_n55625_;
  assign new_n55627_ = ~new_n54790_ & new_n55018_;
  assign new_n55628_ = ~new_n55014_ & new_n55627_;
  assign new_n55629_ = ~new_n55015_ & ~new_n55018_;
  assign new_n55630_ = ~new_n55628_ & ~new_n55629_;
  assign new_n55631_ = ~new_n55248_ & ~new_n55630_;
  assign new_n55632_ = ~new_n54780_ & ~new_n55247_;
  assign new_n55633_ = ~new_n55246_ & new_n55632_;
  assign new_n55634_ = ~new_n55631_ & ~new_n55633_;
  assign new_n55635_ = ~\b[19]  & ~new_n55634_;
  assign new_n55636_ = ~new_n54799_ & new_n55013_;
  assign new_n55637_ = ~new_n55009_ & new_n55636_;
  assign new_n55638_ = ~new_n55010_ & ~new_n55013_;
  assign new_n55639_ = ~new_n55637_ & ~new_n55638_;
  assign new_n55640_ = ~new_n55248_ & ~new_n55639_;
  assign new_n55641_ = ~new_n54789_ & ~new_n55247_;
  assign new_n55642_ = ~new_n55246_ & new_n55641_;
  assign new_n55643_ = ~new_n55640_ & ~new_n55642_;
  assign new_n55644_ = ~\b[18]  & ~new_n55643_;
  assign new_n55645_ = ~new_n54808_ & new_n55008_;
  assign new_n55646_ = ~new_n55004_ & new_n55645_;
  assign new_n55647_ = ~new_n55005_ & ~new_n55008_;
  assign new_n55648_ = ~new_n55646_ & ~new_n55647_;
  assign new_n55649_ = ~new_n55248_ & ~new_n55648_;
  assign new_n55650_ = ~new_n54798_ & ~new_n55247_;
  assign new_n55651_ = ~new_n55246_ & new_n55650_;
  assign new_n55652_ = ~new_n55649_ & ~new_n55651_;
  assign new_n55653_ = ~\b[17]  & ~new_n55652_;
  assign new_n55654_ = ~new_n54817_ & new_n55003_;
  assign new_n55655_ = ~new_n54999_ & new_n55654_;
  assign new_n55656_ = ~new_n55000_ & ~new_n55003_;
  assign new_n55657_ = ~new_n55655_ & ~new_n55656_;
  assign new_n55658_ = ~new_n55248_ & ~new_n55657_;
  assign new_n55659_ = ~new_n54807_ & ~new_n55247_;
  assign new_n55660_ = ~new_n55246_ & new_n55659_;
  assign new_n55661_ = ~new_n55658_ & ~new_n55660_;
  assign new_n55662_ = ~\b[16]  & ~new_n55661_;
  assign new_n55663_ = ~new_n54826_ & new_n54998_;
  assign new_n55664_ = ~new_n54994_ & new_n55663_;
  assign new_n55665_ = ~new_n54995_ & ~new_n54998_;
  assign new_n55666_ = ~new_n55664_ & ~new_n55665_;
  assign new_n55667_ = ~new_n55248_ & ~new_n55666_;
  assign new_n55668_ = ~new_n54816_ & ~new_n55247_;
  assign new_n55669_ = ~new_n55246_ & new_n55668_;
  assign new_n55670_ = ~new_n55667_ & ~new_n55669_;
  assign new_n55671_ = ~\b[15]  & ~new_n55670_;
  assign new_n55672_ = ~new_n54835_ & new_n54993_;
  assign new_n55673_ = ~new_n54989_ & new_n55672_;
  assign new_n55674_ = ~new_n54990_ & ~new_n54993_;
  assign new_n55675_ = ~new_n55673_ & ~new_n55674_;
  assign new_n55676_ = ~new_n55248_ & ~new_n55675_;
  assign new_n55677_ = ~new_n54825_ & ~new_n55247_;
  assign new_n55678_ = ~new_n55246_ & new_n55677_;
  assign new_n55679_ = ~new_n55676_ & ~new_n55678_;
  assign new_n55680_ = ~\b[14]  & ~new_n55679_;
  assign new_n55681_ = ~new_n54844_ & new_n54988_;
  assign new_n55682_ = ~new_n54984_ & new_n55681_;
  assign new_n55683_ = ~new_n54985_ & ~new_n54988_;
  assign new_n55684_ = ~new_n55682_ & ~new_n55683_;
  assign new_n55685_ = ~new_n55248_ & ~new_n55684_;
  assign new_n55686_ = ~new_n54834_ & ~new_n55247_;
  assign new_n55687_ = ~new_n55246_ & new_n55686_;
  assign new_n55688_ = ~new_n55685_ & ~new_n55687_;
  assign new_n55689_ = ~\b[13]  & ~new_n55688_;
  assign new_n55690_ = ~new_n54853_ & new_n54983_;
  assign new_n55691_ = ~new_n54979_ & new_n55690_;
  assign new_n55692_ = ~new_n54980_ & ~new_n54983_;
  assign new_n55693_ = ~new_n55691_ & ~new_n55692_;
  assign new_n55694_ = ~new_n55248_ & ~new_n55693_;
  assign new_n55695_ = ~new_n54843_ & ~new_n55247_;
  assign new_n55696_ = ~new_n55246_ & new_n55695_;
  assign new_n55697_ = ~new_n55694_ & ~new_n55696_;
  assign new_n55698_ = ~\b[12]  & ~new_n55697_;
  assign new_n55699_ = ~new_n54862_ & new_n54978_;
  assign new_n55700_ = ~new_n54974_ & new_n55699_;
  assign new_n55701_ = ~new_n54975_ & ~new_n54978_;
  assign new_n55702_ = ~new_n55700_ & ~new_n55701_;
  assign new_n55703_ = ~new_n55248_ & ~new_n55702_;
  assign new_n55704_ = ~new_n54852_ & ~new_n55247_;
  assign new_n55705_ = ~new_n55246_ & new_n55704_;
  assign new_n55706_ = ~new_n55703_ & ~new_n55705_;
  assign new_n55707_ = ~\b[11]  & ~new_n55706_;
  assign new_n55708_ = ~new_n54871_ & new_n54973_;
  assign new_n55709_ = ~new_n54969_ & new_n55708_;
  assign new_n55710_ = ~new_n54970_ & ~new_n54973_;
  assign new_n55711_ = ~new_n55709_ & ~new_n55710_;
  assign new_n55712_ = ~new_n55248_ & ~new_n55711_;
  assign new_n55713_ = ~new_n54861_ & ~new_n55247_;
  assign new_n55714_ = ~new_n55246_ & new_n55713_;
  assign new_n55715_ = ~new_n55712_ & ~new_n55714_;
  assign new_n55716_ = ~\b[10]  & ~new_n55715_;
  assign new_n55717_ = ~new_n54880_ & new_n54968_;
  assign new_n55718_ = ~new_n54964_ & new_n55717_;
  assign new_n55719_ = ~new_n54965_ & ~new_n54968_;
  assign new_n55720_ = ~new_n55718_ & ~new_n55719_;
  assign new_n55721_ = ~new_n55248_ & ~new_n55720_;
  assign new_n55722_ = ~new_n54870_ & ~new_n55247_;
  assign new_n55723_ = ~new_n55246_ & new_n55722_;
  assign new_n55724_ = ~new_n55721_ & ~new_n55723_;
  assign new_n55725_ = ~\b[9]  & ~new_n55724_;
  assign new_n55726_ = ~new_n54889_ & new_n54963_;
  assign new_n55727_ = ~new_n54959_ & new_n55726_;
  assign new_n55728_ = ~new_n54960_ & ~new_n54963_;
  assign new_n55729_ = ~new_n55727_ & ~new_n55728_;
  assign new_n55730_ = ~new_n55248_ & ~new_n55729_;
  assign new_n55731_ = ~new_n54879_ & ~new_n55247_;
  assign new_n55732_ = ~new_n55246_ & new_n55731_;
  assign new_n55733_ = ~new_n55730_ & ~new_n55732_;
  assign new_n55734_ = ~\b[8]  & ~new_n55733_;
  assign new_n55735_ = ~new_n54898_ & new_n54958_;
  assign new_n55736_ = ~new_n54954_ & new_n55735_;
  assign new_n55737_ = ~new_n54955_ & ~new_n54958_;
  assign new_n55738_ = ~new_n55736_ & ~new_n55737_;
  assign new_n55739_ = ~new_n55248_ & ~new_n55738_;
  assign new_n55740_ = ~new_n54888_ & ~new_n55247_;
  assign new_n55741_ = ~new_n55246_ & new_n55740_;
  assign new_n55742_ = ~new_n55739_ & ~new_n55741_;
  assign new_n55743_ = ~\b[7]  & ~new_n55742_;
  assign new_n55744_ = ~new_n54907_ & new_n54953_;
  assign new_n55745_ = ~new_n54949_ & new_n55744_;
  assign new_n55746_ = ~new_n54950_ & ~new_n54953_;
  assign new_n55747_ = ~new_n55745_ & ~new_n55746_;
  assign new_n55748_ = ~new_n55248_ & ~new_n55747_;
  assign new_n55749_ = ~new_n54897_ & ~new_n55247_;
  assign new_n55750_ = ~new_n55246_ & new_n55749_;
  assign new_n55751_ = ~new_n55748_ & ~new_n55750_;
  assign new_n55752_ = ~\b[6]  & ~new_n55751_;
  assign new_n55753_ = ~new_n54916_ & new_n54948_;
  assign new_n55754_ = ~new_n54944_ & new_n55753_;
  assign new_n55755_ = ~new_n54945_ & ~new_n54948_;
  assign new_n55756_ = ~new_n55754_ & ~new_n55755_;
  assign new_n55757_ = ~new_n55248_ & ~new_n55756_;
  assign new_n55758_ = ~new_n54906_ & ~new_n55247_;
  assign new_n55759_ = ~new_n55246_ & new_n55758_;
  assign new_n55760_ = ~new_n55757_ & ~new_n55759_;
  assign new_n55761_ = ~\b[5]  & ~new_n55760_;
  assign new_n55762_ = ~new_n54924_ & new_n54943_;
  assign new_n55763_ = ~new_n54939_ & new_n55762_;
  assign new_n55764_ = ~new_n54940_ & ~new_n54943_;
  assign new_n55765_ = ~new_n55763_ & ~new_n55764_;
  assign new_n55766_ = ~new_n55248_ & ~new_n55765_;
  assign new_n55767_ = ~new_n54915_ & ~new_n55247_;
  assign new_n55768_ = ~new_n55246_ & new_n55767_;
  assign new_n55769_ = ~new_n55766_ & ~new_n55768_;
  assign new_n55770_ = ~\b[4]  & ~new_n55769_;
  assign new_n55771_ = ~new_n54934_ & new_n54938_;
  assign new_n55772_ = ~new_n54933_ & new_n55771_;
  assign new_n55773_ = ~new_n54935_ & ~new_n54938_;
  assign new_n55774_ = ~new_n55772_ & ~new_n55773_;
  assign new_n55775_ = ~new_n55248_ & ~new_n55774_;
  assign new_n55776_ = ~new_n54923_ & ~new_n55247_;
  assign new_n55777_ = ~new_n55246_ & new_n55776_;
  assign new_n55778_ = ~new_n55775_ & ~new_n55777_;
  assign new_n55779_ = ~\b[3]  & ~new_n55778_;
  assign new_n55780_ = new_n26919_ & ~new_n54931_;
  assign new_n55781_ = ~new_n54929_ & new_n55780_;
  assign new_n55782_ = ~new_n54933_ & ~new_n55781_;
  assign new_n55783_ = ~new_n55248_ & new_n55782_;
  assign new_n55784_ = ~new_n54928_ & ~new_n55247_;
  assign new_n55785_ = ~new_n55246_ & new_n55784_;
  assign new_n55786_ = ~new_n55783_ & ~new_n55785_;
  assign new_n55787_ = ~\b[2]  & ~new_n55786_;
  assign new_n55788_ = \b[0]  & ~new_n55248_;
  assign new_n55789_ = \a[2]  & ~new_n55788_;
  assign new_n55790_ = new_n26919_ & ~new_n55248_;
  assign new_n55791_ = ~new_n55789_ & ~new_n55790_;
  assign new_n55792_ = \b[1]  & ~new_n55791_;
  assign new_n55793_ = ~\b[1]  & ~new_n55790_;
  assign new_n55794_ = ~new_n55789_ & new_n55793_;
  assign new_n55795_ = ~new_n55792_ & ~new_n55794_;
  assign new_n55796_ = ~new_n27783_ & ~new_n55795_;
  assign new_n55797_ = ~\b[1]  & ~new_n55791_;
  assign new_n55798_ = ~new_n55796_ & ~new_n55797_;
  assign new_n55799_ = \b[2]  & ~new_n55785_;
  assign new_n55800_ = ~new_n55783_ & new_n55799_;
  assign new_n55801_ = ~new_n55787_ & ~new_n55800_;
  assign new_n55802_ = ~new_n55798_ & new_n55801_;
  assign new_n55803_ = ~new_n55787_ & ~new_n55802_;
  assign new_n55804_ = \b[3]  & ~new_n55777_;
  assign new_n55805_ = ~new_n55775_ & new_n55804_;
  assign new_n55806_ = ~new_n55779_ & ~new_n55805_;
  assign new_n55807_ = ~new_n55803_ & new_n55806_;
  assign new_n55808_ = ~new_n55779_ & ~new_n55807_;
  assign new_n55809_ = \b[4]  & ~new_n55768_;
  assign new_n55810_ = ~new_n55766_ & new_n55809_;
  assign new_n55811_ = ~new_n55770_ & ~new_n55810_;
  assign new_n55812_ = ~new_n55808_ & new_n55811_;
  assign new_n55813_ = ~new_n55770_ & ~new_n55812_;
  assign new_n55814_ = \b[5]  & ~new_n55759_;
  assign new_n55815_ = ~new_n55757_ & new_n55814_;
  assign new_n55816_ = ~new_n55761_ & ~new_n55815_;
  assign new_n55817_ = ~new_n55813_ & new_n55816_;
  assign new_n55818_ = ~new_n55761_ & ~new_n55817_;
  assign new_n55819_ = \b[6]  & ~new_n55750_;
  assign new_n55820_ = ~new_n55748_ & new_n55819_;
  assign new_n55821_ = ~new_n55752_ & ~new_n55820_;
  assign new_n55822_ = ~new_n55818_ & new_n55821_;
  assign new_n55823_ = ~new_n55752_ & ~new_n55822_;
  assign new_n55824_ = \b[7]  & ~new_n55741_;
  assign new_n55825_ = ~new_n55739_ & new_n55824_;
  assign new_n55826_ = ~new_n55743_ & ~new_n55825_;
  assign new_n55827_ = ~new_n55823_ & new_n55826_;
  assign new_n55828_ = ~new_n55743_ & ~new_n55827_;
  assign new_n55829_ = \b[8]  & ~new_n55732_;
  assign new_n55830_ = ~new_n55730_ & new_n55829_;
  assign new_n55831_ = ~new_n55734_ & ~new_n55830_;
  assign new_n55832_ = ~new_n55828_ & new_n55831_;
  assign new_n55833_ = ~new_n55734_ & ~new_n55832_;
  assign new_n55834_ = \b[9]  & ~new_n55723_;
  assign new_n55835_ = ~new_n55721_ & new_n55834_;
  assign new_n55836_ = ~new_n55725_ & ~new_n55835_;
  assign new_n55837_ = ~new_n55833_ & new_n55836_;
  assign new_n55838_ = ~new_n55725_ & ~new_n55837_;
  assign new_n55839_ = \b[10]  & ~new_n55714_;
  assign new_n55840_ = ~new_n55712_ & new_n55839_;
  assign new_n55841_ = ~new_n55716_ & ~new_n55840_;
  assign new_n55842_ = ~new_n55838_ & new_n55841_;
  assign new_n55843_ = ~new_n55716_ & ~new_n55842_;
  assign new_n55844_ = \b[11]  & ~new_n55705_;
  assign new_n55845_ = ~new_n55703_ & new_n55844_;
  assign new_n55846_ = ~new_n55707_ & ~new_n55845_;
  assign new_n55847_ = ~new_n55843_ & new_n55846_;
  assign new_n55848_ = ~new_n55707_ & ~new_n55847_;
  assign new_n55849_ = \b[12]  & ~new_n55696_;
  assign new_n55850_ = ~new_n55694_ & new_n55849_;
  assign new_n55851_ = ~new_n55698_ & ~new_n55850_;
  assign new_n55852_ = ~new_n55848_ & new_n55851_;
  assign new_n55853_ = ~new_n55698_ & ~new_n55852_;
  assign new_n55854_ = \b[13]  & ~new_n55687_;
  assign new_n55855_ = ~new_n55685_ & new_n55854_;
  assign new_n55856_ = ~new_n55689_ & ~new_n55855_;
  assign new_n55857_ = ~new_n55853_ & new_n55856_;
  assign new_n55858_ = ~new_n55689_ & ~new_n55857_;
  assign new_n55859_ = \b[14]  & ~new_n55678_;
  assign new_n55860_ = ~new_n55676_ & new_n55859_;
  assign new_n55861_ = ~new_n55680_ & ~new_n55860_;
  assign new_n55862_ = ~new_n55858_ & new_n55861_;
  assign new_n55863_ = ~new_n55680_ & ~new_n55862_;
  assign new_n55864_ = \b[15]  & ~new_n55669_;
  assign new_n55865_ = ~new_n55667_ & new_n55864_;
  assign new_n55866_ = ~new_n55671_ & ~new_n55865_;
  assign new_n55867_ = ~new_n55863_ & new_n55866_;
  assign new_n55868_ = ~new_n55671_ & ~new_n55867_;
  assign new_n55869_ = \b[16]  & ~new_n55660_;
  assign new_n55870_ = ~new_n55658_ & new_n55869_;
  assign new_n55871_ = ~new_n55662_ & ~new_n55870_;
  assign new_n55872_ = ~new_n55868_ & new_n55871_;
  assign new_n55873_ = ~new_n55662_ & ~new_n55872_;
  assign new_n55874_ = \b[17]  & ~new_n55651_;
  assign new_n55875_ = ~new_n55649_ & new_n55874_;
  assign new_n55876_ = ~new_n55653_ & ~new_n55875_;
  assign new_n55877_ = ~new_n55873_ & new_n55876_;
  assign new_n55878_ = ~new_n55653_ & ~new_n55877_;
  assign new_n55879_ = \b[18]  & ~new_n55642_;
  assign new_n55880_ = ~new_n55640_ & new_n55879_;
  assign new_n55881_ = ~new_n55644_ & ~new_n55880_;
  assign new_n55882_ = ~new_n55878_ & new_n55881_;
  assign new_n55883_ = ~new_n55644_ & ~new_n55882_;
  assign new_n55884_ = \b[19]  & ~new_n55633_;
  assign new_n55885_ = ~new_n55631_ & new_n55884_;
  assign new_n55886_ = ~new_n55635_ & ~new_n55885_;
  assign new_n55887_ = ~new_n55883_ & new_n55886_;
  assign new_n55888_ = ~new_n55635_ & ~new_n55887_;
  assign new_n55889_ = \b[20]  & ~new_n55624_;
  assign new_n55890_ = ~new_n55622_ & new_n55889_;
  assign new_n55891_ = ~new_n55626_ & ~new_n55890_;
  assign new_n55892_ = ~new_n55888_ & new_n55891_;
  assign new_n55893_ = ~new_n55626_ & ~new_n55892_;
  assign new_n55894_ = \b[21]  & ~new_n55615_;
  assign new_n55895_ = ~new_n55613_ & new_n55894_;
  assign new_n55896_ = ~new_n55617_ & ~new_n55895_;
  assign new_n55897_ = ~new_n55893_ & new_n55896_;
  assign new_n55898_ = ~new_n55617_ & ~new_n55897_;
  assign new_n55899_ = \b[22]  & ~new_n55606_;
  assign new_n55900_ = ~new_n55604_ & new_n55899_;
  assign new_n55901_ = ~new_n55608_ & ~new_n55900_;
  assign new_n55902_ = ~new_n55898_ & new_n55901_;
  assign new_n55903_ = ~new_n55608_ & ~new_n55902_;
  assign new_n55904_ = \b[23]  & ~new_n55597_;
  assign new_n55905_ = ~new_n55595_ & new_n55904_;
  assign new_n55906_ = ~new_n55599_ & ~new_n55905_;
  assign new_n55907_ = ~new_n55903_ & new_n55906_;
  assign new_n55908_ = ~new_n55599_ & ~new_n55907_;
  assign new_n55909_ = \b[24]  & ~new_n55588_;
  assign new_n55910_ = ~new_n55586_ & new_n55909_;
  assign new_n55911_ = ~new_n55590_ & ~new_n55910_;
  assign new_n55912_ = ~new_n55908_ & new_n55911_;
  assign new_n55913_ = ~new_n55590_ & ~new_n55912_;
  assign new_n55914_ = \b[25]  & ~new_n55579_;
  assign new_n55915_ = ~new_n55577_ & new_n55914_;
  assign new_n55916_ = ~new_n55581_ & ~new_n55915_;
  assign new_n55917_ = ~new_n55913_ & new_n55916_;
  assign new_n55918_ = ~new_n55581_ & ~new_n55917_;
  assign new_n55919_ = \b[26]  & ~new_n55570_;
  assign new_n55920_ = ~new_n55568_ & new_n55919_;
  assign new_n55921_ = ~new_n55572_ & ~new_n55920_;
  assign new_n55922_ = ~new_n55918_ & new_n55921_;
  assign new_n55923_ = ~new_n55572_ & ~new_n55922_;
  assign new_n55924_ = \b[27]  & ~new_n55561_;
  assign new_n55925_ = ~new_n55559_ & new_n55924_;
  assign new_n55926_ = ~new_n55563_ & ~new_n55925_;
  assign new_n55927_ = ~new_n55923_ & new_n55926_;
  assign new_n55928_ = ~new_n55563_ & ~new_n55927_;
  assign new_n55929_ = \b[28]  & ~new_n55552_;
  assign new_n55930_ = ~new_n55550_ & new_n55929_;
  assign new_n55931_ = ~new_n55554_ & ~new_n55930_;
  assign new_n55932_ = ~new_n55928_ & new_n55931_;
  assign new_n55933_ = ~new_n55554_ & ~new_n55932_;
  assign new_n55934_ = \b[29]  & ~new_n55543_;
  assign new_n55935_ = ~new_n55541_ & new_n55934_;
  assign new_n55936_ = ~new_n55545_ & ~new_n55935_;
  assign new_n55937_ = ~new_n55933_ & new_n55936_;
  assign new_n55938_ = ~new_n55545_ & ~new_n55937_;
  assign new_n55939_ = \b[30]  & ~new_n55534_;
  assign new_n55940_ = ~new_n55532_ & new_n55939_;
  assign new_n55941_ = ~new_n55536_ & ~new_n55940_;
  assign new_n55942_ = ~new_n55938_ & new_n55941_;
  assign new_n55943_ = ~new_n55536_ & ~new_n55942_;
  assign new_n55944_ = \b[31]  & ~new_n55525_;
  assign new_n55945_ = ~new_n55523_ & new_n55944_;
  assign new_n55946_ = ~new_n55527_ & ~new_n55945_;
  assign new_n55947_ = ~new_n55943_ & new_n55946_;
  assign new_n55948_ = ~new_n55527_ & ~new_n55947_;
  assign new_n55949_ = \b[32]  & ~new_n55516_;
  assign new_n55950_ = ~new_n55514_ & new_n55949_;
  assign new_n55951_ = ~new_n55518_ & ~new_n55950_;
  assign new_n55952_ = ~new_n55948_ & new_n55951_;
  assign new_n55953_ = ~new_n55518_ & ~new_n55952_;
  assign new_n55954_ = \b[33]  & ~new_n55507_;
  assign new_n55955_ = ~new_n55505_ & new_n55954_;
  assign new_n55956_ = ~new_n55509_ & ~new_n55955_;
  assign new_n55957_ = ~new_n55953_ & new_n55956_;
  assign new_n55958_ = ~new_n55509_ & ~new_n55957_;
  assign new_n55959_ = \b[34]  & ~new_n55498_;
  assign new_n55960_ = ~new_n55496_ & new_n55959_;
  assign new_n55961_ = ~new_n55500_ & ~new_n55960_;
  assign new_n55962_ = ~new_n55958_ & new_n55961_;
  assign new_n55963_ = ~new_n55500_ & ~new_n55962_;
  assign new_n55964_ = \b[35]  & ~new_n55489_;
  assign new_n55965_ = ~new_n55487_ & new_n55964_;
  assign new_n55966_ = ~new_n55491_ & ~new_n55965_;
  assign new_n55967_ = ~new_n55963_ & new_n55966_;
  assign new_n55968_ = ~new_n55491_ & ~new_n55967_;
  assign new_n55969_ = \b[36]  & ~new_n55480_;
  assign new_n55970_ = ~new_n55478_ & new_n55969_;
  assign new_n55971_ = ~new_n55482_ & ~new_n55970_;
  assign new_n55972_ = ~new_n55968_ & new_n55971_;
  assign new_n55973_ = ~new_n55482_ & ~new_n55972_;
  assign new_n55974_ = \b[37]  & ~new_n55471_;
  assign new_n55975_ = ~new_n55469_ & new_n55974_;
  assign new_n55976_ = ~new_n55473_ & ~new_n55975_;
  assign new_n55977_ = ~new_n55973_ & new_n55976_;
  assign new_n55978_ = ~new_n55473_ & ~new_n55977_;
  assign new_n55979_ = \b[38]  & ~new_n55462_;
  assign new_n55980_ = ~new_n55460_ & new_n55979_;
  assign new_n55981_ = ~new_n55464_ & ~new_n55980_;
  assign new_n55982_ = ~new_n55978_ & new_n55981_;
  assign new_n55983_ = ~new_n55464_ & ~new_n55982_;
  assign new_n55984_ = \b[39]  & ~new_n55453_;
  assign new_n55985_ = ~new_n55451_ & new_n55984_;
  assign new_n55986_ = ~new_n55455_ & ~new_n55985_;
  assign new_n55987_ = ~new_n55983_ & new_n55986_;
  assign new_n55988_ = ~new_n55455_ & ~new_n55987_;
  assign new_n55989_ = \b[40]  & ~new_n55444_;
  assign new_n55990_ = ~new_n55442_ & new_n55989_;
  assign new_n55991_ = ~new_n55446_ & ~new_n55990_;
  assign new_n55992_ = ~new_n55988_ & new_n55991_;
  assign new_n55993_ = ~new_n55446_ & ~new_n55992_;
  assign new_n55994_ = \b[41]  & ~new_n55435_;
  assign new_n55995_ = ~new_n55433_ & new_n55994_;
  assign new_n55996_ = ~new_n55437_ & ~new_n55995_;
  assign new_n55997_ = ~new_n55993_ & new_n55996_;
  assign new_n55998_ = ~new_n55437_ & ~new_n55997_;
  assign new_n55999_ = \b[42]  & ~new_n55426_;
  assign new_n56000_ = ~new_n55424_ & new_n55999_;
  assign new_n56001_ = ~new_n55428_ & ~new_n56000_;
  assign new_n56002_ = ~new_n55998_ & new_n56001_;
  assign new_n56003_ = ~new_n55428_ & ~new_n56002_;
  assign new_n56004_ = \b[43]  & ~new_n55417_;
  assign new_n56005_ = ~new_n55415_ & new_n56004_;
  assign new_n56006_ = ~new_n55419_ & ~new_n56005_;
  assign new_n56007_ = ~new_n56003_ & new_n56006_;
  assign new_n56008_ = ~new_n55419_ & ~new_n56007_;
  assign new_n56009_ = \b[44]  & ~new_n55408_;
  assign new_n56010_ = ~new_n55406_ & new_n56009_;
  assign new_n56011_ = ~new_n55410_ & ~new_n56010_;
  assign new_n56012_ = ~new_n56008_ & new_n56011_;
  assign new_n56013_ = ~new_n55410_ & ~new_n56012_;
  assign new_n56014_ = \b[45]  & ~new_n55399_;
  assign new_n56015_ = ~new_n55397_ & new_n56014_;
  assign new_n56016_ = ~new_n55401_ & ~new_n56015_;
  assign new_n56017_ = ~new_n56013_ & new_n56016_;
  assign new_n56018_ = ~new_n55401_ & ~new_n56017_;
  assign new_n56019_ = \b[46]  & ~new_n55390_;
  assign new_n56020_ = ~new_n55388_ & new_n56019_;
  assign new_n56021_ = ~new_n55392_ & ~new_n56020_;
  assign new_n56022_ = ~new_n56018_ & new_n56021_;
  assign new_n56023_ = ~new_n55392_ & ~new_n56022_;
  assign new_n56024_ = \b[47]  & ~new_n55381_;
  assign new_n56025_ = ~new_n55379_ & new_n56024_;
  assign new_n56026_ = ~new_n55383_ & ~new_n56025_;
  assign new_n56027_ = ~new_n56023_ & new_n56026_;
  assign new_n56028_ = ~new_n55383_ & ~new_n56027_;
  assign new_n56029_ = \b[48]  & ~new_n55372_;
  assign new_n56030_ = ~new_n55370_ & new_n56029_;
  assign new_n56031_ = ~new_n55374_ & ~new_n56030_;
  assign new_n56032_ = ~new_n56028_ & new_n56031_;
  assign new_n56033_ = ~new_n55374_ & ~new_n56032_;
  assign new_n56034_ = \b[49]  & ~new_n55363_;
  assign new_n56035_ = ~new_n55361_ & new_n56034_;
  assign new_n56036_ = ~new_n55365_ & ~new_n56035_;
  assign new_n56037_ = ~new_n56033_ & new_n56036_;
  assign new_n56038_ = ~new_n55365_ & ~new_n56037_;
  assign new_n56039_ = \b[50]  & ~new_n55354_;
  assign new_n56040_ = ~new_n55352_ & new_n56039_;
  assign new_n56041_ = ~new_n55356_ & ~new_n56040_;
  assign new_n56042_ = ~new_n56038_ & new_n56041_;
  assign new_n56043_ = ~new_n55356_ & ~new_n56042_;
  assign new_n56044_ = \b[51]  & ~new_n55345_;
  assign new_n56045_ = ~new_n55343_ & new_n56044_;
  assign new_n56046_ = ~new_n55347_ & ~new_n56045_;
  assign new_n56047_ = ~new_n56043_ & new_n56046_;
  assign new_n56048_ = ~new_n55347_ & ~new_n56047_;
  assign new_n56049_ = \b[52]  & ~new_n55336_;
  assign new_n56050_ = ~new_n55334_ & new_n56049_;
  assign new_n56051_ = ~new_n55338_ & ~new_n56050_;
  assign new_n56052_ = ~new_n56048_ & new_n56051_;
  assign new_n56053_ = ~new_n55338_ & ~new_n56052_;
  assign new_n56054_ = \b[53]  & ~new_n55327_;
  assign new_n56055_ = ~new_n55325_ & new_n56054_;
  assign new_n56056_ = ~new_n55329_ & ~new_n56055_;
  assign new_n56057_ = ~new_n56053_ & new_n56056_;
  assign new_n56058_ = ~new_n55329_ & ~new_n56057_;
  assign new_n56059_ = \b[54]  & ~new_n55318_;
  assign new_n56060_ = ~new_n55316_ & new_n56059_;
  assign new_n56061_ = ~new_n55320_ & ~new_n56060_;
  assign new_n56062_ = ~new_n56058_ & new_n56061_;
  assign new_n56063_ = ~new_n55320_ & ~new_n56062_;
  assign new_n56064_ = \b[55]  & ~new_n55309_;
  assign new_n56065_ = ~new_n55307_ & new_n56064_;
  assign new_n56066_ = ~new_n55311_ & ~new_n56065_;
  assign new_n56067_ = ~new_n56063_ & new_n56066_;
  assign new_n56068_ = ~new_n55311_ & ~new_n56067_;
  assign new_n56069_ = \b[56]  & ~new_n55300_;
  assign new_n56070_ = ~new_n55298_ & new_n56069_;
  assign new_n56071_ = ~new_n55302_ & ~new_n56070_;
  assign new_n56072_ = ~new_n56068_ & new_n56071_;
  assign new_n56073_ = ~new_n55302_ & ~new_n56072_;
  assign new_n56074_ = \b[57]  & ~new_n55291_;
  assign new_n56075_ = ~new_n55289_ & new_n56074_;
  assign new_n56076_ = ~new_n55293_ & ~new_n56075_;
  assign new_n56077_ = ~new_n56073_ & new_n56076_;
  assign new_n56078_ = ~new_n55293_ & ~new_n56077_;
  assign new_n56079_ = \b[58]  & ~new_n55282_;
  assign new_n56080_ = ~new_n55280_ & new_n56079_;
  assign new_n56081_ = ~new_n55284_ & ~new_n56080_;
  assign new_n56082_ = ~new_n56078_ & new_n56081_;
  assign new_n56083_ = ~new_n55284_ & ~new_n56082_;
  assign new_n56084_ = \b[59]  & ~new_n55273_;
  assign new_n56085_ = ~new_n55271_ & new_n56084_;
  assign new_n56086_ = ~new_n55275_ & ~new_n56085_;
  assign new_n56087_ = ~new_n56083_ & new_n56086_;
  assign new_n56088_ = ~new_n55275_ & ~new_n56087_;
  assign new_n56089_ = \b[60]  & ~new_n55264_;
  assign new_n56090_ = ~new_n55262_ & new_n56089_;
  assign new_n56091_ = ~new_n55266_ & ~new_n56090_;
  assign new_n56092_ = ~new_n56088_ & new_n56091_;
  assign new_n56093_ = ~new_n55266_ & ~new_n56092_;
  assign new_n56094_ = \b[61]  & ~new_n55255_;
  assign new_n56095_ = ~new_n55253_ & new_n56094_;
  assign new_n56096_ = ~new_n55257_ & ~new_n56095_;
  assign new_n56097_ = ~new_n56093_ & new_n56096_;
  assign new_n56098_ = ~new_n55257_ & ~new_n56097_;
  assign new_n56099_ = ~new_n54403_ & ~new_n55243_;
  assign new_n56100_ = ~new_n55241_ & new_n56099_;
  assign new_n56101_ = ~new_n55229_ & new_n56100_;
  assign new_n56102_ = ~new_n55241_ & ~new_n55243_;
  assign new_n56103_ = ~new_n55230_ & ~new_n56102_;
  assign new_n56104_ = ~new_n56101_ & ~new_n56103_;
  assign new_n56105_ = ~new_n55248_ & ~new_n56104_;
  assign new_n56106_ = ~new_n55240_ & ~new_n55247_;
  assign new_n56107_ = ~new_n55246_ & new_n56106_;
  assign new_n56108_ = ~new_n56105_ & ~new_n56107_;
  assign new_n56109_ = ~\b[62]  & ~new_n56108_;
  assign new_n56110_ = \b[62]  & ~new_n56107_;
  assign new_n56111_ = ~new_n56105_ & new_n56110_;
  assign new_n56112_ = ~\b[63]  & ~new_n56111_;
  assign new_n56113_ = ~new_n56109_ & new_n56112_;
  assign new_n56114_ = ~new_n56098_ & new_n56113_;
  assign new_n56115_ = new_n279_ & ~new_n56108_;
  assign new_n56116_ = ~new_n56114_ & ~new_n56115_;
  assign new_n56117_ = ~new_n55257_ & ~new_n56111_;
  assign new_n56118_ = ~new_n56109_ & new_n56117_;
  assign new_n56119_ = ~new_n56097_ & new_n56118_;
  assign new_n56120_ = ~new_n56109_ & ~new_n56111_;
  assign new_n56121_ = ~new_n56098_ & ~new_n56120_;
  assign new_n56122_ = ~new_n56119_ & ~new_n56121_;
  assign new_n56123_ = ~new_n56116_ & ~new_n56122_;
  assign new_n56124_ = ~new_n56108_ & ~new_n56115_;
  assign new_n56125_ = ~new_n56114_ & new_n56124_;
  assign new_n56126_ = ~new_n56123_ & ~new_n56125_;
  assign new_n56127_ = ~\b[63]  & ~new_n56126_;
  assign new_n56128_ = ~new_n55266_ & new_n56096_;
  assign new_n56129_ = ~new_n56092_ & new_n56128_;
  assign new_n56130_ = ~new_n56093_ & ~new_n56096_;
  assign new_n56131_ = ~new_n56129_ & ~new_n56130_;
  assign new_n56132_ = ~new_n56116_ & ~new_n56131_;
  assign new_n56133_ = ~new_n55256_ & ~new_n56115_;
  assign new_n56134_ = ~new_n56114_ & new_n56133_;
  assign new_n56135_ = ~new_n56132_ & ~new_n56134_;
  assign new_n56136_ = ~\b[62]  & ~new_n56135_;
  assign new_n56137_ = ~new_n55275_ & new_n56091_;
  assign new_n56138_ = ~new_n56087_ & new_n56137_;
  assign new_n56139_ = ~new_n56088_ & ~new_n56091_;
  assign new_n56140_ = ~new_n56138_ & ~new_n56139_;
  assign new_n56141_ = ~new_n56116_ & ~new_n56140_;
  assign new_n56142_ = ~new_n55265_ & ~new_n56115_;
  assign new_n56143_ = ~new_n56114_ & new_n56142_;
  assign new_n56144_ = ~new_n56141_ & ~new_n56143_;
  assign new_n56145_ = ~\b[61]  & ~new_n56144_;
  assign new_n56146_ = ~new_n55284_ & new_n56086_;
  assign new_n56147_ = ~new_n56082_ & new_n56146_;
  assign new_n56148_ = ~new_n56083_ & ~new_n56086_;
  assign new_n56149_ = ~new_n56147_ & ~new_n56148_;
  assign new_n56150_ = ~new_n56116_ & ~new_n56149_;
  assign new_n56151_ = ~new_n55274_ & ~new_n56115_;
  assign new_n56152_ = ~new_n56114_ & new_n56151_;
  assign new_n56153_ = ~new_n56150_ & ~new_n56152_;
  assign new_n56154_ = ~\b[60]  & ~new_n56153_;
  assign new_n56155_ = ~new_n55293_ & new_n56081_;
  assign new_n56156_ = ~new_n56077_ & new_n56155_;
  assign new_n56157_ = ~new_n56078_ & ~new_n56081_;
  assign new_n56158_ = ~new_n56156_ & ~new_n56157_;
  assign new_n56159_ = ~new_n56116_ & ~new_n56158_;
  assign new_n56160_ = ~new_n55283_ & ~new_n56115_;
  assign new_n56161_ = ~new_n56114_ & new_n56160_;
  assign new_n56162_ = ~new_n56159_ & ~new_n56161_;
  assign new_n56163_ = ~\b[59]  & ~new_n56162_;
  assign new_n56164_ = ~new_n55302_ & new_n56076_;
  assign new_n56165_ = ~new_n56072_ & new_n56164_;
  assign new_n56166_ = ~new_n56073_ & ~new_n56076_;
  assign new_n56167_ = ~new_n56165_ & ~new_n56166_;
  assign new_n56168_ = ~new_n56116_ & ~new_n56167_;
  assign new_n56169_ = ~new_n55292_ & ~new_n56115_;
  assign new_n56170_ = ~new_n56114_ & new_n56169_;
  assign new_n56171_ = ~new_n56168_ & ~new_n56170_;
  assign new_n56172_ = ~\b[58]  & ~new_n56171_;
  assign new_n56173_ = ~new_n55311_ & new_n56071_;
  assign new_n56174_ = ~new_n56067_ & new_n56173_;
  assign new_n56175_ = ~new_n56068_ & ~new_n56071_;
  assign new_n56176_ = ~new_n56174_ & ~new_n56175_;
  assign new_n56177_ = ~new_n56116_ & ~new_n56176_;
  assign new_n56178_ = ~new_n55301_ & ~new_n56115_;
  assign new_n56179_ = ~new_n56114_ & new_n56178_;
  assign new_n56180_ = ~new_n56177_ & ~new_n56179_;
  assign new_n56181_ = ~\b[57]  & ~new_n56180_;
  assign new_n56182_ = ~new_n55320_ & new_n56066_;
  assign new_n56183_ = ~new_n56062_ & new_n56182_;
  assign new_n56184_ = ~new_n56063_ & ~new_n56066_;
  assign new_n56185_ = ~new_n56183_ & ~new_n56184_;
  assign new_n56186_ = ~new_n56116_ & ~new_n56185_;
  assign new_n56187_ = ~new_n55310_ & ~new_n56115_;
  assign new_n56188_ = ~new_n56114_ & new_n56187_;
  assign new_n56189_ = ~new_n56186_ & ~new_n56188_;
  assign new_n56190_ = ~\b[56]  & ~new_n56189_;
  assign new_n56191_ = ~new_n55329_ & new_n56061_;
  assign new_n56192_ = ~new_n56057_ & new_n56191_;
  assign new_n56193_ = ~new_n56058_ & ~new_n56061_;
  assign new_n56194_ = ~new_n56192_ & ~new_n56193_;
  assign new_n56195_ = ~new_n56116_ & ~new_n56194_;
  assign new_n56196_ = ~new_n55319_ & ~new_n56115_;
  assign new_n56197_ = ~new_n56114_ & new_n56196_;
  assign new_n56198_ = ~new_n56195_ & ~new_n56197_;
  assign new_n56199_ = ~\b[55]  & ~new_n56198_;
  assign new_n56200_ = ~new_n55338_ & new_n56056_;
  assign new_n56201_ = ~new_n56052_ & new_n56200_;
  assign new_n56202_ = ~new_n56053_ & ~new_n56056_;
  assign new_n56203_ = ~new_n56201_ & ~new_n56202_;
  assign new_n56204_ = ~new_n56116_ & ~new_n56203_;
  assign new_n56205_ = ~new_n55328_ & ~new_n56115_;
  assign new_n56206_ = ~new_n56114_ & new_n56205_;
  assign new_n56207_ = ~new_n56204_ & ~new_n56206_;
  assign new_n56208_ = ~\b[54]  & ~new_n56207_;
  assign new_n56209_ = ~new_n55347_ & new_n56051_;
  assign new_n56210_ = ~new_n56047_ & new_n56209_;
  assign new_n56211_ = ~new_n56048_ & ~new_n56051_;
  assign new_n56212_ = ~new_n56210_ & ~new_n56211_;
  assign new_n56213_ = ~new_n56116_ & ~new_n56212_;
  assign new_n56214_ = ~new_n55337_ & ~new_n56115_;
  assign new_n56215_ = ~new_n56114_ & new_n56214_;
  assign new_n56216_ = ~new_n56213_ & ~new_n56215_;
  assign new_n56217_ = ~\b[53]  & ~new_n56216_;
  assign new_n56218_ = ~new_n55356_ & new_n56046_;
  assign new_n56219_ = ~new_n56042_ & new_n56218_;
  assign new_n56220_ = ~new_n56043_ & ~new_n56046_;
  assign new_n56221_ = ~new_n56219_ & ~new_n56220_;
  assign new_n56222_ = ~new_n56116_ & ~new_n56221_;
  assign new_n56223_ = ~new_n55346_ & ~new_n56115_;
  assign new_n56224_ = ~new_n56114_ & new_n56223_;
  assign new_n56225_ = ~new_n56222_ & ~new_n56224_;
  assign new_n56226_ = ~\b[52]  & ~new_n56225_;
  assign new_n56227_ = ~new_n55365_ & new_n56041_;
  assign new_n56228_ = ~new_n56037_ & new_n56227_;
  assign new_n56229_ = ~new_n56038_ & ~new_n56041_;
  assign new_n56230_ = ~new_n56228_ & ~new_n56229_;
  assign new_n56231_ = ~new_n56116_ & ~new_n56230_;
  assign new_n56232_ = ~new_n55355_ & ~new_n56115_;
  assign new_n56233_ = ~new_n56114_ & new_n56232_;
  assign new_n56234_ = ~new_n56231_ & ~new_n56233_;
  assign new_n56235_ = ~\b[51]  & ~new_n56234_;
  assign new_n56236_ = ~new_n55374_ & new_n56036_;
  assign new_n56237_ = ~new_n56032_ & new_n56236_;
  assign new_n56238_ = ~new_n56033_ & ~new_n56036_;
  assign new_n56239_ = ~new_n56237_ & ~new_n56238_;
  assign new_n56240_ = ~new_n56116_ & ~new_n56239_;
  assign new_n56241_ = ~new_n55364_ & ~new_n56115_;
  assign new_n56242_ = ~new_n56114_ & new_n56241_;
  assign new_n56243_ = ~new_n56240_ & ~new_n56242_;
  assign new_n56244_ = ~\b[50]  & ~new_n56243_;
  assign new_n56245_ = ~new_n55383_ & new_n56031_;
  assign new_n56246_ = ~new_n56027_ & new_n56245_;
  assign new_n56247_ = ~new_n56028_ & ~new_n56031_;
  assign new_n56248_ = ~new_n56246_ & ~new_n56247_;
  assign new_n56249_ = ~new_n56116_ & ~new_n56248_;
  assign new_n56250_ = ~new_n55373_ & ~new_n56115_;
  assign new_n56251_ = ~new_n56114_ & new_n56250_;
  assign new_n56252_ = ~new_n56249_ & ~new_n56251_;
  assign new_n56253_ = ~\b[49]  & ~new_n56252_;
  assign new_n56254_ = ~new_n55392_ & new_n56026_;
  assign new_n56255_ = ~new_n56022_ & new_n56254_;
  assign new_n56256_ = ~new_n56023_ & ~new_n56026_;
  assign new_n56257_ = ~new_n56255_ & ~new_n56256_;
  assign new_n56258_ = ~new_n56116_ & ~new_n56257_;
  assign new_n56259_ = ~new_n55382_ & ~new_n56115_;
  assign new_n56260_ = ~new_n56114_ & new_n56259_;
  assign new_n56261_ = ~new_n56258_ & ~new_n56260_;
  assign new_n56262_ = ~\b[48]  & ~new_n56261_;
  assign new_n56263_ = ~new_n55401_ & new_n56021_;
  assign new_n56264_ = ~new_n56017_ & new_n56263_;
  assign new_n56265_ = ~new_n56018_ & ~new_n56021_;
  assign new_n56266_ = ~new_n56264_ & ~new_n56265_;
  assign new_n56267_ = ~new_n56116_ & ~new_n56266_;
  assign new_n56268_ = ~new_n55391_ & ~new_n56115_;
  assign new_n56269_ = ~new_n56114_ & new_n56268_;
  assign new_n56270_ = ~new_n56267_ & ~new_n56269_;
  assign new_n56271_ = ~\b[47]  & ~new_n56270_;
  assign new_n56272_ = ~new_n55410_ & new_n56016_;
  assign new_n56273_ = ~new_n56012_ & new_n56272_;
  assign new_n56274_ = ~new_n56013_ & ~new_n56016_;
  assign new_n56275_ = ~new_n56273_ & ~new_n56274_;
  assign new_n56276_ = ~new_n56116_ & ~new_n56275_;
  assign new_n56277_ = ~new_n55400_ & ~new_n56115_;
  assign new_n56278_ = ~new_n56114_ & new_n56277_;
  assign new_n56279_ = ~new_n56276_ & ~new_n56278_;
  assign new_n56280_ = ~\b[46]  & ~new_n56279_;
  assign new_n56281_ = ~new_n55419_ & new_n56011_;
  assign new_n56282_ = ~new_n56007_ & new_n56281_;
  assign new_n56283_ = ~new_n56008_ & ~new_n56011_;
  assign new_n56284_ = ~new_n56282_ & ~new_n56283_;
  assign new_n56285_ = ~new_n56116_ & ~new_n56284_;
  assign new_n56286_ = ~new_n55409_ & ~new_n56115_;
  assign new_n56287_ = ~new_n56114_ & new_n56286_;
  assign new_n56288_ = ~new_n56285_ & ~new_n56287_;
  assign new_n56289_ = ~\b[45]  & ~new_n56288_;
  assign new_n56290_ = ~new_n55428_ & new_n56006_;
  assign new_n56291_ = ~new_n56002_ & new_n56290_;
  assign new_n56292_ = ~new_n56003_ & ~new_n56006_;
  assign new_n56293_ = ~new_n56291_ & ~new_n56292_;
  assign new_n56294_ = ~new_n56116_ & ~new_n56293_;
  assign new_n56295_ = ~new_n55418_ & ~new_n56115_;
  assign new_n56296_ = ~new_n56114_ & new_n56295_;
  assign new_n56297_ = ~new_n56294_ & ~new_n56296_;
  assign new_n56298_ = ~\b[44]  & ~new_n56297_;
  assign new_n56299_ = ~new_n55437_ & new_n56001_;
  assign new_n56300_ = ~new_n55997_ & new_n56299_;
  assign new_n56301_ = ~new_n55998_ & ~new_n56001_;
  assign new_n56302_ = ~new_n56300_ & ~new_n56301_;
  assign new_n56303_ = ~new_n56116_ & ~new_n56302_;
  assign new_n56304_ = ~new_n55427_ & ~new_n56115_;
  assign new_n56305_ = ~new_n56114_ & new_n56304_;
  assign new_n56306_ = ~new_n56303_ & ~new_n56305_;
  assign new_n56307_ = ~\b[43]  & ~new_n56306_;
  assign new_n56308_ = ~new_n55446_ & new_n55996_;
  assign new_n56309_ = ~new_n55992_ & new_n56308_;
  assign new_n56310_ = ~new_n55993_ & ~new_n55996_;
  assign new_n56311_ = ~new_n56309_ & ~new_n56310_;
  assign new_n56312_ = ~new_n56116_ & ~new_n56311_;
  assign new_n56313_ = ~new_n55436_ & ~new_n56115_;
  assign new_n56314_ = ~new_n56114_ & new_n56313_;
  assign new_n56315_ = ~new_n56312_ & ~new_n56314_;
  assign new_n56316_ = ~\b[42]  & ~new_n56315_;
  assign new_n56317_ = ~new_n55455_ & new_n55991_;
  assign new_n56318_ = ~new_n55987_ & new_n56317_;
  assign new_n56319_ = ~new_n55988_ & ~new_n55991_;
  assign new_n56320_ = ~new_n56318_ & ~new_n56319_;
  assign new_n56321_ = ~new_n56116_ & ~new_n56320_;
  assign new_n56322_ = ~new_n55445_ & ~new_n56115_;
  assign new_n56323_ = ~new_n56114_ & new_n56322_;
  assign new_n56324_ = ~new_n56321_ & ~new_n56323_;
  assign new_n56325_ = ~\b[41]  & ~new_n56324_;
  assign new_n56326_ = ~new_n55464_ & new_n55986_;
  assign new_n56327_ = ~new_n55982_ & new_n56326_;
  assign new_n56328_ = ~new_n55983_ & ~new_n55986_;
  assign new_n56329_ = ~new_n56327_ & ~new_n56328_;
  assign new_n56330_ = ~new_n56116_ & ~new_n56329_;
  assign new_n56331_ = ~new_n55454_ & ~new_n56115_;
  assign new_n56332_ = ~new_n56114_ & new_n56331_;
  assign new_n56333_ = ~new_n56330_ & ~new_n56332_;
  assign new_n56334_ = ~\b[40]  & ~new_n56333_;
  assign new_n56335_ = ~new_n55473_ & new_n55981_;
  assign new_n56336_ = ~new_n55977_ & new_n56335_;
  assign new_n56337_ = ~new_n55978_ & ~new_n55981_;
  assign new_n56338_ = ~new_n56336_ & ~new_n56337_;
  assign new_n56339_ = ~new_n56116_ & ~new_n56338_;
  assign new_n56340_ = ~new_n55463_ & ~new_n56115_;
  assign new_n56341_ = ~new_n56114_ & new_n56340_;
  assign new_n56342_ = ~new_n56339_ & ~new_n56341_;
  assign new_n56343_ = ~\b[39]  & ~new_n56342_;
  assign new_n56344_ = ~new_n55482_ & new_n55976_;
  assign new_n56345_ = ~new_n55972_ & new_n56344_;
  assign new_n56346_ = ~new_n55973_ & ~new_n55976_;
  assign new_n56347_ = ~new_n56345_ & ~new_n56346_;
  assign new_n56348_ = ~new_n56116_ & ~new_n56347_;
  assign new_n56349_ = ~new_n55472_ & ~new_n56115_;
  assign new_n56350_ = ~new_n56114_ & new_n56349_;
  assign new_n56351_ = ~new_n56348_ & ~new_n56350_;
  assign new_n56352_ = ~\b[38]  & ~new_n56351_;
  assign new_n56353_ = ~new_n55491_ & new_n55971_;
  assign new_n56354_ = ~new_n55967_ & new_n56353_;
  assign new_n56355_ = ~new_n55968_ & ~new_n55971_;
  assign new_n56356_ = ~new_n56354_ & ~new_n56355_;
  assign new_n56357_ = ~new_n56116_ & ~new_n56356_;
  assign new_n56358_ = ~new_n55481_ & ~new_n56115_;
  assign new_n56359_ = ~new_n56114_ & new_n56358_;
  assign new_n56360_ = ~new_n56357_ & ~new_n56359_;
  assign new_n56361_ = ~\b[37]  & ~new_n56360_;
  assign new_n56362_ = ~new_n55500_ & new_n55966_;
  assign new_n56363_ = ~new_n55962_ & new_n56362_;
  assign new_n56364_ = ~new_n55963_ & ~new_n55966_;
  assign new_n56365_ = ~new_n56363_ & ~new_n56364_;
  assign new_n56366_ = ~new_n56116_ & ~new_n56365_;
  assign new_n56367_ = ~new_n55490_ & ~new_n56115_;
  assign new_n56368_ = ~new_n56114_ & new_n56367_;
  assign new_n56369_ = ~new_n56366_ & ~new_n56368_;
  assign new_n56370_ = ~\b[36]  & ~new_n56369_;
  assign new_n56371_ = ~new_n55509_ & new_n55961_;
  assign new_n56372_ = ~new_n55957_ & new_n56371_;
  assign new_n56373_ = ~new_n55958_ & ~new_n55961_;
  assign new_n56374_ = ~new_n56372_ & ~new_n56373_;
  assign new_n56375_ = ~new_n56116_ & ~new_n56374_;
  assign new_n56376_ = ~new_n55499_ & ~new_n56115_;
  assign new_n56377_ = ~new_n56114_ & new_n56376_;
  assign new_n56378_ = ~new_n56375_ & ~new_n56377_;
  assign new_n56379_ = ~\b[35]  & ~new_n56378_;
  assign new_n56380_ = ~new_n55518_ & new_n55956_;
  assign new_n56381_ = ~new_n55952_ & new_n56380_;
  assign new_n56382_ = ~new_n55953_ & ~new_n55956_;
  assign new_n56383_ = ~new_n56381_ & ~new_n56382_;
  assign new_n56384_ = ~new_n56116_ & ~new_n56383_;
  assign new_n56385_ = ~new_n55508_ & ~new_n56115_;
  assign new_n56386_ = ~new_n56114_ & new_n56385_;
  assign new_n56387_ = ~new_n56384_ & ~new_n56386_;
  assign new_n56388_ = ~\b[34]  & ~new_n56387_;
  assign new_n56389_ = ~new_n55527_ & new_n55951_;
  assign new_n56390_ = ~new_n55947_ & new_n56389_;
  assign new_n56391_ = ~new_n55948_ & ~new_n55951_;
  assign new_n56392_ = ~new_n56390_ & ~new_n56391_;
  assign new_n56393_ = ~new_n56116_ & ~new_n56392_;
  assign new_n56394_ = ~new_n55517_ & ~new_n56115_;
  assign new_n56395_ = ~new_n56114_ & new_n56394_;
  assign new_n56396_ = ~new_n56393_ & ~new_n56395_;
  assign new_n56397_ = ~\b[33]  & ~new_n56396_;
  assign new_n56398_ = ~new_n55536_ & new_n55946_;
  assign new_n56399_ = ~new_n55942_ & new_n56398_;
  assign new_n56400_ = ~new_n55943_ & ~new_n55946_;
  assign new_n56401_ = ~new_n56399_ & ~new_n56400_;
  assign new_n56402_ = ~new_n56116_ & ~new_n56401_;
  assign new_n56403_ = ~new_n55526_ & ~new_n56115_;
  assign new_n56404_ = ~new_n56114_ & new_n56403_;
  assign new_n56405_ = ~new_n56402_ & ~new_n56404_;
  assign new_n56406_ = ~\b[32]  & ~new_n56405_;
  assign new_n56407_ = ~new_n55545_ & new_n55941_;
  assign new_n56408_ = ~new_n55937_ & new_n56407_;
  assign new_n56409_ = ~new_n55938_ & ~new_n55941_;
  assign new_n56410_ = ~new_n56408_ & ~new_n56409_;
  assign new_n56411_ = ~new_n56116_ & ~new_n56410_;
  assign new_n56412_ = ~new_n55535_ & ~new_n56115_;
  assign new_n56413_ = ~new_n56114_ & new_n56412_;
  assign new_n56414_ = ~new_n56411_ & ~new_n56413_;
  assign new_n56415_ = ~\b[31]  & ~new_n56414_;
  assign new_n56416_ = ~new_n55554_ & new_n55936_;
  assign new_n56417_ = ~new_n55932_ & new_n56416_;
  assign new_n56418_ = ~new_n55933_ & ~new_n55936_;
  assign new_n56419_ = ~new_n56417_ & ~new_n56418_;
  assign new_n56420_ = ~new_n56116_ & ~new_n56419_;
  assign new_n56421_ = ~new_n55544_ & ~new_n56115_;
  assign new_n56422_ = ~new_n56114_ & new_n56421_;
  assign new_n56423_ = ~new_n56420_ & ~new_n56422_;
  assign new_n56424_ = ~\b[30]  & ~new_n56423_;
  assign new_n56425_ = ~new_n55563_ & new_n55931_;
  assign new_n56426_ = ~new_n55927_ & new_n56425_;
  assign new_n56427_ = ~new_n55928_ & ~new_n55931_;
  assign new_n56428_ = ~new_n56426_ & ~new_n56427_;
  assign new_n56429_ = ~new_n56116_ & ~new_n56428_;
  assign new_n56430_ = ~new_n55553_ & ~new_n56115_;
  assign new_n56431_ = ~new_n56114_ & new_n56430_;
  assign new_n56432_ = ~new_n56429_ & ~new_n56431_;
  assign new_n56433_ = ~\b[29]  & ~new_n56432_;
  assign new_n56434_ = ~new_n55572_ & new_n55926_;
  assign new_n56435_ = ~new_n55922_ & new_n56434_;
  assign new_n56436_ = ~new_n55923_ & ~new_n55926_;
  assign new_n56437_ = ~new_n56435_ & ~new_n56436_;
  assign new_n56438_ = ~new_n56116_ & ~new_n56437_;
  assign new_n56439_ = ~new_n55562_ & ~new_n56115_;
  assign new_n56440_ = ~new_n56114_ & new_n56439_;
  assign new_n56441_ = ~new_n56438_ & ~new_n56440_;
  assign new_n56442_ = ~\b[28]  & ~new_n56441_;
  assign new_n56443_ = ~new_n55581_ & new_n55921_;
  assign new_n56444_ = ~new_n55917_ & new_n56443_;
  assign new_n56445_ = ~new_n55918_ & ~new_n55921_;
  assign new_n56446_ = ~new_n56444_ & ~new_n56445_;
  assign new_n56447_ = ~new_n56116_ & ~new_n56446_;
  assign new_n56448_ = ~new_n55571_ & ~new_n56115_;
  assign new_n56449_ = ~new_n56114_ & new_n56448_;
  assign new_n56450_ = ~new_n56447_ & ~new_n56449_;
  assign new_n56451_ = ~\b[27]  & ~new_n56450_;
  assign new_n56452_ = ~new_n55590_ & new_n55916_;
  assign new_n56453_ = ~new_n55912_ & new_n56452_;
  assign new_n56454_ = ~new_n55913_ & ~new_n55916_;
  assign new_n56455_ = ~new_n56453_ & ~new_n56454_;
  assign new_n56456_ = ~new_n56116_ & ~new_n56455_;
  assign new_n56457_ = ~new_n55580_ & ~new_n56115_;
  assign new_n56458_ = ~new_n56114_ & new_n56457_;
  assign new_n56459_ = ~new_n56456_ & ~new_n56458_;
  assign new_n56460_ = ~\b[26]  & ~new_n56459_;
  assign new_n56461_ = ~new_n55599_ & new_n55911_;
  assign new_n56462_ = ~new_n55907_ & new_n56461_;
  assign new_n56463_ = ~new_n55908_ & ~new_n55911_;
  assign new_n56464_ = ~new_n56462_ & ~new_n56463_;
  assign new_n56465_ = ~new_n56116_ & ~new_n56464_;
  assign new_n56466_ = ~new_n55589_ & ~new_n56115_;
  assign new_n56467_ = ~new_n56114_ & new_n56466_;
  assign new_n56468_ = ~new_n56465_ & ~new_n56467_;
  assign new_n56469_ = ~\b[25]  & ~new_n56468_;
  assign new_n56470_ = ~new_n55608_ & new_n55906_;
  assign new_n56471_ = ~new_n55902_ & new_n56470_;
  assign new_n56472_ = ~new_n55903_ & ~new_n55906_;
  assign new_n56473_ = ~new_n56471_ & ~new_n56472_;
  assign new_n56474_ = ~new_n56116_ & ~new_n56473_;
  assign new_n56475_ = ~new_n55598_ & ~new_n56115_;
  assign new_n56476_ = ~new_n56114_ & new_n56475_;
  assign new_n56477_ = ~new_n56474_ & ~new_n56476_;
  assign new_n56478_ = ~\b[24]  & ~new_n56477_;
  assign new_n56479_ = ~new_n55617_ & new_n55901_;
  assign new_n56480_ = ~new_n55897_ & new_n56479_;
  assign new_n56481_ = ~new_n55898_ & ~new_n55901_;
  assign new_n56482_ = ~new_n56480_ & ~new_n56481_;
  assign new_n56483_ = ~new_n56116_ & ~new_n56482_;
  assign new_n56484_ = ~new_n55607_ & ~new_n56115_;
  assign new_n56485_ = ~new_n56114_ & new_n56484_;
  assign new_n56486_ = ~new_n56483_ & ~new_n56485_;
  assign new_n56487_ = ~\b[23]  & ~new_n56486_;
  assign new_n56488_ = ~new_n55626_ & new_n55896_;
  assign new_n56489_ = ~new_n55892_ & new_n56488_;
  assign new_n56490_ = ~new_n55893_ & ~new_n55896_;
  assign new_n56491_ = ~new_n56489_ & ~new_n56490_;
  assign new_n56492_ = ~new_n56116_ & ~new_n56491_;
  assign new_n56493_ = ~new_n55616_ & ~new_n56115_;
  assign new_n56494_ = ~new_n56114_ & new_n56493_;
  assign new_n56495_ = ~new_n56492_ & ~new_n56494_;
  assign new_n56496_ = ~\b[22]  & ~new_n56495_;
  assign new_n56497_ = ~new_n55635_ & new_n55891_;
  assign new_n56498_ = ~new_n55887_ & new_n56497_;
  assign new_n56499_ = ~new_n55888_ & ~new_n55891_;
  assign new_n56500_ = ~new_n56498_ & ~new_n56499_;
  assign new_n56501_ = ~new_n56116_ & ~new_n56500_;
  assign new_n56502_ = ~new_n55625_ & ~new_n56115_;
  assign new_n56503_ = ~new_n56114_ & new_n56502_;
  assign new_n56504_ = ~new_n56501_ & ~new_n56503_;
  assign new_n56505_ = ~\b[21]  & ~new_n56504_;
  assign new_n56506_ = ~new_n55644_ & new_n55886_;
  assign new_n56507_ = ~new_n55882_ & new_n56506_;
  assign new_n56508_ = ~new_n55883_ & ~new_n55886_;
  assign new_n56509_ = ~new_n56507_ & ~new_n56508_;
  assign new_n56510_ = ~new_n56116_ & ~new_n56509_;
  assign new_n56511_ = ~new_n55634_ & ~new_n56115_;
  assign new_n56512_ = ~new_n56114_ & new_n56511_;
  assign new_n56513_ = ~new_n56510_ & ~new_n56512_;
  assign new_n56514_ = ~\b[20]  & ~new_n56513_;
  assign new_n56515_ = ~new_n55653_ & new_n55881_;
  assign new_n56516_ = ~new_n55877_ & new_n56515_;
  assign new_n56517_ = ~new_n55878_ & ~new_n55881_;
  assign new_n56518_ = ~new_n56516_ & ~new_n56517_;
  assign new_n56519_ = ~new_n56116_ & ~new_n56518_;
  assign new_n56520_ = ~new_n55643_ & ~new_n56115_;
  assign new_n56521_ = ~new_n56114_ & new_n56520_;
  assign new_n56522_ = ~new_n56519_ & ~new_n56521_;
  assign new_n56523_ = ~\b[19]  & ~new_n56522_;
  assign new_n56524_ = ~new_n55662_ & new_n55876_;
  assign new_n56525_ = ~new_n55872_ & new_n56524_;
  assign new_n56526_ = ~new_n55873_ & ~new_n55876_;
  assign new_n56527_ = ~new_n56525_ & ~new_n56526_;
  assign new_n56528_ = ~new_n56116_ & ~new_n56527_;
  assign new_n56529_ = ~new_n55652_ & ~new_n56115_;
  assign new_n56530_ = ~new_n56114_ & new_n56529_;
  assign new_n56531_ = ~new_n56528_ & ~new_n56530_;
  assign new_n56532_ = ~\b[18]  & ~new_n56531_;
  assign new_n56533_ = ~new_n55671_ & new_n55871_;
  assign new_n56534_ = ~new_n55867_ & new_n56533_;
  assign new_n56535_ = ~new_n55868_ & ~new_n55871_;
  assign new_n56536_ = ~new_n56534_ & ~new_n56535_;
  assign new_n56537_ = ~new_n56116_ & ~new_n56536_;
  assign new_n56538_ = ~new_n55661_ & ~new_n56115_;
  assign new_n56539_ = ~new_n56114_ & new_n56538_;
  assign new_n56540_ = ~new_n56537_ & ~new_n56539_;
  assign new_n56541_ = ~\b[17]  & ~new_n56540_;
  assign new_n56542_ = ~new_n55680_ & new_n55866_;
  assign new_n56543_ = ~new_n55862_ & new_n56542_;
  assign new_n56544_ = ~new_n55863_ & ~new_n55866_;
  assign new_n56545_ = ~new_n56543_ & ~new_n56544_;
  assign new_n56546_ = ~new_n56116_ & ~new_n56545_;
  assign new_n56547_ = ~new_n55670_ & ~new_n56115_;
  assign new_n56548_ = ~new_n56114_ & new_n56547_;
  assign new_n56549_ = ~new_n56546_ & ~new_n56548_;
  assign new_n56550_ = ~\b[16]  & ~new_n56549_;
  assign new_n56551_ = ~new_n55689_ & new_n55861_;
  assign new_n56552_ = ~new_n55857_ & new_n56551_;
  assign new_n56553_ = ~new_n55858_ & ~new_n55861_;
  assign new_n56554_ = ~new_n56552_ & ~new_n56553_;
  assign new_n56555_ = ~new_n56116_ & ~new_n56554_;
  assign new_n56556_ = ~new_n55679_ & ~new_n56115_;
  assign new_n56557_ = ~new_n56114_ & new_n56556_;
  assign new_n56558_ = ~new_n56555_ & ~new_n56557_;
  assign new_n56559_ = ~\b[15]  & ~new_n56558_;
  assign new_n56560_ = ~new_n55698_ & new_n55856_;
  assign new_n56561_ = ~new_n55852_ & new_n56560_;
  assign new_n56562_ = ~new_n55853_ & ~new_n55856_;
  assign new_n56563_ = ~new_n56561_ & ~new_n56562_;
  assign new_n56564_ = ~new_n56116_ & ~new_n56563_;
  assign new_n56565_ = ~new_n55688_ & ~new_n56115_;
  assign new_n56566_ = ~new_n56114_ & new_n56565_;
  assign new_n56567_ = ~new_n56564_ & ~new_n56566_;
  assign new_n56568_ = ~\b[14]  & ~new_n56567_;
  assign new_n56569_ = ~new_n55707_ & new_n55851_;
  assign new_n56570_ = ~new_n55847_ & new_n56569_;
  assign new_n56571_ = ~new_n55848_ & ~new_n55851_;
  assign new_n56572_ = ~new_n56570_ & ~new_n56571_;
  assign new_n56573_ = ~new_n56116_ & ~new_n56572_;
  assign new_n56574_ = ~new_n55697_ & ~new_n56115_;
  assign new_n56575_ = ~new_n56114_ & new_n56574_;
  assign new_n56576_ = ~new_n56573_ & ~new_n56575_;
  assign new_n56577_ = ~\b[13]  & ~new_n56576_;
  assign new_n56578_ = ~new_n55716_ & new_n55846_;
  assign new_n56579_ = ~new_n55842_ & new_n56578_;
  assign new_n56580_ = ~new_n55843_ & ~new_n55846_;
  assign new_n56581_ = ~new_n56579_ & ~new_n56580_;
  assign new_n56582_ = ~new_n56116_ & ~new_n56581_;
  assign new_n56583_ = ~new_n55706_ & ~new_n56115_;
  assign new_n56584_ = ~new_n56114_ & new_n56583_;
  assign new_n56585_ = ~new_n56582_ & ~new_n56584_;
  assign new_n56586_ = ~\b[12]  & ~new_n56585_;
  assign new_n56587_ = ~new_n55725_ & new_n55841_;
  assign new_n56588_ = ~new_n55837_ & new_n56587_;
  assign new_n56589_ = ~new_n55838_ & ~new_n55841_;
  assign new_n56590_ = ~new_n56588_ & ~new_n56589_;
  assign new_n56591_ = ~new_n56116_ & ~new_n56590_;
  assign new_n56592_ = ~new_n55715_ & ~new_n56115_;
  assign new_n56593_ = ~new_n56114_ & new_n56592_;
  assign new_n56594_ = ~new_n56591_ & ~new_n56593_;
  assign new_n56595_ = ~\b[11]  & ~new_n56594_;
  assign new_n56596_ = ~new_n55734_ & new_n55836_;
  assign new_n56597_ = ~new_n55832_ & new_n56596_;
  assign new_n56598_ = ~new_n55833_ & ~new_n55836_;
  assign new_n56599_ = ~new_n56597_ & ~new_n56598_;
  assign new_n56600_ = ~new_n56116_ & ~new_n56599_;
  assign new_n56601_ = ~new_n55724_ & ~new_n56115_;
  assign new_n56602_ = ~new_n56114_ & new_n56601_;
  assign new_n56603_ = ~new_n56600_ & ~new_n56602_;
  assign new_n56604_ = ~\b[10]  & ~new_n56603_;
  assign new_n56605_ = ~new_n55743_ & new_n55831_;
  assign new_n56606_ = ~new_n55827_ & new_n56605_;
  assign new_n56607_ = ~new_n55828_ & ~new_n55831_;
  assign new_n56608_ = ~new_n56606_ & ~new_n56607_;
  assign new_n56609_ = ~new_n56116_ & ~new_n56608_;
  assign new_n56610_ = ~new_n55733_ & ~new_n56115_;
  assign new_n56611_ = ~new_n56114_ & new_n56610_;
  assign new_n56612_ = ~new_n56609_ & ~new_n56611_;
  assign new_n56613_ = ~\b[9]  & ~new_n56612_;
  assign new_n56614_ = ~new_n55752_ & new_n55826_;
  assign new_n56615_ = ~new_n55822_ & new_n56614_;
  assign new_n56616_ = ~new_n55823_ & ~new_n55826_;
  assign new_n56617_ = ~new_n56615_ & ~new_n56616_;
  assign new_n56618_ = ~new_n56116_ & ~new_n56617_;
  assign new_n56619_ = ~new_n55742_ & ~new_n56115_;
  assign new_n56620_ = ~new_n56114_ & new_n56619_;
  assign new_n56621_ = ~new_n56618_ & ~new_n56620_;
  assign new_n56622_ = ~\b[8]  & ~new_n56621_;
  assign new_n56623_ = ~new_n55761_ & new_n55821_;
  assign new_n56624_ = ~new_n55817_ & new_n56623_;
  assign new_n56625_ = ~new_n55818_ & ~new_n55821_;
  assign new_n56626_ = ~new_n56624_ & ~new_n56625_;
  assign new_n56627_ = ~new_n56116_ & ~new_n56626_;
  assign new_n56628_ = ~new_n55751_ & ~new_n56115_;
  assign new_n56629_ = ~new_n56114_ & new_n56628_;
  assign new_n56630_ = ~new_n56627_ & ~new_n56629_;
  assign new_n56631_ = ~\b[7]  & ~new_n56630_;
  assign new_n56632_ = ~new_n55770_ & new_n55816_;
  assign new_n56633_ = ~new_n55812_ & new_n56632_;
  assign new_n56634_ = ~new_n55813_ & ~new_n55816_;
  assign new_n56635_ = ~new_n56633_ & ~new_n56634_;
  assign new_n56636_ = ~new_n56116_ & ~new_n56635_;
  assign new_n56637_ = ~new_n55760_ & ~new_n56115_;
  assign new_n56638_ = ~new_n56114_ & new_n56637_;
  assign new_n56639_ = ~new_n56636_ & ~new_n56638_;
  assign new_n56640_ = ~\b[6]  & ~new_n56639_;
  assign new_n56641_ = ~new_n55779_ & new_n55811_;
  assign new_n56642_ = ~new_n55807_ & new_n56641_;
  assign new_n56643_ = ~new_n55808_ & ~new_n55811_;
  assign new_n56644_ = ~new_n56642_ & ~new_n56643_;
  assign new_n56645_ = ~new_n56116_ & ~new_n56644_;
  assign new_n56646_ = ~new_n55769_ & ~new_n56115_;
  assign new_n56647_ = ~new_n56114_ & new_n56646_;
  assign new_n56648_ = ~new_n56645_ & ~new_n56647_;
  assign new_n56649_ = ~\b[5]  & ~new_n56648_;
  assign new_n56650_ = ~new_n55787_ & new_n55806_;
  assign new_n56651_ = ~new_n55802_ & new_n56650_;
  assign new_n56652_ = ~new_n55803_ & ~new_n55806_;
  assign new_n56653_ = ~new_n56651_ & ~new_n56652_;
  assign new_n56654_ = ~new_n56116_ & ~new_n56653_;
  assign new_n56655_ = ~new_n55778_ & ~new_n56115_;
  assign new_n56656_ = ~new_n56114_ & new_n56655_;
  assign new_n56657_ = ~new_n56654_ & ~new_n56656_;
  assign new_n56658_ = ~\b[4]  & ~new_n56657_;
  assign new_n56659_ = ~new_n55797_ & new_n55801_;
  assign new_n56660_ = ~new_n55796_ & new_n56659_;
  assign new_n56661_ = ~new_n55798_ & ~new_n55801_;
  assign new_n56662_ = ~new_n56660_ & ~new_n56661_;
  assign new_n56663_ = ~new_n56116_ & ~new_n56662_;
  assign new_n56664_ = ~new_n55786_ & ~new_n56115_;
  assign new_n56665_ = ~new_n56114_ & new_n56664_;
  assign new_n56666_ = ~new_n56663_ & ~new_n56665_;
  assign new_n56667_ = ~\b[3]  & ~new_n56666_;
  assign new_n56668_ = new_n27783_ & ~new_n55794_;
  assign new_n56669_ = ~new_n55792_ & new_n56668_;
  assign new_n56670_ = ~new_n55796_ & ~new_n56669_;
  assign new_n56671_ = ~new_n56116_ & new_n56670_;
  assign new_n56672_ = ~new_n55791_ & ~new_n56115_;
  assign new_n56673_ = ~new_n56114_ & new_n56672_;
  assign new_n56674_ = ~new_n56671_ & ~new_n56673_;
  assign new_n56675_ = ~\b[2]  & ~new_n56674_;
  assign new_n56676_ = \b[0]  & ~new_n56116_;
  assign new_n56677_ = \a[1]  & ~new_n56676_;
  assign new_n56678_ = new_n27783_ & ~new_n56116_;
  assign new_n56679_ = ~new_n56677_ & ~new_n56678_;
  assign new_n56680_ = \b[1]  & ~new_n56679_;
  assign new_n56681_ = ~\b[1]  & ~new_n56678_;
  assign new_n56682_ = ~new_n56677_ & new_n56681_;
  assign new_n56683_ = ~new_n56680_ & ~new_n56682_;
  assign new_n56684_ = ~new_n28345_ & ~new_n56683_;
  assign new_n56685_ = ~\b[1]  & ~new_n56679_;
  assign new_n56686_ = ~new_n56684_ & ~new_n56685_;
  assign new_n56687_ = \b[2]  & ~new_n56673_;
  assign new_n56688_ = ~new_n56671_ & new_n56687_;
  assign new_n56689_ = ~new_n56675_ & ~new_n56688_;
  assign new_n56690_ = ~new_n56686_ & new_n56689_;
  assign new_n56691_ = ~new_n56675_ & ~new_n56690_;
  assign new_n56692_ = \b[3]  & ~new_n56665_;
  assign new_n56693_ = ~new_n56663_ & new_n56692_;
  assign new_n56694_ = ~new_n56667_ & ~new_n56693_;
  assign new_n56695_ = ~new_n56691_ & new_n56694_;
  assign new_n56696_ = ~new_n56667_ & ~new_n56695_;
  assign new_n56697_ = \b[4]  & ~new_n56656_;
  assign new_n56698_ = ~new_n56654_ & new_n56697_;
  assign new_n56699_ = ~new_n56658_ & ~new_n56698_;
  assign new_n56700_ = ~new_n56696_ & new_n56699_;
  assign new_n56701_ = ~new_n56658_ & ~new_n56700_;
  assign new_n56702_ = \b[5]  & ~new_n56647_;
  assign new_n56703_ = ~new_n56645_ & new_n56702_;
  assign new_n56704_ = ~new_n56649_ & ~new_n56703_;
  assign new_n56705_ = ~new_n56701_ & new_n56704_;
  assign new_n56706_ = ~new_n56649_ & ~new_n56705_;
  assign new_n56707_ = \b[6]  & ~new_n56638_;
  assign new_n56708_ = ~new_n56636_ & new_n56707_;
  assign new_n56709_ = ~new_n56640_ & ~new_n56708_;
  assign new_n56710_ = ~new_n56706_ & new_n56709_;
  assign new_n56711_ = ~new_n56640_ & ~new_n56710_;
  assign new_n56712_ = \b[7]  & ~new_n56629_;
  assign new_n56713_ = ~new_n56627_ & new_n56712_;
  assign new_n56714_ = ~new_n56631_ & ~new_n56713_;
  assign new_n56715_ = ~new_n56711_ & new_n56714_;
  assign new_n56716_ = ~new_n56631_ & ~new_n56715_;
  assign new_n56717_ = \b[8]  & ~new_n56620_;
  assign new_n56718_ = ~new_n56618_ & new_n56717_;
  assign new_n56719_ = ~new_n56622_ & ~new_n56718_;
  assign new_n56720_ = ~new_n56716_ & new_n56719_;
  assign new_n56721_ = ~new_n56622_ & ~new_n56720_;
  assign new_n56722_ = \b[9]  & ~new_n56611_;
  assign new_n56723_ = ~new_n56609_ & new_n56722_;
  assign new_n56724_ = ~new_n56613_ & ~new_n56723_;
  assign new_n56725_ = ~new_n56721_ & new_n56724_;
  assign new_n56726_ = ~new_n56613_ & ~new_n56725_;
  assign new_n56727_ = \b[10]  & ~new_n56602_;
  assign new_n56728_ = ~new_n56600_ & new_n56727_;
  assign new_n56729_ = ~new_n56604_ & ~new_n56728_;
  assign new_n56730_ = ~new_n56726_ & new_n56729_;
  assign new_n56731_ = ~new_n56604_ & ~new_n56730_;
  assign new_n56732_ = \b[11]  & ~new_n56593_;
  assign new_n56733_ = ~new_n56591_ & new_n56732_;
  assign new_n56734_ = ~new_n56595_ & ~new_n56733_;
  assign new_n56735_ = ~new_n56731_ & new_n56734_;
  assign new_n56736_ = ~new_n56595_ & ~new_n56735_;
  assign new_n56737_ = \b[12]  & ~new_n56584_;
  assign new_n56738_ = ~new_n56582_ & new_n56737_;
  assign new_n56739_ = ~new_n56586_ & ~new_n56738_;
  assign new_n56740_ = ~new_n56736_ & new_n56739_;
  assign new_n56741_ = ~new_n56586_ & ~new_n56740_;
  assign new_n56742_ = \b[13]  & ~new_n56575_;
  assign new_n56743_ = ~new_n56573_ & new_n56742_;
  assign new_n56744_ = ~new_n56577_ & ~new_n56743_;
  assign new_n56745_ = ~new_n56741_ & new_n56744_;
  assign new_n56746_ = ~new_n56577_ & ~new_n56745_;
  assign new_n56747_ = \b[14]  & ~new_n56566_;
  assign new_n56748_ = ~new_n56564_ & new_n56747_;
  assign new_n56749_ = ~new_n56568_ & ~new_n56748_;
  assign new_n56750_ = ~new_n56746_ & new_n56749_;
  assign new_n56751_ = ~new_n56568_ & ~new_n56750_;
  assign new_n56752_ = \b[15]  & ~new_n56557_;
  assign new_n56753_ = ~new_n56555_ & new_n56752_;
  assign new_n56754_ = ~new_n56559_ & ~new_n56753_;
  assign new_n56755_ = ~new_n56751_ & new_n56754_;
  assign new_n56756_ = ~new_n56559_ & ~new_n56755_;
  assign new_n56757_ = \b[16]  & ~new_n56548_;
  assign new_n56758_ = ~new_n56546_ & new_n56757_;
  assign new_n56759_ = ~new_n56550_ & ~new_n56758_;
  assign new_n56760_ = ~new_n56756_ & new_n56759_;
  assign new_n56761_ = ~new_n56550_ & ~new_n56760_;
  assign new_n56762_ = \b[17]  & ~new_n56539_;
  assign new_n56763_ = ~new_n56537_ & new_n56762_;
  assign new_n56764_ = ~new_n56541_ & ~new_n56763_;
  assign new_n56765_ = ~new_n56761_ & new_n56764_;
  assign new_n56766_ = ~new_n56541_ & ~new_n56765_;
  assign new_n56767_ = \b[18]  & ~new_n56530_;
  assign new_n56768_ = ~new_n56528_ & new_n56767_;
  assign new_n56769_ = ~new_n56532_ & ~new_n56768_;
  assign new_n56770_ = ~new_n56766_ & new_n56769_;
  assign new_n56771_ = ~new_n56532_ & ~new_n56770_;
  assign new_n56772_ = \b[19]  & ~new_n56521_;
  assign new_n56773_ = ~new_n56519_ & new_n56772_;
  assign new_n56774_ = ~new_n56523_ & ~new_n56773_;
  assign new_n56775_ = ~new_n56771_ & new_n56774_;
  assign new_n56776_ = ~new_n56523_ & ~new_n56775_;
  assign new_n56777_ = \b[20]  & ~new_n56512_;
  assign new_n56778_ = ~new_n56510_ & new_n56777_;
  assign new_n56779_ = ~new_n56514_ & ~new_n56778_;
  assign new_n56780_ = ~new_n56776_ & new_n56779_;
  assign new_n56781_ = ~new_n56514_ & ~new_n56780_;
  assign new_n56782_ = \b[21]  & ~new_n56503_;
  assign new_n56783_ = ~new_n56501_ & new_n56782_;
  assign new_n56784_ = ~new_n56505_ & ~new_n56783_;
  assign new_n56785_ = ~new_n56781_ & new_n56784_;
  assign new_n56786_ = ~new_n56505_ & ~new_n56785_;
  assign new_n56787_ = \b[22]  & ~new_n56494_;
  assign new_n56788_ = ~new_n56492_ & new_n56787_;
  assign new_n56789_ = ~new_n56496_ & ~new_n56788_;
  assign new_n56790_ = ~new_n56786_ & new_n56789_;
  assign new_n56791_ = ~new_n56496_ & ~new_n56790_;
  assign new_n56792_ = \b[23]  & ~new_n56485_;
  assign new_n56793_ = ~new_n56483_ & new_n56792_;
  assign new_n56794_ = ~new_n56487_ & ~new_n56793_;
  assign new_n56795_ = ~new_n56791_ & new_n56794_;
  assign new_n56796_ = ~new_n56487_ & ~new_n56795_;
  assign new_n56797_ = \b[24]  & ~new_n56476_;
  assign new_n56798_ = ~new_n56474_ & new_n56797_;
  assign new_n56799_ = ~new_n56478_ & ~new_n56798_;
  assign new_n56800_ = ~new_n56796_ & new_n56799_;
  assign new_n56801_ = ~new_n56478_ & ~new_n56800_;
  assign new_n56802_ = \b[25]  & ~new_n56467_;
  assign new_n56803_ = ~new_n56465_ & new_n56802_;
  assign new_n56804_ = ~new_n56469_ & ~new_n56803_;
  assign new_n56805_ = ~new_n56801_ & new_n56804_;
  assign new_n56806_ = ~new_n56469_ & ~new_n56805_;
  assign new_n56807_ = \b[26]  & ~new_n56458_;
  assign new_n56808_ = ~new_n56456_ & new_n56807_;
  assign new_n56809_ = ~new_n56460_ & ~new_n56808_;
  assign new_n56810_ = ~new_n56806_ & new_n56809_;
  assign new_n56811_ = ~new_n56460_ & ~new_n56810_;
  assign new_n56812_ = \b[27]  & ~new_n56449_;
  assign new_n56813_ = ~new_n56447_ & new_n56812_;
  assign new_n56814_ = ~new_n56451_ & ~new_n56813_;
  assign new_n56815_ = ~new_n56811_ & new_n56814_;
  assign new_n56816_ = ~new_n56451_ & ~new_n56815_;
  assign new_n56817_ = \b[28]  & ~new_n56440_;
  assign new_n56818_ = ~new_n56438_ & new_n56817_;
  assign new_n56819_ = ~new_n56442_ & ~new_n56818_;
  assign new_n56820_ = ~new_n56816_ & new_n56819_;
  assign new_n56821_ = ~new_n56442_ & ~new_n56820_;
  assign new_n56822_ = \b[29]  & ~new_n56431_;
  assign new_n56823_ = ~new_n56429_ & new_n56822_;
  assign new_n56824_ = ~new_n56433_ & ~new_n56823_;
  assign new_n56825_ = ~new_n56821_ & new_n56824_;
  assign new_n56826_ = ~new_n56433_ & ~new_n56825_;
  assign new_n56827_ = \b[30]  & ~new_n56422_;
  assign new_n56828_ = ~new_n56420_ & new_n56827_;
  assign new_n56829_ = ~new_n56424_ & ~new_n56828_;
  assign new_n56830_ = ~new_n56826_ & new_n56829_;
  assign new_n56831_ = ~new_n56424_ & ~new_n56830_;
  assign new_n56832_ = \b[31]  & ~new_n56413_;
  assign new_n56833_ = ~new_n56411_ & new_n56832_;
  assign new_n56834_ = ~new_n56415_ & ~new_n56833_;
  assign new_n56835_ = ~new_n56831_ & new_n56834_;
  assign new_n56836_ = ~new_n56415_ & ~new_n56835_;
  assign new_n56837_ = \b[32]  & ~new_n56404_;
  assign new_n56838_ = ~new_n56402_ & new_n56837_;
  assign new_n56839_ = ~new_n56406_ & ~new_n56838_;
  assign new_n56840_ = ~new_n56836_ & new_n56839_;
  assign new_n56841_ = ~new_n56406_ & ~new_n56840_;
  assign new_n56842_ = \b[33]  & ~new_n56395_;
  assign new_n56843_ = ~new_n56393_ & new_n56842_;
  assign new_n56844_ = ~new_n56397_ & ~new_n56843_;
  assign new_n56845_ = ~new_n56841_ & new_n56844_;
  assign new_n56846_ = ~new_n56397_ & ~new_n56845_;
  assign new_n56847_ = \b[34]  & ~new_n56386_;
  assign new_n56848_ = ~new_n56384_ & new_n56847_;
  assign new_n56849_ = ~new_n56388_ & ~new_n56848_;
  assign new_n56850_ = ~new_n56846_ & new_n56849_;
  assign new_n56851_ = ~new_n56388_ & ~new_n56850_;
  assign new_n56852_ = \b[35]  & ~new_n56377_;
  assign new_n56853_ = ~new_n56375_ & new_n56852_;
  assign new_n56854_ = ~new_n56379_ & ~new_n56853_;
  assign new_n56855_ = ~new_n56851_ & new_n56854_;
  assign new_n56856_ = ~new_n56379_ & ~new_n56855_;
  assign new_n56857_ = \b[36]  & ~new_n56368_;
  assign new_n56858_ = ~new_n56366_ & new_n56857_;
  assign new_n56859_ = ~new_n56370_ & ~new_n56858_;
  assign new_n56860_ = ~new_n56856_ & new_n56859_;
  assign new_n56861_ = ~new_n56370_ & ~new_n56860_;
  assign new_n56862_ = \b[37]  & ~new_n56359_;
  assign new_n56863_ = ~new_n56357_ & new_n56862_;
  assign new_n56864_ = ~new_n56361_ & ~new_n56863_;
  assign new_n56865_ = ~new_n56861_ & new_n56864_;
  assign new_n56866_ = ~new_n56361_ & ~new_n56865_;
  assign new_n56867_ = \b[38]  & ~new_n56350_;
  assign new_n56868_ = ~new_n56348_ & new_n56867_;
  assign new_n56869_ = ~new_n56352_ & ~new_n56868_;
  assign new_n56870_ = ~new_n56866_ & new_n56869_;
  assign new_n56871_ = ~new_n56352_ & ~new_n56870_;
  assign new_n56872_ = \b[39]  & ~new_n56341_;
  assign new_n56873_ = ~new_n56339_ & new_n56872_;
  assign new_n56874_ = ~new_n56343_ & ~new_n56873_;
  assign new_n56875_ = ~new_n56871_ & new_n56874_;
  assign new_n56876_ = ~new_n56343_ & ~new_n56875_;
  assign new_n56877_ = \b[40]  & ~new_n56332_;
  assign new_n56878_ = ~new_n56330_ & new_n56877_;
  assign new_n56879_ = ~new_n56334_ & ~new_n56878_;
  assign new_n56880_ = ~new_n56876_ & new_n56879_;
  assign new_n56881_ = ~new_n56334_ & ~new_n56880_;
  assign new_n56882_ = \b[41]  & ~new_n56323_;
  assign new_n56883_ = ~new_n56321_ & new_n56882_;
  assign new_n56884_ = ~new_n56325_ & ~new_n56883_;
  assign new_n56885_ = ~new_n56881_ & new_n56884_;
  assign new_n56886_ = ~new_n56325_ & ~new_n56885_;
  assign new_n56887_ = \b[42]  & ~new_n56314_;
  assign new_n56888_ = ~new_n56312_ & new_n56887_;
  assign new_n56889_ = ~new_n56316_ & ~new_n56888_;
  assign new_n56890_ = ~new_n56886_ & new_n56889_;
  assign new_n56891_ = ~new_n56316_ & ~new_n56890_;
  assign new_n56892_ = \b[43]  & ~new_n56305_;
  assign new_n56893_ = ~new_n56303_ & new_n56892_;
  assign new_n56894_ = ~new_n56307_ & ~new_n56893_;
  assign new_n56895_ = ~new_n56891_ & new_n56894_;
  assign new_n56896_ = ~new_n56307_ & ~new_n56895_;
  assign new_n56897_ = \b[44]  & ~new_n56296_;
  assign new_n56898_ = ~new_n56294_ & new_n56897_;
  assign new_n56899_ = ~new_n56298_ & ~new_n56898_;
  assign new_n56900_ = ~new_n56896_ & new_n56899_;
  assign new_n56901_ = ~new_n56298_ & ~new_n56900_;
  assign new_n56902_ = \b[45]  & ~new_n56287_;
  assign new_n56903_ = ~new_n56285_ & new_n56902_;
  assign new_n56904_ = ~new_n56289_ & ~new_n56903_;
  assign new_n56905_ = ~new_n56901_ & new_n56904_;
  assign new_n56906_ = ~new_n56289_ & ~new_n56905_;
  assign new_n56907_ = \b[46]  & ~new_n56278_;
  assign new_n56908_ = ~new_n56276_ & new_n56907_;
  assign new_n56909_ = ~new_n56280_ & ~new_n56908_;
  assign new_n56910_ = ~new_n56906_ & new_n56909_;
  assign new_n56911_ = ~new_n56280_ & ~new_n56910_;
  assign new_n56912_ = \b[47]  & ~new_n56269_;
  assign new_n56913_ = ~new_n56267_ & new_n56912_;
  assign new_n56914_ = ~new_n56271_ & ~new_n56913_;
  assign new_n56915_ = ~new_n56911_ & new_n56914_;
  assign new_n56916_ = ~new_n56271_ & ~new_n56915_;
  assign new_n56917_ = \b[48]  & ~new_n56260_;
  assign new_n56918_ = ~new_n56258_ & new_n56917_;
  assign new_n56919_ = ~new_n56262_ & ~new_n56918_;
  assign new_n56920_ = ~new_n56916_ & new_n56919_;
  assign new_n56921_ = ~new_n56262_ & ~new_n56920_;
  assign new_n56922_ = \b[49]  & ~new_n56251_;
  assign new_n56923_ = ~new_n56249_ & new_n56922_;
  assign new_n56924_ = ~new_n56253_ & ~new_n56923_;
  assign new_n56925_ = ~new_n56921_ & new_n56924_;
  assign new_n56926_ = ~new_n56253_ & ~new_n56925_;
  assign new_n56927_ = \b[50]  & ~new_n56242_;
  assign new_n56928_ = ~new_n56240_ & new_n56927_;
  assign new_n56929_ = ~new_n56244_ & ~new_n56928_;
  assign new_n56930_ = ~new_n56926_ & new_n56929_;
  assign new_n56931_ = ~new_n56244_ & ~new_n56930_;
  assign new_n56932_ = \b[51]  & ~new_n56233_;
  assign new_n56933_ = ~new_n56231_ & new_n56932_;
  assign new_n56934_ = ~new_n56235_ & ~new_n56933_;
  assign new_n56935_ = ~new_n56931_ & new_n56934_;
  assign new_n56936_ = ~new_n56235_ & ~new_n56935_;
  assign new_n56937_ = \b[52]  & ~new_n56224_;
  assign new_n56938_ = ~new_n56222_ & new_n56937_;
  assign new_n56939_ = ~new_n56226_ & ~new_n56938_;
  assign new_n56940_ = ~new_n56936_ & new_n56939_;
  assign new_n56941_ = ~new_n56226_ & ~new_n56940_;
  assign new_n56942_ = \b[53]  & ~new_n56215_;
  assign new_n56943_ = ~new_n56213_ & new_n56942_;
  assign new_n56944_ = ~new_n56217_ & ~new_n56943_;
  assign new_n56945_ = ~new_n56941_ & new_n56944_;
  assign new_n56946_ = ~new_n56217_ & ~new_n56945_;
  assign new_n56947_ = \b[54]  & ~new_n56206_;
  assign new_n56948_ = ~new_n56204_ & new_n56947_;
  assign new_n56949_ = ~new_n56208_ & ~new_n56948_;
  assign new_n56950_ = ~new_n56946_ & new_n56949_;
  assign new_n56951_ = ~new_n56208_ & ~new_n56950_;
  assign new_n56952_ = \b[55]  & ~new_n56197_;
  assign new_n56953_ = ~new_n56195_ & new_n56952_;
  assign new_n56954_ = ~new_n56199_ & ~new_n56953_;
  assign new_n56955_ = ~new_n56951_ & new_n56954_;
  assign new_n56956_ = ~new_n56199_ & ~new_n56955_;
  assign new_n56957_ = \b[56]  & ~new_n56188_;
  assign new_n56958_ = ~new_n56186_ & new_n56957_;
  assign new_n56959_ = ~new_n56190_ & ~new_n56958_;
  assign new_n56960_ = ~new_n56956_ & new_n56959_;
  assign new_n56961_ = ~new_n56190_ & ~new_n56960_;
  assign new_n56962_ = \b[57]  & ~new_n56179_;
  assign new_n56963_ = ~new_n56177_ & new_n56962_;
  assign new_n56964_ = ~new_n56181_ & ~new_n56963_;
  assign new_n56965_ = ~new_n56961_ & new_n56964_;
  assign new_n56966_ = ~new_n56181_ & ~new_n56965_;
  assign new_n56967_ = \b[58]  & ~new_n56170_;
  assign new_n56968_ = ~new_n56168_ & new_n56967_;
  assign new_n56969_ = ~new_n56172_ & ~new_n56968_;
  assign new_n56970_ = ~new_n56966_ & new_n56969_;
  assign new_n56971_ = ~new_n56172_ & ~new_n56970_;
  assign new_n56972_ = \b[59]  & ~new_n56161_;
  assign new_n56973_ = ~new_n56159_ & new_n56972_;
  assign new_n56974_ = ~new_n56163_ & ~new_n56973_;
  assign new_n56975_ = ~new_n56971_ & new_n56974_;
  assign new_n56976_ = ~new_n56163_ & ~new_n56975_;
  assign new_n56977_ = \b[60]  & ~new_n56152_;
  assign new_n56978_ = ~new_n56150_ & new_n56977_;
  assign new_n56979_ = ~new_n56154_ & ~new_n56978_;
  assign new_n56980_ = ~new_n56976_ & new_n56979_;
  assign new_n56981_ = ~new_n56154_ & ~new_n56980_;
  assign new_n56982_ = \b[61]  & ~new_n56143_;
  assign new_n56983_ = ~new_n56141_ & new_n56982_;
  assign new_n56984_ = ~new_n56145_ & ~new_n56983_;
  assign new_n56985_ = ~new_n56981_ & new_n56984_;
  assign new_n56986_ = ~new_n56145_ & ~new_n56985_;
  assign new_n56987_ = \b[62]  & ~new_n56134_;
  assign new_n56988_ = ~new_n56132_ & new_n56987_;
  assign new_n56989_ = ~new_n56136_ & ~new_n56988_;
  assign new_n56990_ = ~new_n56986_ & new_n56989_;
  assign new_n56991_ = ~new_n56136_ & ~new_n56990_;
  assign new_n56992_ = \b[63]  & ~new_n56125_;
  assign new_n56993_ = ~new_n56123_ & new_n56992_;
  assign new_n56994_ = ~new_n56127_ & ~new_n56993_;
  assign new_n56995_ = ~new_n56991_ & new_n56994_;
  assign new_n56996_ = ~new_n56127_ & ~new_n56995_;
  assign new_n56997_ = \b[0]  & ~new_n56996_;
  assign new_n56998_ = \a[0]  & ~new_n56997_;
  assign new_n56999_ = new_n28345_ & ~new_n56996_;
  assign \remainder[0]  = new_n56998_ | new_n56999_;
  assign new_n57001_ = new_n28345_ & ~new_n56682_;
  assign new_n57002_ = ~new_n56680_ & new_n57001_;
  assign new_n57003_ = ~new_n56684_ & ~new_n57002_;
  assign new_n57004_ = ~new_n56996_ & new_n57003_;
  assign new_n57005_ = ~new_n56127_ & ~new_n56679_;
  assign new_n57006_ = ~new_n56995_ & new_n57005_;
  assign \remainder[1]  = new_n57004_ | new_n57006_;
  assign new_n57008_ = ~new_n56685_ & new_n56689_;
  assign new_n57009_ = ~new_n56684_ & new_n57008_;
  assign new_n57010_ = ~new_n56686_ & ~new_n56689_;
  assign new_n57011_ = ~new_n57009_ & ~new_n57010_;
  assign new_n57012_ = ~new_n56996_ & ~new_n57011_;
  assign new_n57013_ = ~new_n56127_ & ~new_n56674_;
  assign new_n57014_ = ~new_n56995_ & new_n57013_;
  assign \remainder[2]  = new_n57012_ | new_n57014_;
  assign new_n57016_ = ~new_n56675_ & new_n56694_;
  assign new_n57017_ = ~new_n56690_ & new_n57016_;
  assign new_n57018_ = ~new_n56691_ & ~new_n56694_;
  assign new_n57019_ = ~new_n57017_ & ~new_n57018_;
  assign new_n57020_ = ~new_n56996_ & ~new_n57019_;
  assign new_n57021_ = ~new_n56127_ & ~new_n56666_;
  assign new_n57022_ = ~new_n56995_ & new_n57021_;
  assign \remainder[3]  = new_n57020_ | new_n57022_;
  assign new_n57024_ = ~new_n56667_ & new_n56699_;
  assign new_n57025_ = ~new_n56695_ & new_n57024_;
  assign new_n57026_ = ~new_n56696_ & ~new_n56699_;
  assign new_n57027_ = ~new_n57025_ & ~new_n57026_;
  assign new_n57028_ = ~new_n56996_ & ~new_n57027_;
  assign new_n57029_ = ~new_n56127_ & ~new_n56657_;
  assign new_n57030_ = ~new_n56995_ & new_n57029_;
  assign \remainder[4]  = new_n57028_ | new_n57030_;
  assign new_n57032_ = ~new_n56658_ & new_n56704_;
  assign new_n57033_ = ~new_n56700_ & new_n57032_;
  assign new_n57034_ = ~new_n56701_ & ~new_n56704_;
  assign new_n57035_ = ~new_n57033_ & ~new_n57034_;
  assign new_n57036_ = ~new_n56996_ & ~new_n57035_;
  assign new_n57037_ = ~new_n56127_ & ~new_n56648_;
  assign new_n57038_ = ~new_n56995_ & new_n57037_;
  assign \remainder[5]  = new_n57036_ | new_n57038_;
  assign new_n57040_ = ~new_n56649_ & new_n56709_;
  assign new_n57041_ = ~new_n56705_ & new_n57040_;
  assign new_n57042_ = ~new_n56706_ & ~new_n56709_;
  assign new_n57043_ = ~new_n57041_ & ~new_n57042_;
  assign new_n57044_ = ~new_n56996_ & ~new_n57043_;
  assign new_n57045_ = ~new_n56127_ & ~new_n56639_;
  assign new_n57046_ = ~new_n56995_ & new_n57045_;
  assign \remainder[6]  = new_n57044_ | new_n57046_;
  assign new_n57048_ = ~new_n56640_ & new_n56714_;
  assign new_n57049_ = ~new_n56710_ & new_n57048_;
  assign new_n57050_ = ~new_n56711_ & ~new_n56714_;
  assign new_n57051_ = ~new_n57049_ & ~new_n57050_;
  assign new_n57052_ = ~new_n56996_ & ~new_n57051_;
  assign new_n57053_ = ~new_n56127_ & ~new_n56630_;
  assign new_n57054_ = ~new_n56995_ & new_n57053_;
  assign \remainder[7]  = new_n57052_ | new_n57054_;
  assign new_n57056_ = ~new_n56631_ & new_n56719_;
  assign new_n57057_ = ~new_n56715_ & new_n57056_;
  assign new_n57058_ = ~new_n56716_ & ~new_n56719_;
  assign new_n57059_ = ~new_n57057_ & ~new_n57058_;
  assign new_n57060_ = ~new_n56996_ & ~new_n57059_;
  assign new_n57061_ = ~new_n56127_ & ~new_n56621_;
  assign new_n57062_ = ~new_n56995_ & new_n57061_;
  assign \remainder[8]  = new_n57060_ | new_n57062_;
  assign new_n57064_ = ~new_n56622_ & new_n56724_;
  assign new_n57065_ = ~new_n56720_ & new_n57064_;
  assign new_n57066_ = ~new_n56721_ & ~new_n56724_;
  assign new_n57067_ = ~new_n57065_ & ~new_n57066_;
  assign new_n57068_ = ~new_n56996_ & ~new_n57067_;
  assign new_n57069_ = ~new_n56127_ & ~new_n56612_;
  assign new_n57070_ = ~new_n56995_ & new_n57069_;
  assign \remainder[9]  = new_n57068_ | new_n57070_;
  assign new_n57072_ = ~new_n56613_ & new_n56729_;
  assign new_n57073_ = ~new_n56725_ & new_n57072_;
  assign new_n57074_ = ~new_n56726_ & ~new_n56729_;
  assign new_n57075_ = ~new_n57073_ & ~new_n57074_;
  assign new_n57076_ = ~new_n56996_ & ~new_n57075_;
  assign new_n57077_ = ~new_n56127_ & ~new_n56603_;
  assign new_n57078_ = ~new_n56995_ & new_n57077_;
  assign \remainder[10]  = new_n57076_ | new_n57078_;
  assign new_n57080_ = ~new_n56604_ & new_n56734_;
  assign new_n57081_ = ~new_n56730_ & new_n57080_;
  assign new_n57082_ = ~new_n56731_ & ~new_n56734_;
  assign new_n57083_ = ~new_n57081_ & ~new_n57082_;
  assign new_n57084_ = ~new_n56996_ & ~new_n57083_;
  assign new_n57085_ = ~new_n56127_ & ~new_n56594_;
  assign new_n57086_ = ~new_n56995_ & new_n57085_;
  assign \remainder[11]  = new_n57084_ | new_n57086_;
  assign new_n57088_ = ~new_n56595_ & new_n56739_;
  assign new_n57089_ = ~new_n56735_ & new_n57088_;
  assign new_n57090_ = ~new_n56736_ & ~new_n56739_;
  assign new_n57091_ = ~new_n57089_ & ~new_n57090_;
  assign new_n57092_ = ~new_n56996_ & ~new_n57091_;
  assign new_n57093_ = ~new_n56127_ & ~new_n56585_;
  assign new_n57094_ = ~new_n56995_ & new_n57093_;
  assign \remainder[12]  = new_n57092_ | new_n57094_;
  assign new_n57096_ = ~new_n56586_ & new_n56744_;
  assign new_n57097_ = ~new_n56740_ & new_n57096_;
  assign new_n57098_ = ~new_n56741_ & ~new_n56744_;
  assign new_n57099_ = ~new_n57097_ & ~new_n57098_;
  assign new_n57100_ = ~new_n56996_ & ~new_n57099_;
  assign new_n57101_ = ~new_n56127_ & ~new_n56576_;
  assign new_n57102_ = ~new_n56995_ & new_n57101_;
  assign \remainder[13]  = new_n57100_ | new_n57102_;
  assign new_n57104_ = ~new_n56577_ & new_n56749_;
  assign new_n57105_ = ~new_n56745_ & new_n57104_;
  assign new_n57106_ = ~new_n56746_ & ~new_n56749_;
  assign new_n57107_ = ~new_n57105_ & ~new_n57106_;
  assign new_n57108_ = ~new_n56996_ & ~new_n57107_;
  assign new_n57109_ = ~new_n56127_ & ~new_n56567_;
  assign new_n57110_ = ~new_n56995_ & new_n57109_;
  assign \remainder[14]  = new_n57108_ | new_n57110_;
  assign new_n57112_ = ~new_n56568_ & new_n56754_;
  assign new_n57113_ = ~new_n56750_ & new_n57112_;
  assign new_n57114_ = ~new_n56751_ & ~new_n56754_;
  assign new_n57115_ = ~new_n57113_ & ~new_n57114_;
  assign new_n57116_ = ~new_n56996_ & ~new_n57115_;
  assign new_n57117_ = ~new_n56127_ & ~new_n56558_;
  assign new_n57118_ = ~new_n56995_ & new_n57117_;
  assign \remainder[15]  = new_n57116_ | new_n57118_;
  assign new_n57120_ = ~new_n56559_ & new_n56759_;
  assign new_n57121_ = ~new_n56755_ & new_n57120_;
  assign new_n57122_ = ~new_n56756_ & ~new_n56759_;
  assign new_n57123_ = ~new_n57121_ & ~new_n57122_;
  assign new_n57124_ = ~new_n56996_ & ~new_n57123_;
  assign new_n57125_ = ~new_n56127_ & ~new_n56549_;
  assign new_n57126_ = ~new_n56995_ & new_n57125_;
  assign \remainder[16]  = new_n57124_ | new_n57126_;
  assign new_n57128_ = ~new_n56550_ & new_n56764_;
  assign new_n57129_ = ~new_n56760_ & new_n57128_;
  assign new_n57130_ = ~new_n56761_ & ~new_n56764_;
  assign new_n57131_ = ~new_n57129_ & ~new_n57130_;
  assign new_n57132_ = ~new_n56996_ & ~new_n57131_;
  assign new_n57133_ = ~new_n56127_ & ~new_n56540_;
  assign new_n57134_ = ~new_n56995_ & new_n57133_;
  assign \remainder[17]  = new_n57132_ | new_n57134_;
  assign new_n57136_ = ~new_n56541_ & new_n56769_;
  assign new_n57137_ = ~new_n56765_ & new_n57136_;
  assign new_n57138_ = ~new_n56766_ & ~new_n56769_;
  assign new_n57139_ = ~new_n57137_ & ~new_n57138_;
  assign new_n57140_ = ~new_n56996_ & ~new_n57139_;
  assign new_n57141_ = ~new_n56127_ & ~new_n56531_;
  assign new_n57142_ = ~new_n56995_ & new_n57141_;
  assign \remainder[18]  = new_n57140_ | new_n57142_;
  assign new_n57144_ = ~new_n56532_ & new_n56774_;
  assign new_n57145_ = ~new_n56770_ & new_n57144_;
  assign new_n57146_ = ~new_n56771_ & ~new_n56774_;
  assign new_n57147_ = ~new_n57145_ & ~new_n57146_;
  assign new_n57148_ = ~new_n56996_ & ~new_n57147_;
  assign new_n57149_ = ~new_n56127_ & ~new_n56522_;
  assign new_n57150_ = ~new_n56995_ & new_n57149_;
  assign \remainder[19]  = new_n57148_ | new_n57150_;
  assign new_n57152_ = ~new_n56523_ & new_n56779_;
  assign new_n57153_ = ~new_n56775_ & new_n57152_;
  assign new_n57154_ = ~new_n56776_ & ~new_n56779_;
  assign new_n57155_ = ~new_n57153_ & ~new_n57154_;
  assign new_n57156_ = ~new_n56996_ & ~new_n57155_;
  assign new_n57157_ = ~new_n56127_ & ~new_n56513_;
  assign new_n57158_ = ~new_n56995_ & new_n57157_;
  assign \remainder[20]  = new_n57156_ | new_n57158_;
  assign new_n57160_ = ~new_n56514_ & new_n56784_;
  assign new_n57161_ = ~new_n56780_ & new_n57160_;
  assign new_n57162_ = ~new_n56781_ & ~new_n56784_;
  assign new_n57163_ = ~new_n57161_ & ~new_n57162_;
  assign new_n57164_ = ~new_n56996_ & ~new_n57163_;
  assign new_n57165_ = ~new_n56127_ & ~new_n56504_;
  assign new_n57166_ = ~new_n56995_ & new_n57165_;
  assign \remainder[21]  = new_n57164_ | new_n57166_;
  assign new_n57168_ = ~new_n56505_ & new_n56789_;
  assign new_n57169_ = ~new_n56785_ & new_n57168_;
  assign new_n57170_ = ~new_n56786_ & ~new_n56789_;
  assign new_n57171_ = ~new_n57169_ & ~new_n57170_;
  assign new_n57172_ = ~new_n56996_ & ~new_n57171_;
  assign new_n57173_ = ~new_n56127_ & ~new_n56495_;
  assign new_n57174_ = ~new_n56995_ & new_n57173_;
  assign \remainder[22]  = new_n57172_ | new_n57174_;
  assign new_n57176_ = ~new_n56496_ & new_n56794_;
  assign new_n57177_ = ~new_n56790_ & new_n57176_;
  assign new_n57178_ = ~new_n56791_ & ~new_n56794_;
  assign new_n57179_ = ~new_n57177_ & ~new_n57178_;
  assign new_n57180_ = ~new_n56996_ & ~new_n57179_;
  assign new_n57181_ = ~new_n56127_ & ~new_n56486_;
  assign new_n57182_ = ~new_n56995_ & new_n57181_;
  assign \remainder[23]  = new_n57180_ | new_n57182_;
  assign new_n57184_ = ~new_n56487_ & new_n56799_;
  assign new_n57185_ = ~new_n56795_ & new_n57184_;
  assign new_n57186_ = ~new_n56796_ & ~new_n56799_;
  assign new_n57187_ = ~new_n57185_ & ~new_n57186_;
  assign new_n57188_ = ~new_n56996_ & ~new_n57187_;
  assign new_n57189_ = ~new_n56127_ & ~new_n56477_;
  assign new_n57190_ = ~new_n56995_ & new_n57189_;
  assign \remainder[24]  = new_n57188_ | new_n57190_;
  assign new_n57192_ = ~new_n56478_ & new_n56804_;
  assign new_n57193_ = ~new_n56800_ & new_n57192_;
  assign new_n57194_ = ~new_n56801_ & ~new_n56804_;
  assign new_n57195_ = ~new_n57193_ & ~new_n57194_;
  assign new_n57196_ = ~new_n56996_ & ~new_n57195_;
  assign new_n57197_ = ~new_n56127_ & ~new_n56468_;
  assign new_n57198_ = ~new_n56995_ & new_n57197_;
  assign \remainder[25]  = new_n57196_ | new_n57198_;
  assign new_n57200_ = ~new_n56469_ & new_n56809_;
  assign new_n57201_ = ~new_n56805_ & new_n57200_;
  assign new_n57202_ = ~new_n56806_ & ~new_n56809_;
  assign new_n57203_ = ~new_n57201_ & ~new_n57202_;
  assign new_n57204_ = ~new_n56996_ & ~new_n57203_;
  assign new_n57205_ = ~new_n56127_ & ~new_n56459_;
  assign new_n57206_ = ~new_n56995_ & new_n57205_;
  assign \remainder[26]  = new_n57204_ | new_n57206_;
  assign new_n57208_ = ~new_n56460_ & new_n56814_;
  assign new_n57209_ = ~new_n56810_ & new_n57208_;
  assign new_n57210_ = ~new_n56811_ & ~new_n56814_;
  assign new_n57211_ = ~new_n57209_ & ~new_n57210_;
  assign new_n57212_ = ~new_n56996_ & ~new_n57211_;
  assign new_n57213_ = ~new_n56127_ & ~new_n56450_;
  assign new_n57214_ = ~new_n56995_ & new_n57213_;
  assign \remainder[27]  = new_n57212_ | new_n57214_;
  assign new_n57216_ = ~new_n56451_ & new_n56819_;
  assign new_n57217_ = ~new_n56815_ & new_n57216_;
  assign new_n57218_ = ~new_n56816_ & ~new_n56819_;
  assign new_n57219_ = ~new_n57217_ & ~new_n57218_;
  assign new_n57220_ = ~new_n56996_ & ~new_n57219_;
  assign new_n57221_ = ~new_n56127_ & ~new_n56441_;
  assign new_n57222_ = ~new_n56995_ & new_n57221_;
  assign \remainder[28]  = new_n57220_ | new_n57222_;
  assign new_n57224_ = ~new_n56442_ & new_n56824_;
  assign new_n57225_ = ~new_n56820_ & new_n57224_;
  assign new_n57226_ = ~new_n56821_ & ~new_n56824_;
  assign new_n57227_ = ~new_n57225_ & ~new_n57226_;
  assign new_n57228_ = ~new_n56996_ & ~new_n57227_;
  assign new_n57229_ = ~new_n56127_ & ~new_n56432_;
  assign new_n57230_ = ~new_n56995_ & new_n57229_;
  assign \remainder[29]  = new_n57228_ | new_n57230_;
  assign new_n57232_ = ~new_n56433_ & new_n56829_;
  assign new_n57233_ = ~new_n56825_ & new_n57232_;
  assign new_n57234_ = ~new_n56826_ & ~new_n56829_;
  assign new_n57235_ = ~new_n57233_ & ~new_n57234_;
  assign new_n57236_ = ~new_n56996_ & ~new_n57235_;
  assign new_n57237_ = ~new_n56127_ & ~new_n56423_;
  assign new_n57238_ = ~new_n56995_ & new_n57237_;
  assign \remainder[30]  = new_n57236_ | new_n57238_;
  assign new_n57240_ = ~new_n56424_ & new_n56834_;
  assign new_n57241_ = ~new_n56830_ & new_n57240_;
  assign new_n57242_ = ~new_n56831_ & ~new_n56834_;
  assign new_n57243_ = ~new_n57241_ & ~new_n57242_;
  assign new_n57244_ = ~new_n56996_ & ~new_n57243_;
  assign new_n57245_ = ~new_n56127_ & ~new_n56414_;
  assign new_n57246_ = ~new_n56995_ & new_n57245_;
  assign \remainder[31]  = new_n57244_ | new_n57246_;
  assign new_n57248_ = ~new_n56415_ & new_n56839_;
  assign new_n57249_ = ~new_n56835_ & new_n57248_;
  assign new_n57250_ = ~new_n56836_ & ~new_n56839_;
  assign new_n57251_ = ~new_n57249_ & ~new_n57250_;
  assign new_n57252_ = ~new_n56996_ & ~new_n57251_;
  assign new_n57253_ = ~new_n56127_ & ~new_n56405_;
  assign new_n57254_ = ~new_n56995_ & new_n57253_;
  assign \remainder[32]  = new_n57252_ | new_n57254_;
  assign new_n57256_ = ~new_n56406_ & new_n56844_;
  assign new_n57257_ = ~new_n56840_ & new_n57256_;
  assign new_n57258_ = ~new_n56841_ & ~new_n56844_;
  assign new_n57259_ = ~new_n57257_ & ~new_n57258_;
  assign new_n57260_ = ~new_n56996_ & ~new_n57259_;
  assign new_n57261_ = ~new_n56127_ & ~new_n56396_;
  assign new_n57262_ = ~new_n56995_ & new_n57261_;
  assign \remainder[33]  = new_n57260_ | new_n57262_;
  assign new_n57264_ = ~new_n56397_ & new_n56849_;
  assign new_n57265_ = ~new_n56845_ & new_n57264_;
  assign new_n57266_ = ~new_n56846_ & ~new_n56849_;
  assign new_n57267_ = ~new_n57265_ & ~new_n57266_;
  assign new_n57268_ = ~new_n56996_ & ~new_n57267_;
  assign new_n57269_ = ~new_n56127_ & ~new_n56387_;
  assign new_n57270_ = ~new_n56995_ & new_n57269_;
  assign \remainder[34]  = new_n57268_ | new_n57270_;
  assign new_n57272_ = ~new_n56388_ & new_n56854_;
  assign new_n57273_ = ~new_n56850_ & new_n57272_;
  assign new_n57274_ = ~new_n56851_ & ~new_n56854_;
  assign new_n57275_ = ~new_n57273_ & ~new_n57274_;
  assign new_n57276_ = ~new_n56996_ & ~new_n57275_;
  assign new_n57277_ = ~new_n56127_ & ~new_n56378_;
  assign new_n57278_ = ~new_n56995_ & new_n57277_;
  assign \remainder[35]  = new_n57276_ | new_n57278_;
  assign new_n57280_ = ~new_n56379_ & new_n56859_;
  assign new_n57281_ = ~new_n56855_ & new_n57280_;
  assign new_n57282_ = ~new_n56856_ & ~new_n56859_;
  assign new_n57283_ = ~new_n57281_ & ~new_n57282_;
  assign new_n57284_ = ~new_n56996_ & ~new_n57283_;
  assign new_n57285_ = ~new_n56127_ & ~new_n56369_;
  assign new_n57286_ = ~new_n56995_ & new_n57285_;
  assign \remainder[36]  = new_n57284_ | new_n57286_;
  assign new_n57288_ = ~new_n56370_ & new_n56864_;
  assign new_n57289_ = ~new_n56860_ & new_n57288_;
  assign new_n57290_ = ~new_n56861_ & ~new_n56864_;
  assign new_n57291_ = ~new_n57289_ & ~new_n57290_;
  assign new_n57292_ = ~new_n56996_ & ~new_n57291_;
  assign new_n57293_ = ~new_n56127_ & ~new_n56360_;
  assign new_n57294_ = ~new_n56995_ & new_n57293_;
  assign \remainder[37]  = new_n57292_ | new_n57294_;
  assign new_n57296_ = ~new_n56361_ & new_n56869_;
  assign new_n57297_ = ~new_n56865_ & new_n57296_;
  assign new_n57298_ = ~new_n56866_ & ~new_n56869_;
  assign new_n57299_ = ~new_n57297_ & ~new_n57298_;
  assign new_n57300_ = ~new_n56996_ & ~new_n57299_;
  assign new_n57301_ = ~new_n56127_ & ~new_n56351_;
  assign new_n57302_ = ~new_n56995_ & new_n57301_;
  assign \remainder[38]  = new_n57300_ | new_n57302_;
  assign new_n57304_ = ~new_n56352_ & new_n56874_;
  assign new_n57305_ = ~new_n56870_ & new_n57304_;
  assign new_n57306_ = ~new_n56871_ & ~new_n56874_;
  assign new_n57307_ = ~new_n57305_ & ~new_n57306_;
  assign new_n57308_ = ~new_n56996_ & ~new_n57307_;
  assign new_n57309_ = ~new_n56127_ & ~new_n56342_;
  assign new_n57310_ = ~new_n56995_ & new_n57309_;
  assign \remainder[39]  = new_n57308_ | new_n57310_;
  assign new_n57312_ = ~new_n56343_ & new_n56879_;
  assign new_n57313_ = ~new_n56875_ & new_n57312_;
  assign new_n57314_ = ~new_n56876_ & ~new_n56879_;
  assign new_n57315_ = ~new_n57313_ & ~new_n57314_;
  assign new_n57316_ = ~new_n56996_ & ~new_n57315_;
  assign new_n57317_ = ~new_n56127_ & ~new_n56333_;
  assign new_n57318_ = ~new_n56995_ & new_n57317_;
  assign \remainder[40]  = new_n57316_ | new_n57318_;
  assign new_n57320_ = ~new_n56334_ & new_n56884_;
  assign new_n57321_ = ~new_n56880_ & new_n57320_;
  assign new_n57322_ = ~new_n56881_ & ~new_n56884_;
  assign new_n57323_ = ~new_n57321_ & ~new_n57322_;
  assign new_n57324_ = ~new_n56996_ & ~new_n57323_;
  assign new_n57325_ = ~new_n56127_ & ~new_n56324_;
  assign new_n57326_ = ~new_n56995_ & new_n57325_;
  assign \remainder[41]  = new_n57324_ | new_n57326_;
  assign new_n57328_ = ~new_n56325_ & new_n56889_;
  assign new_n57329_ = ~new_n56885_ & new_n57328_;
  assign new_n57330_ = ~new_n56886_ & ~new_n56889_;
  assign new_n57331_ = ~new_n57329_ & ~new_n57330_;
  assign new_n57332_ = ~new_n56996_ & ~new_n57331_;
  assign new_n57333_ = ~new_n56127_ & ~new_n56315_;
  assign new_n57334_ = ~new_n56995_ & new_n57333_;
  assign \remainder[42]  = new_n57332_ | new_n57334_;
  assign new_n57336_ = ~new_n56316_ & new_n56894_;
  assign new_n57337_ = ~new_n56890_ & new_n57336_;
  assign new_n57338_ = ~new_n56891_ & ~new_n56894_;
  assign new_n57339_ = ~new_n57337_ & ~new_n57338_;
  assign new_n57340_ = ~new_n56996_ & ~new_n57339_;
  assign new_n57341_ = ~new_n56127_ & ~new_n56306_;
  assign new_n57342_ = ~new_n56995_ & new_n57341_;
  assign \remainder[43]  = new_n57340_ | new_n57342_;
  assign new_n57344_ = ~new_n56307_ & new_n56899_;
  assign new_n57345_ = ~new_n56895_ & new_n57344_;
  assign new_n57346_ = ~new_n56896_ & ~new_n56899_;
  assign new_n57347_ = ~new_n57345_ & ~new_n57346_;
  assign new_n57348_ = ~new_n56996_ & ~new_n57347_;
  assign new_n57349_ = ~new_n56127_ & ~new_n56297_;
  assign new_n57350_ = ~new_n56995_ & new_n57349_;
  assign \remainder[44]  = new_n57348_ | new_n57350_;
  assign new_n57352_ = ~new_n56298_ & new_n56904_;
  assign new_n57353_ = ~new_n56900_ & new_n57352_;
  assign new_n57354_ = ~new_n56901_ & ~new_n56904_;
  assign new_n57355_ = ~new_n57353_ & ~new_n57354_;
  assign new_n57356_ = ~new_n56996_ & ~new_n57355_;
  assign new_n57357_ = ~new_n56127_ & ~new_n56288_;
  assign new_n57358_ = ~new_n56995_ & new_n57357_;
  assign \remainder[45]  = new_n57356_ | new_n57358_;
  assign new_n57360_ = ~new_n56289_ & new_n56909_;
  assign new_n57361_ = ~new_n56905_ & new_n57360_;
  assign new_n57362_ = ~new_n56906_ & ~new_n56909_;
  assign new_n57363_ = ~new_n57361_ & ~new_n57362_;
  assign new_n57364_ = ~new_n56996_ & ~new_n57363_;
  assign new_n57365_ = ~new_n56127_ & ~new_n56279_;
  assign new_n57366_ = ~new_n56995_ & new_n57365_;
  assign \remainder[46]  = new_n57364_ | new_n57366_;
  assign new_n57368_ = ~new_n56280_ & new_n56914_;
  assign new_n57369_ = ~new_n56910_ & new_n57368_;
  assign new_n57370_ = ~new_n56911_ & ~new_n56914_;
  assign new_n57371_ = ~new_n57369_ & ~new_n57370_;
  assign new_n57372_ = ~new_n56996_ & ~new_n57371_;
  assign new_n57373_ = ~new_n56127_ & ~new_n56270_;
  assign new_n57374_ = ~new_n56995_ & new_n57373_;
  assign \remainder[47]  = new_n57372_ | new_n57374_;
  assign new_n57376_ = ~new_n56271_ & new_n56919_;
  assign new_n57377_ = ~new_n56915_ & new_n57376_;
  assign new_n57378_ = ~new_n56916_ & ~new_n56919_;
  assign new_n57379_ = ~new_n57377_ & ~new_n57378_;
  assign new_n57380_ = ~new_n56996_ & ~new_n57379_;
  assign new_n57381_ = ~new_n56127_ & ~new_n56261_;
  assign new_n57382_ = ~new_n56995_ & new_n57381_;
  assign \remainder[48]  = new_n57380_ | new_n57382_;
  assign new_n57384_ = ~new_n56262_ & new_n56924_;
  assign new_n57385_ = ~new_n56920_ & new_n57384_;
  assign new_n57386_ = ~new_n56921_ & ~new_n56924_;
  assign new_n57387_ = ~new_n57385_ & ~new_n57386_;
  assign new_n57388_ = ~new_n56996_ & ~new_n57387_;
  assign new_n57389_ = ~new_n56127_ & ~new_n56252_;
  assign new_n57390_ = ~new_n56995_ & new_n57389_;
  assign \remainder[49]  = new_n57388_ | new_n57390_;
  assign new_n57392_ = ~new_n56253_ & new_n56929_;
  assign new_n57393_ = ~new_n56925_ & new_n57392_;
  assign new_n57394_ = ~new_n56926_ & ~new_n56929_;
  assign new_n57395_ = ~new_n57393_ & ~new_n57394_;
  assign new_n57396_ = ~new_n56996_ & ~new_n57395_;
  assign new_n57397_ = ~new_n56127_ & ~new_n56243_;
  assign new_n57398_ = ~new_n56995_ & new_n57397_;
  assign \remainder[50]  = new_n57396_ | new_n57398_;
  assign new_n57400_ = ~new_n56244_ & new_n56934_;
  assign new_n57401_ = ~new_n56930_ & new_n57400_;
  assign new_n57402_ = ~new_n56931_ & ~new_n56934_;
  assign new_n57403_ = ~new_n57401_ & ~new_n57402_;
  assign new_n57404_ = ~new_n56996_ & ~new_n57403_;
  assign new_n57405_ = ~new_n56127_ & ~new_n56234_;
  assign new_n57406_ = ~new_n56995_ & new_n57405_;
  assign \remainder[51]  = new_n57404_ | new_n57406_;
  assign new_n57408_ = ~new_n56235_ & new_n56939_;
  assign new_n57409_ = ~new_n56935_ & new_n57408_;
  assign new_n57410_ = ~new_n56936_ & ~new_n56939_;
  assign new_n57411_ = ~new_n57409_ & ~new_n57410_;
  assign new_n57412_ = ~new_n56996_ & ~new_n57411_;
  assign new_n57413_ = ~new_n56127_ & ~new_n56225_;
  assign new_n57414_ = ~new_n56995_ & new_n57413_;
  assign \remainder[52]  = new_n57412_ | new_n57414_;
  assign new_n57416_ = ~new_n56226_ & new_n56944_;
  assign new_n57417_ = ~new_n56940_ & new_n57416_;
  assign new_n57418_ = ~new_n56941_ & ~new_n56944_;
  assign new_n57419_ = ~new_n57417_ & ~new_n57418_;
  assign new_n57420_ = ~new_n56996_ & ~new_n57419_;
  assign new_n57421_ = ~new_n56127_ & ~new_n56216_;
  assign new_n57422_ = ~new_n56995_ & new_n57421_;
  assign \remainder[53]  = new_n57420_ | new_n57422_;
  assign new_n57424_ = ~new_n56217_ & new_n56949_;
  assign new_n57425_ = ~new_n56945_ & new_n57424_;
  assign new_n57426_ = ~new_n56946_ & ~new_n56949_;
  assign new_n57427_ = ~new_n57425_ & ~new_n57426_;
  assign new_n57428_ = ~new_n56996_ & ~new_n57427_;
  assign new_n57429_ = ~new_n56127_ & ~new_n56207_;
  assign new_n57430_ = ~new_n56995_ & new_n57429_;
  assign \remainder[54]  = new_n57428_ | new_n57430_;
  assign new_n57432_ = ~new_n56208_ & new_n56954_;
  assign new_n57433_ = ~new_n56950_ & new_n57432_;
  assign new_n57434_ = ~new_n56951_ & ~new_n56954_;
  assign new_n57435_ = ~new_n57433_ & ~new_n57434_;
  assign new_n57436_ = ~new_n56996_ & ~new_n57435_;
  assign new_n57437_ = ~new_n56127_ & ~new_n56198_;
  assign new_n57438_ = ~new_n56995_ & new_n57437_;
  assign \remainder[55]  = new_n57436_ | new_n57438_;
  assign new_n57440_ = ~new_n56199_ & new_n56959_;
  assign new_n57441_ = ~new_n56955_ & new_n57440_;
  assign new_n57442_ = ~new_n56956_ & ~new_n56959_;
  assign new_n57443_ = ~new_n57441_ & ~new_n57442_;
  assign new_n57444_ = ~new_n56996_ & ~new_n57443_;
  assign new_n57445_ = ~new_n56127_ & ~new_n56189_;
  assign new_n57446_ = ~new_n56995_ & new_n57445_;
  assign \remainder[56]  = new_n57444_ | new_n57446_;
  assign new_n57448_ = ~new_n56190_ & new_n56964_;
  assign new_n57449_ = ~new_n56960_ & new_n57448_;
  assign new_n57450_ = ~new_n56961_ & ~new_n56964_;
  assign new_n57451_ = ~new_n57449_ & ~new_n57450_;
  assign new_n57452_ = ~new_n56996_ & ~new_n57451_;
  assign new_n57453_ = ~new_n56127_ & ~new_n56180_;
  assign new_n57454_ = ~new_n56995_ & new_n57453_;
  assign \remainder[57]  = new_n57452_ | new_n57454_;
  assign new_n57456_ = ~new_n56181_ & new_n56969_;
  assign new_n57457_ = ~new_n56965_ & new_n57456_;
  assign new_n57458_ = ~new_n56966_ & ~new_n56969_;
  assign new_n57459_ = ~new_n57457_ & ~new_n57458_;
  assign new_n57460_ = ~new_n56996_ & ~new_n57459_;
  assign new_n57461_ = ~new_n56127_ & ~new_n56171_;
  assign new_n57462_ = ~new_n56995_ & new_n57461_;
  assign \remainder[58]  = new_n57460_ | new_n57462_;
  assign new_n57464_ = ~new_n56172_ & new_n56974_;
  assign new_n57465_ = ~new_n56970_ & new_n57464_;
  assign new_n57466_ = ~new_n56971_ & ~new_n56974_;
  assign new_n57467_ = ~new_n57465_ & ~new_n57466_;
  assign new_n57468_ = ~new_n56996_ & ~new_n57467_;
  assign new_n57469_ = ~new_n56127_ & ~new_n56162_;
  assign new_n57470_ = ~new_n56995_ & new_n57469_;
  assign \remainder[59]  = new_n57468_ | new_n57470_;
  assign new_n57472_ = ~new_n56163_ & new_n56979_;
  assign new_n57473_ = ~new_n56975_ & new_n57472_;
  assign new_n57474_ = ~new_n56976_ & ~new_n56979_;
  assign new_n57475_ = ~new_n57473_ & ~new_n57474_;
  assign new_n57476_ = ~new_n56996_ & ~new_n57475_;
  assign new_n57477_ = ~new_n56127_ & ~new_n56153_;
  assign new_n57478_ = ~new_n56995_ & new_n57477_;
  assign \remainder[60]  = new_n57476_ | new_n57478_;
  assign new_n57480_ = ~new_n56154_ & new_n56984_;
  assign new_n57481_ = ~new_n56980_ & new_n57480_;
  assign new_n57482_ = ~new_n56981_ & ~new_n56984_;
  assign new_n57483_ = ~new_n57481_ & ~new_n57482_;
  assign new_n57484_ = ~new_n56996_ & ~new_n57483_;
  assign new_n57485_ = ~new_n56127_ & ~new_n56144_;
  assign new_n57486_ = ~new_n56995_ & new_n57485_;
  assign \remainder[61]  = new_n57484_ | new_n57486_;
  assign new_n57488_ = ~new_n56145_ & new_n56989_;
  assign new_n57489_ = ~new_n56985_ & new_n57488_;
  assign new_n57490_ = ~new_n56986_ & ~new_n56989_;
  assign new_n57491_ = ~new_n57489_ & ~new_n57490_;
  assign new_n57492_ = ~new_n56996_ & ~new_n57491_;
  assign new_n57493_ = ~new_n56127_ & ~new_n56135_;
  assign new_n57494_ = ~new_n56995_ & new_n57493_;
  assign \remainder[62]  = new_n57492_ | new_n57494_;
  assign new_n57496_ = ~new_n56136_ & new_n56994_;
  assign new_n57497_ = ~new_n56990_ & new_n57496_;
  assign new_n57498_ = ~new_n56991_ & ~new_n56994_;
  assign new_n57499_ = ~new_n57497_ & ~new_n57498_;
  assign new_n57500_ = ~new_n56996_ & ~new_n57499_;
  assign new_n57501_ = ~new_n56126_ & ~new_n56127_;
  assign new_n57502_ = ~new_n56995_ & new_n57501_;
  assign \remainder[63]  = new_n57500_ | new_n57502_;
endmodule


