// Benchmark "testing" written by ABC on Thu Oct  8 22:16:59 2020

module testing ( 
    A302, A301, A300, A299, A298, A269, A268, A267, A266, A265, A236, A235,
    A234, A233, A232, A203, A202, A201, A200, A199, A166, A167, A168, A169,
    A170,
    A142, A141, A140, A139, A138, A109, A108, A107, A106, A105, A76, A75,
    A74, A73, A72, A43, A42, A41, A40, A39, A6, A7, A8, A9, A10  );
  input  A302, A301, A300, A299, A298, A269, A268, A267, A266, A265,
    A236, A235, A234, A233, A232, A203, A202, A201, A200, A199, A166, A167,
    A168, A169, A170;
  output A142, A141, A140, A139, A138, A109, A108, A107, A106, A105, A76, A75,
    A74, A73, A72, A43, A42, A41, A40, A39, A6, A7, A8, A9, A10;
  wire new_A198_, new_A197_, new_A196_, new_A195_, new_A194_, new_A193_,
    new_A192_, new_A191_, new_A190_, new_A189_, new_A188_, new_A187_,
    new_A186_, new_A185_, new_A184_, new_A183_, new_A182_, new_A181_,
    new_A180_, new_A179_, new_A178_, new_A177_, new_A176_, new_A175_,
    new_A174_, new_A173_, new_A172_, new_A171_, new_A204_, new_A205_,
    new_A206_, new_A207_, new_A208_, new_A209_, new_A210_, new_A211_,
    new_A212_, new_A213_, new_A214_, new_A215_, new_A216_, new_A217_,
    new_A218_, new_A219_, new_A220_, new_A221_, new_A222_, new_A223_,
    new_A224_, new_A225_, new_A226_, new_A227_, new_A228_, new_A229_,
    new_A230_, new_A231_, new_A237_, new_A238_, new_A239_, new_A240_,
    new_A241_, new_A242_, new_A243_, new_A244_, new_A245_, new_A246_,
    new_A247_, new_A248_, new_A249_, new_A250_, new_A251_, new_A252_,
    new_A253_, new_A254_, new_A255_, new_A256_, new_A257_, new_A258_,
    new_A259_, new_A260_, new_A261_, new_A262_, new_A263_, new_A264_,
    new_A270_, new_A271_, new_A272_, new_A273_, new_A274_, new_A275_,
    new_A276_, new_A277_, new_A278_, new_A279_, new_A280_, new_A281_,
    new_A282_, new_A283_, new_A284_, new_A285_, new_A286_, new_A287_,
    new_A288_, new_A289_, new_A290_, new_A291_, new_A292_, new_A293_,
    new_A294_, new_A295_, new_A296_, new_A297_, new_A303_, new_A304_,
    new_A305_, new_A306_, new_A307_, new_A308_, new_A309_, new_A310_,
    new_A311_, new_A312_, new_A313_, new_A314_, new_A315_, new_A316_,
    new_A317_, new_A318_, new_A319_, new_A320_, new_A321_, new_A322_,
    new_A323_, new_A324_, new_A325_, new_A326_, new_A327_, new_A328_,
    new_A329_, new_A330_, new_A165_, new_A164_, new_A163_, new_A162_,
    new_A161_, new_A160_, new_A159_, new_A158_, new_A157_, new_A156_,
    new_A155_, new_A154_, new_A153_, new_A152_, new_A151_, new_A150_,
    new_A149_, new_A148_, new_A147_, new_A146_, new_A145_, new_A144_,
    new_A143_, new_A137_, new_A136_, new_A135_, new_A134_, new_A133_,
    new_A132_, new_A131_, new_A130_, new_A129_, new_A128_, new_A127_,
    new_A126_, new_A125_, new_A124_, new_A123_, new_A122_, new_A121_,
    new_A120_, new_A119_, new_A118_, new_A117_, new_A116_, new_A115_,
    new_A114_, new_A113_, new_A112_, new_A111_, new_A110_, new_A104_,
    new_A103_, new_A102_, new_A101_, new_A100_, new_A99_, new_A98_,
    new_A97_, new_A96_, new_A95_, new_A94_, new_A93_, new_A92_, new_A91_,
    new_A90_, new_A89_, new_A88_, new_A87_, new_A86_, new_A85_, new_A84_,
    new_A83_, new_A82_, new_A81_, new_A80_, new_A79_, new_A78_, new_A77_,
    new_A71_, new_A70_, new_A69_, new_A68_, new_A67_, new_A66_, new_A65_,
    new_A64_, new_A63_, new_A62_, new_A61_, new_A60_, new_A59_, new_A58_,
    new_A57_, new_A56_, new_A55_, new_A54_, new_A53_, new_A52_, new_A51_,
    new_A50_, new_A49_, new_A48_, new_A47_, new_A46_, new_A45_, new_A44_,
    new_A38_, new_A37_, new_A36_, new_A35_, new_A34_, new_A1_, new_A2_,
    new_A3_, new_A4_, new_A5_, new_A11_, new_A12_, new_A13_, new_A14_,
    new_A15_, new_A16_, new_A17_, new_A18_, new_A19_, new_A20_, new_A21_,
    new_A22_, new_A23_, new_A24_, new_A25_, new_A26_, new_A27_, new_A28_,
    new_A29_, new_A30_, new_A31_, new_A32_, new_A33_;
  assign new_A198_ = new_A176_ & new_A191_;
  assign new_A197_ = ~new_A176_ & ~new_A198_;
  assign new_A196_ = new_A176_ | new_A191_;
  assign new_A195_ = ~A169 | ~A170;
  assign new_A194_ = new_A176_ | new_A191_;
  assign new_A193_ = ~new_A192_ & ~new_A176_;
  assign new_A192_ = new_A176_ & new_A191_;
  assign new_A191_ = ~A167 | ~A168;
  assign new_A190_ = A168 & new_A180_;
  assign new_A189_ = A169 | new_A176_;
  assign new_A188_ = A169 | A170;
  assign new_A187_ = ~new_A197_ | ~new_A196_;
  assign new_A186_ = new_A195_ & new_A188_;
  assign new_A185_ = A169 ^ new_A176_;
  assign new_A184_ = ~new_A193_ | ~new_A194_;
  assign new_A183_ = ~A168 ^ new_A180_;
  assign new_A182_ = new_A190_ | A167;
  assign new_A181_ = new_A187_ & A168;
  assign new_A180_ = new_A189_ & new_A188_;
  assign new_A179_ = new_A184_ & A168;
  assign new_A178_ = new_A186_ & new_A185_;
  assign new_A177_ = new_A178_ ^ A168;
  assign new_A176_ = A166 ^ A167;
  assign new_A175_ = new_A176_ & new_A183_;
  assign new_A174_ = new_A176_ & new_A182_;
  assign new_A173_ = new_A181_ | new_A180_;
  assign new_A172_ = new_A179_ | new_A178_;
  assign new_A171_ = new_A177_ & new_A176_;
  assign new_A204_ = new_A210_ & new_A209_;
  assign new_A205_ = new_A212_ | new_A211_;
  assign new_A206_ = new_A214_ | new_A213_;
  assign new_A207_ = new_A209_ & new_A215_;
  assign new_A208_ = new_A209_ & new_A216_;
  assign new_A209_ = A199 ^ A200;
  assign new_A210_ = new_A211_ ^ A201;
  assign new_A211_ = new_A219_ & new_A218_;
  assign new_A212_ = new_A217_ & A201;
  assign new_A213_ = new_A222_ & new_A221_;
  assign new_A214_ = new_A220_ & A201;
  assign new_A215_ = new_A223_ | A200;
  assign new_A216_ = ~A201 ^ new_A213_;
  assign new_A217_ = ~new_A226_ | ~new_A227_;
  assign new_A218_ = A202 ^ new_A209_;
  assign new_A219_ = new_A228_ & new_A221_;
  assign new_A220_ = ~new_A230_ | ~new_A229_;
  assign new_A221_ = A202 | A203;
  assign new_A222_ = A202 | new_A209_;
  assign new_A223_ = A201 & new_A213_;
  assign new_A224_ = ~A200 | ~A201;
  assign new_A225_ = new_A209_ & new_A224_;
  assign new_A226_ = ~new_A225_ & ~new_A209_;
  assign new_A227_ = new_A209_ | new_A224_;
  assign new_A228_ = ~A202 | ~A203;
  assign new_A229_ = new_A209_ | new_A224_;
  assign new_A230_ = ~new_A209_ & ~new_A231_;
  assign new_A231_ = new_A209_ & new_A224_;
  assign new_A237_ = new_A243_ & new_A242_;
  assign new_A238_ = new_A245_ | new_A244_;
  assign new_A239_ = new_A247_ | new_A246_;
  assign new_A240_ = new_A242_ & new_A248_;
  assign new_A241_ = new_A242_ & new_A249_;
  assign new_A242_ = A232 ^ A233;
  assign new_A243_ = new_A244_ ^ A234;
  assign new_A244_ = new_A252_ & new_A251_;
  assign new_A245_ = new_A250_ & A234;
  assign new_A246_ = new_A255_ & new_A254_;
  assign new_A247_ = new_A253_ & A234;
  assign new_A248_ = new_A256_ | A233;
  assign new_A249_ = ~A234 ^ new_A246_;
  assign new_A250_ = ~new_A259_ | ~new_A260_;
  assign new_A251_ = A235 ^ new_A242_;
  assign new_A252_ = new_A261_ & new_A254_;
  assign new_A253_ = ~new_A263_ | ~new_A262_;
  assign new_A254_ = A235 | A236;
  assign new_A255_ = A235 | new_A242_;
  assign new_A256_ = A234 & new_A246_;
  assign new_A257_ = ~A233 | ~A234;
  assign new_A258_ = new_A242_ & new_A257_;
  assign new_A259_ = ~new_A258_ & ~new_A242_;
  assign new_A260_ = new_A242_ | new_A257_;
  assign new_A261_ = ~A235 | ~A236;
  assign new_A262_ = new_A242_ | new_A257_;
  assign new_A263_ = ~new_A242_ & ~new_A264_;
  assign new_A264_ = new_A242_ & new_A257_;
  assign new_A270_ = new_A276_ & new_A275_;
  assign new_A271_ = new_A278_ | new_A277_;
  assign new_A272_ = new_A280_ | new_A279_;
  assign new_A273_ = new_A275_ & new_A281_;
  assign new_A274_ = new_A275_ & new_A282_;
  assign new_A275_ = A265 ^ A266;
  assign new_A276_ = new_A277_ ^ A267;
  assign new_A277_ = new_A285_ & new_A284_;
  assign new_A278_ = new_A283_ & A267;
  assign new_A279_ = new_A288_ & new_A287_;
  assign new_A280_ = new_A286_ & A267;
  assign new_A281_ = new_A289_ | A266;
  assign new_A282_ = ~A267 ^ new_A279_;
  assign new_A283_ = ~new_A292_ | ~new_A293_;
  assign new_A284_ = A268 ^ new_A275_;
  assign new_A285_ = new_A294_ & new_A287_;
  assign new_A286_ = ~new_A296_ | ~new_A295_;
  assign new_A287_ = A268 | A269;
  assign new_A288_ = A268 | new_A275_;
  assign new_A289_ = A267 & new_A279_;
  assign new_A290_ = ~A266 | ~A267;
  assign new_A291_ = new_A275_ & new_A290_;
  assign new_A292_ = ~new_A291_ & ~new_A275_;
  assign new_A293_ = new_A275_ | new_A290_;
  assign new_A294_ = ~A268 | ~A269;
  assign new_A295_ = new_A275_ | new_A290_;
  assign new_A296_ = ~new_A275_ & ~new_A297_;
  assign new_A297_ = new_A275_ & new_A290_;
  assign new_A303_ = new_A309_ & new_A308_;
  assign new_A304_ = new_A311_ | new_A310_;
  assign new_A305_ = new_A313_ | new_A312_;
  assign new_A306_ = new_A308_ & new_A314_;
  assign new_A307_ = new_A308_ & new_A315_;
  assign new_A308_ = A298 ^ A299;
  assign new_A309_ = new_A310_ ^ A300;
  assign new_A310_ = new_A318_ & new_A317_;
  assign new_A311_ = new_A316_ & A300;
  assign new_A312_ = new_A321_ & new_A320_;
  assign new_A313_ = new_A319_ & A300;
  assign new_A314_ = new_A322_ | A299;
  assign new_A315_ = ~A300 ^ new_A312_;
  assign new_A316_ = ~new_A325_ | ~new_A326_;
  assign new_A317_ = A301 ^ new_A308_;
  assign new_A318_ = new_A327_ & new_A320_;
  assign new_A319_ = ~new_A329_ | ~new_A328_;
  assign new_A320_ = A301 | A302;
  assign new_A321_ = A301 | new_A308_;
  assign new_A322_ = A300 & new_A312_;
  assign new_A323_ = ~A299 | ~A300;
  assign new_A324_ = new_A308_ & new_A323_;
  assign new_A325_ = ~new_A324_ & ~new_A308_;
  assign new_A326_ = new_A308_ | new_A323_;
  assign new_A327_ = ~A301 | ~A302;
  assign new_A328_ = new_A308_ | new_A323_;
  assign new_A329_ = ~new_A308_ & ~new_A330_;
  assign new_A330_ = new_A308_ & new_A323_;
  assign new_A165_ = new_A143_ & new_A158_;
  assign new_A164_ = ~new_A143_ & ~new_A165_;
  assign new_A163_ = new_A143_ | new_A158_;
  assign new_A162_ = ~new_A136_ | ~new_A137_;
  assign new_A161_ = new_A143_ | new_A158_;
  assign new_A160_ = ~new_A159_ & ~new_A143_;
  assign new_A159_ = new_A143_ & new_A158_;
  assign new_A158_ = ~new_A134_ | ~new_A135_;
  assign new_A157_ = new_A135_ & new_A147_;
  assign new_A156_ = new_A136_ | new_A143_;
  assign new_A155_ = new_A136_ | new_A137_;
  assign new_A154_ = ~new_A164_ | ~new_A163_;
  assign new_A153_ = new_A162_ & new_A155_;
  assign new_A152_ = new_A136_ ^ new_A143_;
  assign new_A151_ = ~new_A160_ | ~new_A161_;
  assign new_A150_ = ~new_A135_ ^ new_A147_;
  assign new_A149_ = new_A157_ | new_A134_;
  assign new_A148_ = new_A154_ & new_A135_;
  assign new_A147_ = new_A156_ & new_A155_;
  assign new_A146_ = new_A151_ & new_A135_;
  assign new_A145_ = new_A153_ & new_A152_;
  assign new_A144_ = new_A145_ ^ new_A135_;
  assign new_A143_ = new_A133_ ^ new_A134_;
  assign A142 = new_A143_ & new_A150_;
  assign A141 = new_A143_ & new_A149_;
  assign A140 = new_A148_ | new_A147_;
  assign A139 = new_A146_ | new_A145_;
  assign A138 = new_A144_ & new_A143_;
  assign new_A137_ = new_A307_;
  assign new_A136_ = new_A274_;
  assign new_A135_ = new_A241_;
  assign new_A134_ = new_A208_;
  assign new_A133_ = new_A171_;
  assign new_A132_ = new_A110_ & new_A125_;
  assign new_A131_ = ~new_A110_ & ~new_A132_;
  assign new_A130_ = new_A110_ | new_A125_;
  assign new_A129_ = ~new_A103_ | ~new_A104_;
  assign new_A128_ = new_A110_ | new_A125_;
  assign new_A127_ = ~new_A126_ & ~new_A110_;
  assign new_A126_ = new_A110_ & new_A125_;
  assign new_A125_ = ~new_A101_ | ~new_A102_;
  assign new_A124_ = new_A102_ & new_A114_;
  assign new_A123_ = new_A103_ | new_A110_;
  assign new_A122_ = new_A103_ | new_A104_;
  assign new_A121_ = ~new_A131_ | ~new_A130_;
  assign new_A120_ = new_A129_ & new_A122_;
  assign new_A119_ = new_A103_ ^ new_A110_;
  assign new_A118_ = ~new_A127_ | ~new_A128_;
  assign new_A117_ = ~new_A102_ ^ new_A114_;
  assign new_A116_ = new_A124_ | new_A101_;
  assign new_A115_ = new_A121_ & new_A102_;
  assign new_A114_ = new_A123_ & new_A122_;
  assign new_A113_ = new_A118_ & new_A102_;
  assign new_A112_ = new_A120_ & new_A119_;
  assign new_A111_ = new_A112_ ^ new_A102_;
  assign new_A110_ = new_A100_ ^ new_A101_;
  assign A109 = new_A110_ & new_A117_;
  assign A108 = new_A110_ & new_A116_;
  assign A107 = new_A115_ | new_A114_;
  assign A106 = new_A113_ | new_A112_;
  assign A105 = new_A111_ & new_A110_;
  assign new_A104_ = new_A306_;
  assign new_A103_ = new_A273_;
  assign new_A102_ = new_A240_;
  assign new_A101_ = new_A207_;
  assign new_A100_ = new_A172_;
  assign new_A99_ = new_A77_ & new_A92_;
  assign new_A98_ = ~new_A77_ & ~new_A99_;
  assign new_A97_ = new_A77_ | new_A92_;
  assign new_A96_ = ~new_A70_ | ~new_A71_;
  assign new_A95_ = new_A77_ | new_A92_;
  assign new_A94_ = ~new_A93_ & ~new_A77_;
  assign new_A93_ = new_A77_ & new_A92_;
  assign new_A92_ = ~new_A68_ | ~new_A69_;
  assign new_A91_ = new_A69_ & new_A81_;
  assign new_A90_ = new_A70_ | new_A77_;
  assign new_A89_ = new_A70_ | new_A71_;
  assign new_A88_ = ~new_A98_ | ~new_A97_;
  assign new_A87_ = new_A96_ & new_A89_;
  assign new_A86_ = new_A70_ ^ new_A77_;
  assign new_A85_ = ~new_A94_ | ~new_A95_;
  assign new_A84_ = ~new_A69_ ^ new_A81_;
  assign new_A83_ = new_A91_ | new_A68_;
  assign new_A82_ = new_A88_ & new_A69_;
  assign new_A81_ = new_A90_ & new_A89_;
  assign new_A80_ = new_A85_ & new_A69_;
  assign new_A79_ = new_A87_ & new_A86_;
  assign new_A78_ = new_A79_ ^ new_A69_;
  assign new_A77_ = new_A67_ ^ new_A68_;
  assign A76 = new_A77_ & new_A84_;
  assign A75 = new_A77_ & new_A83_;
  assign A74 = new_A82_ | new_A81_;
  assign A73 = new_A80_ | new_A79_;
  assign A72 = new_A78_ & new_A77_;
  assign new_A71_ = new_A305_;
  assign new_A70_ = new_A272_;
  assign new_A69_ = new_A239_;
  assign new_A68_ = new_A206_;
  assign new_A67_ = new_A173_;
  assign new_A66_ = new_A44_ & new_A59_;
  assign new_A65_ = ~new_A44_ & ~new_A66_;
  assign new_A64_ = new_A44_ | new_A59_;
  assign new_A63_ = ~new_A37_ | ~new_A38_;
  assign new_A62_ = new_A44_ | new_A59_;
  assign new_A61_ = ~new_A60_ & ~new_A44_;
  assign new_A60_ = new_A44_ & new_A59_;
  assign new_A59_ = ~new_A35_ | ~new_A36_;
  assign new_A58_ = new_A36_ & new_A48_;
  assign new_A57_ = new_A37_ | new_A44_;
  assign new_A56_ = new_A37_ | new_A38_;
  assign new_A55_ = ~new_A65_ | ~new_A64_;
  assign new_A54_ = new_A63_ & new_A56_;
  assign new_A53_ = new_A37_ ^ new_A44_;
  assign new_A52_ = ~new_A61_ | ~new_A62_;
  assign new_A51_ = ~new_A36_ ^ new_A48_;
  assign new_A50_ = new_A58_ | new_A35_;
  assign new_A49_ = new_A55_ & new_A36_;
  assign new_A48_ = new_A57_ & new_A56_;
  assign new_A47_ = new_A52_ & new_A36_;
  assign new_A46_ = new_A54_ & new_A53_;
  assign new_A45_ = new_A46_ ^ new_A36_;
  assign new_A44_ = new_A34_ ^ new_A35_;
  assign A43 = new_A44_ & new_A51_;
  assign A42 = new_A44_ & new_A50_;
  assign A41 = new_A49_ | new_A48_;
  assign A40 = new_A47_ | new_A46_;
  assign A39 = new_A45_ & new_A44_;
  assign new_A38_ = new_A304_;
  assign new_A37_ = new_A271_;
  assign new_A36_ = new_A238_;
  assign new_A35_ = new_A205_;
  assign new_A34_ = new_A174_;
  assign new_A1_ = new_A303_;
  assign new_A2_ = new_A270_;
  assign new_A3_ = new_A237_;
  assign new_A4_ = new_A204_;
  assign new_A5_ = new_A175_;
  assign A6 = new_A12_ & new_A11_;
  assign A7 = new_A14_ | new_A13_;
  assign A8 = new_A16_ | new_A15_;
  assign A9 = new_A11_ & new_A17_;
  assign A10 = new_A11_ & new_A18_;
  assign new_A11_ = new_A1_ ^ new_A2_;
  assign new_A12_ = new_A13_ ^ new_A3_;
  assign new_A13_ = new_A21_ & new_A20_;
  assign new_A14_ = new_A19_ & new_A3_;
  assign new_A15_ = new_A24_ & new_A23_;
  assign new_A16_ = new_A22_ & new_A3_;
  assign new_A17_ = new_A25_ | new_A2_;
  assign new_A18_ = ~new_A3_ ^ new_A15_;
  assign new_A19_ = ~new_A28_ | ~new_A29_;
  assign new_A20_ = new_A4_ ^ new_A11_;
  assign new_A21_ = new_A30_ & new_A23_;
  assign new_A22_ = ~new_A32_ | ~new_A31_;
  assign new_A23_ = new_A4_ | new_A5_;
  assign new_A24_ = new_A4_ | new_A11_;
  assign new_A25_ = new_A3_ & new_A15_;
  assign new_A26_ = ~new_A2_ | ~new_A3_;
  assign new_A27_ = new_A11_ & new_A26_;
  assign new_A28_ = ~new_A27_ & ~new_A11_;
  assign new_A29_ = new_A11_ | new_A26_;
  assign new_A30_ = ~new_A4_ | ~new_A5_;
  assign new_A31_ = new_A11_ | new_A26_;
  assign new_A32_ = ~new_A11_ & ~new_A33_;
  assign new_A33_ = new_A11_ & new_A26_;
endmodule


