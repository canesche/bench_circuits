module top ( clock, 
    pg310, pg102, pg560, pg39, pg314, pg89, pg306, pg107, pg301, pg702,
    pg639, pclk, pg94, pg40, pg559, pg98, pg23, pg45, pg46, pg32, pg47,
    pg319, pg557, pg22, pg558, pg567, pg38, pg41, pg562, pg37, pg42, pg561,
    pg705, pg36, pg564, pg44, pg563,
    pg6282, pg6360, pg6370, pg4809, pg6362, pg6372, pg6364, pg5692, pg6284,
    pg6374, pg4098, pg4108, pg4109, pg4307, pg5137, pg2584, pg1293, pg3222,
    pg4104, pg4105, pg5469, pg4106, pg6728, pg4107, pg4422, pg3600, pg4100,
    pg1290, pg4099, pg4101, pg4110, pg4321, pg4102, pg5468, pg4103, pg4112,
    pg4121, pg6366, pg6368  );
  input  clock;
  input  pg310, pg102, pg560, pg39, pg314, pg89, pg306, pg107, pg301,
    pg702, pg639, pclk, pg94, pg40, pg559, pg98, pg23, pg45, pg46, pg32,
    pg47, pg319, pg557, pg22, pg558, pg567, pg38, pg41, pg562, pg37, pg42,
    pg561, pg705, pg36, pg564, pg44, pg563;
  output pg6282, pg6360, pg6370, pg4809, pg6362, pg6372, pg6364, pg5692,
    pg6284, pg6374, pg4098, pg4108, pg4109, pg4307, pg5137, pg2584, pg1293,
    pg3222, pg4104, pg4105, pg5469, pg4106, pg6728, pg4107, pg4422, pg3600,
    pg4100, pg1290, pg4099, pg4101, pg4110, pg4321, pg4102, pg5468, pg4103,
    pg4112, pg4121, pg6366, pg6368;
  reg ng230, ng197, ng434, ng25, ng205, ng266, ng204, ng524, ng699, ng658,
    ng666, ng414, ng1, ng598, ng578, ng406, ng582, ng691, ng668, ng548,
    ng485, ng694, ng422, ng500, ng19, ng532, ng210, ng236, ng677, ng512,
    ng465, ng676, ng622, ng278, ng461, ng650, ng7, ng18, ng508, ng260,
    ng689, ng692, ng24, ng277, ng453, ng445, ng2, ng279, ng594, ng269,
    ng293, ng628, ng667, ng286, ng574, ng687, ng254, ng672, ng489, ng207,
    ng441, ng6, ng290, ng680, ng616, ng554, ng625, ng426, ng402, ng218,
    ng496, ng208, ng634, ng418, ng242, ng48, ng276, ng449, ng471, ng590,
    ng437, ng528, ng486, ng551, ng685, ng281, ng430, ng698, ng545, ng682,
    ng3, ng15, ng410, ng654, ng683, ng11, ng282, ng669, ng212, ng10, ng663,
    ng606, ng43, ng520, ng297, ng14, ng280, ng646, ng206, ng211, ng541,
    ng283, ng642, ng610, ng619, ng697, ng586, ng504, ng613, ng602, ng209,
    ng631, ng662, ng571, ng536, ng28, ng638, ng675, ng457, ng33, ng29,
    ng516, ng688, ng492, ng478;
  wire new_n483_, new_n484_1_, new_n485_, new_n486_, new_n487_, new_n488_,
    new_n489_1_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_1_,
    new_n495_, new_n496_, new_n497_, new_n498_, new_n499_1_, new_n500_,
    new_n501_, new_n502_, new_n503_, new_n504_1_, new_n505_, new_n506_,
    new_n507_, new_n508_, new_n509_1_, new_n510_, new_n511_, new_n512_,
    new_n513_, new_n514_1_, new_n515_, new_n516_, new_n517_, new_n519_1_,
    new_n520_, new_n522_, new_n524_1_, new_n525_, new_n527_, new_n529_1_,
    new_n531_, new_n533_, new_n534_1_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_1_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_1_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_1_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_1_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_1_, new_n560_, new_n561_,
    new_n563_, new_n566_, new_n568_, new_n570_, new_n572_, new_n573_,
    new_n574_1_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_1_,
    new_n580_, new_n581_, new_n582_, new_n584_1_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_1_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_1_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_1_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_1_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_1_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_1_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_1_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_1_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_1_, new_n630_, new_n631_, new_n633_, new_n634_1_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_1_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_1_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_1_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_1_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_1_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_1_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_1_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_1_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_1_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_1_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_1_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_1_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_1_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_1_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_1_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_1_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_1_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_1_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_1_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_1_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_1_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_1_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_1_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_1_, new_n756_,
    new_n757_, new_n758_, new_n759_1_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_1_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_1_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_1_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_1_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_1_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_1_, new_n790_, new_n792_, new_n793_,
    new_n794_1_, new_n795_, new_n796_, new_n797_, new_n799_1_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_1_, new_n805_, new_n808_,
    new_n809_1_, new_n810_, new_n811_, new_n813_, new_n814_1_, new_n815_,
    new_n816_, new_n817_, new_n820_, new_n821_, new_n823_, new_n824_1_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n850_, new_n851_,
    new_n853_, new_n854_, new_n855_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n921_, new_n922_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n988_,
    new_n989_, new_n991_, new_n992_, new_n994_, new_n995_, new_n996_,
    new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_,
    new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_,
    new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_,
    new_n1015_, new_n1016_, new_n1017_, new_n1019_, new_n1020_, new_n1021_,
    new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_,
    new_n1028_, new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_,
    new_n1035_, new_n1037_, new_n1038_, new_n1039_, new_n1041_, new_n1042_,
    new_n1044_, new_n1045_, new_n1047_, new_n1048_, new_n1050_, new_n1051_,
    new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_,
    new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_,
    new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_,
    new_n1070_, new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_,
    new_n1076_, new_n1078_, new_n1079_, new_n1080_, new_n1082_, new_n1083_,
    new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1090_,
    new_n1091_, new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_,
    new_n1098_, new_n1099_, new_n1100_, new_n1102_, new_n1103_, new_n1104_,
    new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_,
    new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_,
    new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_,
    new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_,
    new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_,
    new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_,
    new_n1141_, new_n1142_, new_n1143_, new_n1145_, new_n1146_, new_n1147_,
    new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1154_,
    new_n1155_, new_n1157_, new_n1158_, new_n1160_, new_n1161_, new_n1163_,
    new_n1164_, new_n1166_, new_n1167_, new_n1169_, new_n1170_, new_n1172_,
    new_n1173_, new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_,
    new_n1180_, new_n1181_, new_n1182_, new_n1184_, new_n1185_, new_n1187_,
    new_n1188_, new_n1190_, new_n1191_, new_n1192_, new_n1194_, new_n1195_,
    new_n1196_, new_n1197_, new_n1199_, new_n1200_, new_n1202_, new_n1203_,
    new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1210_,
    new_n1211_, new_n1213_, new_n1214_, new_n1216_, new_n1217_, new_n1218_,
    new_n1220_, new_n1221_, new_n1223_, new_n1224_, new_n1225_, new_n1227_,
    new_n1228_, new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_,
    new_n1236_, new_n1238_, new_n1239_, new_n1240_, new_n1242_, new_n1243_,
    new_n1245_, new_n1246_, new_n1248_, new_n1249_, new_n1250_, new_n1251_,
    new_n1253_, new_n1254_, new_n1256_, new_n1257_, new_n1258_, new_n1259_,
    new_n1261_, new_n1262_, new_n1264_, new_n1265_, new_n1267_, new_n1268_,
    new_n1270_, new_n1271_, new_n1273_, new_n1274_, new_n1276_, new_n1277_,
    new_n1278_, new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_,
    new_n1284_, new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_,
    new_n1290_, new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_,
    new_n1296_, new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_,
    new_n1302_, new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1308_,
    new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_,
    new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1320_,
    new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_,
    new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_,
    new_n1333_, new_n1334_, new_n1335_, new_n1337_, new_n1338_, new_n1340_,
    new_n1341_, new_n1342_, new_n1343_, new_n1345_, new_n1346_, new_n1347_,
    new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_, new_n1353_,
    new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1358_, new_n1359_,
    new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_,
    new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_, new_n1371_,
    new_n1373_, new_n1374_, new_n1375_, new_n1376_, new_n1377_, new_n1378_,
    new_n1379_, new_n1380_, new_n1382_, new_n1383_, new_n1385_, new_n1387_,
    new_n1388_, new_n1390_, new_n1391_, new_n1392_, new_n1394_, new_n1395_,
    new_n1396_, new_n1397_, new_n1398_, new_n1399_, new_n1400_, new_n1401_,
    new_n1402_, new_n1403_, new_n1404_, new_n1405_, new_n1406_, new_n1407_,
    new_n1408_, new_n1409_, new_n1410_, new_n1411_, new_n1412_, new_n1413_,
    new_n1414_, new_n1415_, new_n1416_, new_n1417_, new_n1418_, new_n1419_,
    new_n1420_, new_n1421_, new_n1422_, new_n1423_, new_n1424_, new_n1425_,
    new_n1426_, new_n1427_, new_n1428_, new_n1430_, new_n1431_, new_n1433_,
    new_n1434_, new_n1436_, new_n1437_, new_n1439_, new_n1440_, new_n1441_,
    new_n1443_, new_n1444_, new_n1446_, new_n1447_, new_n1448_, new_n1449_,
    new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1455_, new_n1456_,
    new_n1458_, new_n1459_, new_n1460_, new_n1462_, new_n1463_, new_n1464_,
    new_n1466_, new_n1467_, new_n1468_, new_n1470_, new_n1471_, new_n1472_,
    new_n1474_, new_n1475_, new_n1477_, new_n1478_, new_n1479_, new_n1480_,
    new_n1483_, new_n1484_, new_n1485_, new_n1487_, new_n1488_, new_n1489_,
    new_n1490_, new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1496_,
    new_n1497_, new_n1498_, new_n1500_, new_n1501_, new_n1503_, new_n1504_,
    new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_,
    new_n1512_, new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_,
    new_n1518_, new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_,
    new_n1524_, new_n1525_, new_n1526_, new_n1527_, new_n1529_, new_n1530_,
    new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_, new_n1536_,
    new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1542_,
    new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_, new_n1548_,
    new_n1549_, new_n1550_, new_n1552_, new_n1553_, new_n1555_, n154, n159,
    n164, n169, n174, n179, n184, n189, n194, n199, n204, n209, n214, n219,
    n224, n229, n234, n239, n244, n249, n254, n259, n264, n269, n274, n279,
    n284, n289, n294, n299, n304, n309, n314, n319, n324, n329, n334, n339,
    n344, n349, n354, n359, n364, n369, n374, n379, n384, n389, n394, n399,
    n404, n409, n414, n419, n424, n429, n434, n439, n444, n449, n454, n459,
    n464, n469, n474, n479, n484, n489, n494, n499, n504, n509, n514, n519,
    n524, n529, n534, n539, n544, n549, n554, n559, n564, n569, n574, n579,
    n584, n589, n594, n599, n604, n609, n614, n619, n624, n629, n634, n639,
    n644, n649, n654, n659, n664, n669, n674, n679, n684, n689, n694, n699,
    n704, n709, n714, n719, n724, n729, n734, n739, n744, n749, n754, n759,
    n764, n769, n774, n779, n784, n789, n794, n799, n804, n809, n814, n819,
    n824;
  assign new_n483_ = ng24 & ng28;
  assign new_n484_1_ = ng28 & ~new_n483_;
  assign new_n485_ = ng24 & ~new_n483_;
  assign new_n486_ = ~new_n484_1_ & ~new_n485_;
  assign new_n487_ = ng18 & ng14;
  assign new_n488_ = ng18 & ~new_n487_;
  assign new_n489_1_ = ng14 & ~new_n487_;
  assign new_n490_ = ~new_n488_ & ~new_n489_1_;
  assign new_n491_ = ~new_n486_ & ~new_n490_;
  assign new_n492_ = ~new_n486_ & ~new_n491_;
  assign new_n493_ = ~new_n490_ & ~new_n491_;
  assign new_n494_1_ = ~new_n492_ & ~new_n493_;
  assign new_n495_ = ng6 & ng10;
  assign new_n496_ = ng10 & ~new_n495_;
  assign new_n497_ = ng6 & ~new_n495_;
  assign new_n498_ = ~new_n496_ & ~new_n497_;
  assign new_n499_1_ = ng1 & ng2;
  assign new_n500_ = ng2 & ~new_n499_1_;
  assign new_n501_ = ng1 & ~new_n499_1_;
  assign new_n502_ = ~new_n500_ & ~new_n501_;
  assign new_n503_ = ~new_n498_ & ~new_n502_;
  assign new_n504_1_ = ~new_n498_ & ~new_n503_;
  assign new_n505_ = ~new_n502_ & ~new_n503_;
  assign new_n506_ = ~new_n504_1_ & ~new_n505_;
  assign new_n507_ = ~new_n494_1_ & ~new_n506_;
  assign new_n508_ = ~new_n494_1_ & ~new_n507_;
  assign new_n509_1_ = ~new_n506_ & ~new_n507_;
  assign new_n510_ = ~new_n508_ & ~new_n509_1_;
  assign new_n511_ = ng48 & ~new_n510_;
  assign new_n512_ = ng48 & ~new_n511_;
  assign new_n513_ = ~new_n510_ & ~new_n511_;
  assign new_n514_1_ = ~new_n512_ & ~new_n513_;
  assign new_n515_ = ~pg41 & new_n514_1_;
  assign new_n516_ = ng676 & ~new_n515_;
  assign new_n517_ = ~pg22 & ng675;
  assign pg6282 = ~new_n516_ | ~new_n517_;
  assign new_n519_1_ = pg41 & ~pg6282;
  assign new_n520_ = ng25 & new_n519_1_;
  assign pg6360 = ~new_n519_1_ | new_n520_;
  assign new_n522_ = ng11 & new_n519_1_;
  assign pg6370 = ~new_n519_1_ | new_n522_;
  assign new_n524_1_ = ~ng489 & ng492;
  assign new_n525_ = ng496 & ~ng486;
  assign pg4809 = ~new_n524_1_ & ~new_n525_;
  assign new_n527_ = ng29 & new_n519_1_;
  assign pg6362 = ~new_n519_1_ | new_n527_;
  assign new_n529_1_ = ng15 & new_n519_1_;
  assign pg6372 = ~new_n519_1_ | new_n529_1_;
  assign new_n531_ = ng3 & new_n519_1_;
  assign pg6364 = ~new_n519_1_ | new_n531_;
  assign new_n533_ = ng7 & ng3;
  assign new_n534_1_ = ng3 & ~new_n533_;
  assign new_n535_ = ng7 & ~new_n533_;
  assign new_n536_ = ~new_n534_1_ & ~new_n535_;
  assign new_n537_ = ng15 & ng11;
  assign new_n538_ = ng11 & ~new_n537_;
  assign new_n539_1_ = ng15 & ~new_n537_;
  assign new_n540_ = ~new_n538_ & ~new_n539_1_;
  assign new_n541_ = ~new_n536_ & ~new_n540_;
  assign new_n542_ = ~new_n536_ & ~new_n541_;
  assign new_n543_ = ~new_n540_ & ~new_n541_;
  assign new_n544_1_ = ~new_n542_ & ~new_n543_;
  assign new_n545_ = ng25 & ng19;
  assign new_n546_ = ng19 & ~new_n545_;
  assign new_n547_ = ng25 & ~new_n545_;
  assign new_n548_ = ~new_n546_ & ~new_n547_;
  assign new_n549_1_ = ng33 & ng29;
  assign new_n550_ = ng29 & ~new_n549_1_;
  assign new_n551_ = ng33 & ~new_n549_1_;
  assign new_n552_ = ~new_n550_ & ~new_n551_;
  assign new_n553_ = ~new_n548_ & ~new_n552_;
  assign new_n554_1_ = ~new_n548_ & ~new_n553_;
  assign new_n555_ = ~new_n552_ & ~new_n553_;
  assign new_n556_ = ~new_n554_1_ & ~new_n555_;
  assign new_n557_ = ~new_n544_1_ & ~new_n556_;
  assign new_n558_ = ~new_n544_1_ & ~new_n557_;
  assign new_n559_1_ = ~new_n556_ & ~new_n557_;
  assign new_n560_ = ~new_n558_ & ~new_n559_1_;
  assign new_n561_ = new_n519_1_ & new_n560_;
  assign pg6284 = ~new_n519_1_ | new_n561_;
  assign new_n563_ = ng19 & new_n519_1_;
  assign pg6374 = ~new_n519_1_ | new_n563_;
  assign pg2584 = ~pg102 & pg89;
  assign new_n566_ = ~pg567 & ng638;
  assign pg4121 = ~ng638 | new_n566_;
  assign new_n568_ = ng33 & new_n519_1_;
  assign pg6366 = ~new_n519_1_ | new_n568_;
  assign new_n570_ = ng7 & new_n519_1_;
  assign pg6368 = ~new_n519_1_ | new_n570_;
  assign new_n572_ = ng689 & ng698;
  assign new_n573_ = ~ng688 & new_n572_;
  assign new_n574_1_ = ng685 & new_n573_;
  assign new_n575_ = pg702 & ng699;
  assign new_n576_ = ~pg41 & new_n575_;
  assign new_n577_ = new_n516_ & new_n576_;
  assign new_n578_ = ng697 & new_n574_1_;
  assign new_n579_1_ = ~ng683 & new_n577_;
  assign new_n580_ = new_n578_ & new_n579_1_;
  assign new_n581_ = ng677 & new_n580_;
  assign new_n582_ = ng197 & ~new_n580_;
  assign n159 = new_n581_ | new_n582_;
  assign new_n584_1_ = ng236 & ng516;
  assign new_n585_ = ng236 & ~new_n584_1_;
  assign new_n586_ = ng516 & ~new_n584_1_;
  assign new_n587_ = ~new_n585_ & ~new_n586_;
  assign new_n588_ = ng242 & ng520;
  assign new_n589_1_ = ng242 & ~new_n588_;
  assign new_n590_ = ng520 & ~new_n588_;
  assign new_n591_ = ~new_n589_1_ & ~new_n590_;
  assign new_n592_ = ng230 & ng512;
  assign new_n593_ = ng230 & ~new_n592_;
  assign new_n594_1_ = ng512 & ~new_n592_;
  assign new_n595_ = ~new_n593_ & ~new_n594_1_;
  assign new_n596_ = new_n587_ & new_n591_;
  assign new_n597_ = new_n595_ & new_n596_;
  assign new_n598_ = ng254 & ng528;
  assign new_n599_1_ = ng254 & ~new_n598_;
  assign new_n600_ = ng528 & ~new_n598_;
  assign new_n601_ = ~new_n599_1_ & ~new_n600_;
  assign new_n602_ = ng532 & ng260;
  assign new_n603_ = ng260 & ~new_n602_;
  assign new_n604_1_ = ng532 & ~new_n602_;
  assign new_n605_ = ~new_n603_ & ~new_n604_1_;
  assign new_n606_ = ng524 & ng290;
  assign new_n607_ = ng290 & ~new_n606_;
  assign new_n608_ = ng524 & ~new_n606_;
  assign new_n609_1_ = ~new_n607_ & ~new_n608_;
  assign new_n610_ = new_n601_ & new_n605_;
  assign new_n611_ = new_n609_1_ & new_n610_;
  assign new_n612_ = ng218 & ng504;
  assign new_n613_ = ng218 & ~new_n612_;
  assign new_n614_1_ = ng504 & ~new_n612_;
  assign new_n615_ = ~new_n613_ & ~new_n614_1_;
  assign new_n616_ = ng508 & ng286;
  assign new_n617_ = ng286 & ~new_n616_;
  assign new_n618_ = ng508 & ~new_n616_;
  assign new_n619_1_ = ~new_n617_ & ~new_n618_;
  assign new_n620_ = ng500 & ng212;
  assign new_n621_ = ng212 & ~new_n620_;
  assign new_n622_ = ng500 & ~new_n620_;
  assign new_n623_ = ~new_n621_ & ~new_n622_;
  assign new_n624_1_ = new_n615_ & new_n619_1_;
  assign new_n625_ = new_n623_ & new_n624_1_;
  assign new_n626_ = new_n597_ & new_n611_;
  assign new_n627_ = new_n625_ & new_n626_;
  assign new_n628_ = ~ng541 & new_n627_;
  assign new_n629_1_ = ~ng536 & new_n628_;
  assign new_n630_ = ng437 & new_n629_1_;
  assign new_n631_ = ng434 & ~new_n629_1_;
  assign n164 = new_n630_ | new_n631_;
  assign new_n633_ = ng683 & ng697;
  assign new_n634_1_ = ng266 & ~ng658;
  assign new_n635_ = ~ng658 & ng662;
  assign new_n636_ = ~new_n634_1_ & ~new_n635_;
  assign new_n637_ = pg41 & ~new_n636_;
  assign new_n638_ = new_n575_ & new_n637_;
  assign new_n639_1_ = new_n574_1_ & new_n633_;
  assign new_n640_ = ng682 & new_n638_;
  assign new_n641_ = new_n639_1_ & new_n640_;
  assign new_n642_ = ~ng677 & new_n641_;
  assign new_n643_ = ng441 & new_n642_;
  assign new_n644_1_ = ng689 & ~ng698;
  assign new_n645_ = new_n575_ & new_n635_;
  assign new_n646_ = pg41 & new_n645_;
  assign new_n647_ = new_n516_ & new_n646_;
  assign new_n648_ = ~ng687 & new_n644_1_;
  assign new_n649_1_ = new_n647_ & new_n648_;
  assign new_n650_ = ng677 & ng682;
  assign new_n651_ = ~ng677 & ng682;
  assign new_n652_ = ~new_n650_ & ~new_n651_;
  assign new_n653_ = new_n649_1_ & ~new_n652_;
  assign new_n654_1_ = ng677 & new_n641_;
  assign new_n655_ = ng422 & new_n654_1_;
  assign new_n656_ = ~ng685 & new_n573_;
  assign new_n657_ = ng697 & new_n647_;
  assign new_n658_ = new_n656_ & new_n657_;
  assign new_n659_1_ = ng682 & new_n658_;
  assign new_n660_ = ~new_n643_ & ~new_n653_;
  assign new_n661_ = ~new_n655_ & ~new_n659_1_;
  assign new_n662_ = new_n660_ & new_n661_;
  assign new_n663_ = ng688 & new_n572_;
  assign new_n664_1_ = ng691 & ng692;
  assign new_n665_ = new_n663_ & new_n664_1_;
  assign new_n666_ = ~ng680 & new_n638_;
  assign new_n667_ = new_n665_ & new_n666_;
  assign new_n668_ = pg559 & new_n667_;
  assign new_n669_1_ = ~ng683 & new_n638_;
  assign new_n670_ = new_n578_ & new_n669_1_;
  assign new_n671_ = ~new_n667_ & ~new_n670_;
  assign new_n672_ = ~new_n642_ & ~new_n649_1_;
  assign new_n673_ = ~new_n654_1_ & ~new_n658_;
  assign new_n674_1_ = new_n672_ & new_n673_;
  assign new_n675_ = ng694 & ~ng682;
  assign new_n676_ = new_n638_ & new_n675_;
  assign new_n677_ = new_n639_1_ & new_n676_;
  assign new_n678_ = ~ng694 & ~ng682;
  assign new_n679_1_ = new_n638_ & new_n678_;
  assign new_n680_ = new_n639_1_ & new_n679_1_;
  assign new_n681_ = ng677 & new_n680_;
  assign new_n682_ = ~ng677 & new_n680_;
  assign new_n683_ = ~ng691 & ~ng692;
  assign new_n684_1_ = new_n638_ & new_n663_;
  assign new_n685_ = ng680 & new_n683_;
  assign new_n686_ = new_n684_1_ & new_n685_;
  assign new_n687_ = ~ng692 & ~ng680;
  assign new_n688_ = ng691 & new_n663_;
  assign new_n689_1_ = new_n638_ & new_n687_;
  assign new_n690_ = new_n688_ & new_n689_1_;
  assign new_n691_ = new_n663_ & new_n687_;
  assign new_n692_ = ~ng691 & new_n638_;
  assign new_n693_ = new_n691_ & new_n692_;
  assign new_n694_1_ = ~new_n686_ & ~new_n690_;
  assign new_n695_ = ~new_n693_ & new_n694_1_;
  assign new_n696_ = ~new_n677_ & ~new_n681_;
  assign new_n697_ = ~new_n682_ & new_n695_;
  assign new_n698_ = new_n696_ & new_n697_;
  assign new_n699_1_ = ~ng697 & new_n573_;
  assign new_n700_ = ~ng685 & new_n647_;
  assign new_n701_ = new_n699_1_ & new_n700_;
  assign new_n702_ = ~ng689 & ~ng698;
  assign new_n703_ = ~ng687 & new_n702_;
  assign new_n704_1_ = ~ng688 & new_n647_;
  assign new_n705_ = new_n703_ & new_n704_1_;
  assign new_n706_ = ~ng688 & new_n702_;
  assign new_n707_ = ng687 & new_n647_;
  assign new_n708_ = new_n706_ & new_n707_;
  assign new_n709_1_ = ng687 & new_n644_1_;
  assign new_n710_ = new_n647_ & new_n709_1_;
  assign new_n711_ = ~new_n701_ & ~new_n705_;
  assign new_n712_ = ~new_n708_ & ~new_n710_;
  assign new_n713_ = new_n711_ & new_n712_;
  assign new_n714_1_ = new_n671_ & new_n674_1_;
  assign new_n715_ = new_n698_ & new_n714_1_;
  assign new_n716_ = new_n713_ & new_n715_;
  assign new_n717_ = ng520 & new_n681_;
  assign new_n718_ = ~new_n668_ & ~new_n716_;
  assign new_n719_1_ = ~new_n717_ & new_n718_;
  assign new_n720_ = ng682 & new_n701_;
  assign new_n721_ = ~ng197 & ng682;
  assign new_n722_ = ng205 & ng206;
  assign new_n723_ = ng204 & new_n722_;
  assign new_n724_1_ = ng207 & ng208;
  assign new_n725_ = new_n723_ & new_n724_1_;
  assign new_n726_ = ng209 & new_n725_;
  assign new_n727_ = ng209 & ~new_n726_;
  assign new_n728_ = new_n725_ & ~new_n726_;
  assign new_n729_1_ = ~new_n727_ & ~new_n728_;
  assign new_n730_ = ~ng210 & ~ng211;
  assign new_n731_ = ng208 & ng209;
  assign new_n732_ = ng208 & ~new_n731_;
  assign new_n733_ = ng209 & ~new_n731_;
  assign new_n734_1_ = ~new_n732_ & ~new_n733_;
  assign new_n735_ = ng205 & ng204;
  assign new_n736_ = ng206 & new_n735_;
  assign new_n737_ = ng207 & ng209;
  assign new_n738_ = ~ng208 & new_n737_;
  assign new_n739_1_ = new_n736_ & new_n738_;
  assign new_n740_ = ~new_n734_1_ & ~new_n739_1_;
  assign new_n741_ = ~ng471 & ~new_n740_;
  assign new_n742_ = new_n730_ & new_n741_;
  assign new_n743_ = new_n729_1_ & ~new_n742_;
  assign new_n744_1_ = ng471 & new_n740_;
  assign new_n745_ = ~ng471 & new_n740_;
  assign new_n746_ = ~new_n744_1_ & new_n745_;
  assign new_n747_ = new_n730_ & new_n746_;
  assign new_n748_ = ng209 & new_n724_1_;
  assign new_n749_1_ = ng205 & new_n748_;
  assign new_n750_ = ng204 & new_n749_1_;
  assign new_n751_ = ng206 & new_n750_;
  assign new_n752_ = ~new_n747_ & ~new_n751_;
  assign new_n753_ = ~new_n743_ & new_n752_;
  assign new_n754_1_ = ng197 & new_n753_;
  assign n754 = new_n721_ | new_n754_1_;
  assign new_n756_ = new_n705_ & n754;
  assign new_n757_ = ~ng269 & ng682;
  assign new_n758_ = ng278 & ng277;
  assign new_n759_1_ = ng276 & new_n758_;
  assign new_n760_ = ng279 & ng280;
  assign new_n761_ = new_n759_1_ & new_n760_;
  assign new_n762_ = ng281 & new_n761_;
  assign new_n763_ = ng281 & ~new_n762_;
  assign new_n764_1_ = new_n761_ & ~new_n762_;
  assign new_n765_ = ~new_n763_ & ~new_n764_1_;
  assign new_n766_ = ~ng282 & ~ng283;
  assign new_n767_ = ng281 & ng280;
  assign new_n768_ = ng280 & ~new_n767_;
  assign new_n769_1_ = ng281 & ~new_n767_;
  assign new_n770_ = ~new_n768_ & ~new_n769_1_;
  assign new_n771_ = ng277 & ng276;
  assign new_n772_ = ng278 & new_n771_;
  assign new_n773_ = ng279 & ng281;
  assign new_n774_1_ = ~ng280 & new_n773_;
  assign new_n775_ = new_n772_ & new_n774_1_;
  assign new_n776_ = ~new_n770_ & ~new_n775_;
  assign new_n777_ = ~ng478 & ~new_n776_;
  assign new_n778_ = new_n766_ & new_n777_;
  assign new_n779_1_ = new_n765_ & ~new_n778_;
  assign new_n780_ = ng478 & new_n776_;
  assign new_n781_ = ~ng478 & new_n776_;
  assign new_n782_ = ~new_n780_ & new_n781_;
  assign new_n783_ = new_n766_ & new_n782_;
  assign new_n784_1_ = ng281 & new_n760_;
  assign new_n785_ = ng277 & new_n784_1_;
  assign new_n786_ = ng276 & new_n785_;
  assign new_n787_ = ng278 & new_n786_;
  assign new_n788_ = ~new_n783_ & ~new_n787_;
  assign new_n789_1_ = ~new_n779_1_ & new_n788_;
  assign new_n790_ = ng269 & new_n789_1_;
  assign n579 = new_n757_ | new_n790_;
  assign new_n792_ = new_n708_ & n579;
  assign new_n793_ = ~new_n652_ & new_n710_;
  assign new_n794_1_ = ~new_n720_ & ~new_n756_;
  assign new_n795_ = ~new_n792_ & ~new_n793_;
  assign new_n796_ = new_n794_1_ & new_n795_;
  assign new_n797_ = new_n662_ & new_n719_1_;
  assign n169 = ~new_n796_ | ~new_n797_;
  assign new_n799_1_ = ~ng197 & ng691;
  assign new_n800_ = ng205 & ~new_n735_;
  assign new_n801_ = ng204 & ~new_n735_;
  assign new_n802_ = ~new_n800_ & ~new_n801_;
  assign new_n803_ = new_n752_ & ~new_n802_;
  assign new_n804_1_ = ~new_n742_ & new_n803_;
  assign new_n805_ = ng197 & new_n804_1_;
  assign n174 = new_n799_1_ | new_n805_;
  assign n179 = pg45 & ~ng266;
  assign new_n808_ = ~ng197 & ng677;
  assign new_n809_1_ = ~ng204 & ~new_n742_;
  assign new_n810_ = new_n752_ & new_n809_1_;
  assign new_n811_ = ng197 & new_n810_;
  assign n184 = new_n808_ | new_n811_;
  assign new_n813_ = new_n577_ & new_n678_;
  assign new_n814_1_ = new_n639_1_ & new_n813_;
  assign new_n815_ = ng677 & new_n814_1_;
  assign new_n816_ = ng683 & new_n815_;
  assign new_n817_ = ng524 & ~new_n815_;
  assign n189 = new_n816_ | new_n817_;
  assign n199 = pg45 & ~ng658;
  assign new_n820_ = ng410 & new_n629_1_;
  assign new_n821_ = ng414 & ~new_n629_1_;
  assign n209 = new_n820_ | new_n821_;
  assign new_n823_ = new_n519_1_ & pg6364;
  assign new_n824_1_ = ng3 & ~new_n519_1_;
  assign n214 = new_n823_ | new_n824_1_;
  assign new_n826_ = pg567 & ng598;
  assign new_n827_ = ng598 & ~new_n826_;
  assign new_n828_ = pg567 & ~new_n826_;
  assign new_n829_ = ~new_n827_ & ~new_n828_;
  assign n219 = ng638 & ~new_n829_;
  assign new_n831_ = ng610 & ng602;
  assign new_n832_ = ng613 & new_n831_;
  assign new_n833_ = ng616 & new_n832_;
  assign new_n834_ = ng619 & new_n833_;
  assign new_n835_ = ng622 & new_n834_;
  assign new_n836_ = ng625 & new_n835_;
  assign new_n837_ = ng628 & new_n836_;
  assign new_n838_ = ng631 & new_n837_;
  assign new_n839_ = ng578 & new_n838_;
  assign new_n840_ = ng582 & new_n839_;
  assign new_n841_ = ng586 & new_n840_;
  assign new_n842_ = ng574 & new_n841_;
  assign new_n843_ = ng590 & new_n842_;
  assign new_n844_ = ng594 & new_n843_;
  assign new_n845_ = pg639 & ~new_n844_;
  assign new_n846_ = ng578 & ~new_n839_;
  assign new_n847_ = new_n838_ & ~new_n839_;
  assign new_n848_ = ~new_n846_ & ~new_n847_;
  assign n224 = new_n845_ & ~new_n848_;
  assign new_n850_ = ng402 & new_n629_1_;
  assign new_n851_ = ng406 & ~new_n629_1_;
  assign n229 = new_n850_ | new_n851_;
  assign new_n853_ = ng582 & ~new_n840_;
  assign new_n854_ = new_n839_ & ~new_n840_;
  assign new_n855_ = ~new_n853_ & ~new_n854_;
  assign n234 = new_n845_ & ~new_n855_;
  assign new_n857_ = ng204 & ng677;
  assign new_n858_ = ~ng204 & ng691;
  assign new_n859_ = ~new_n857_ & ~new_n858_;
  assign new_n860_ = ng205 & new_n859_;
  assign new_n861_ = ng204 & ng692;
  assign new_n862_ = ~ng204 & ng680;
  assign new_n863_ = ~new_n861_ & ~new_n862_;
  assign new_n864_ = ~ng205 & new_n863_;
  assign new_n865_ = ~new_n860_ & ~new_n864_;
  assign new_n866_ = ng206 & new_n865_;
  assign new_n867_ = ng204 & ng694;
  assign new_n868_ = ~ng204 & ng682;
  assign new_n869_ = ~new_n867_ & ~new_n868_;
  assign new_n870_ = ng205 & new_n869_;
  assign new_n871_ = ng204 & ng683;
  assign new_n872_ = ~ng204 & ng697;
  assign new_n873_ = ~new_n871_ & ~new_n872_;
  assign new_n874_ = ~ng205 & new_n873_;
  assign new_n875_ = ~new_n870_ & ~new_n874_;
  assign new_n876_ = ~ng206 & new_n875_;
  assign new_n877_ = ~new_n866_ & ~new_n876_;
  assign new_n878_ = ng207 & new_n877_;
  assign new_n879_ = ~ng207 & new_n877_;
  assign new_n880_ = ~new_n878_ & ~new_n879_;
  assign new_n881_ = ng471 & new_n880_;
  assign new_n882_ = new_n880_ & ~new_n881_;
  assign new_n883_ = ng471 & ~new_n881_;
  assign new_n884_ = ~new_n882_ & ~new_n883_;
  assign new_n885_ = ng210 & ~ng211;
  assign new_n886_ = new_n734_1_ & ~new_n884_;
  assign new_n887_ = new_n885_ & new_n886_;
  assign new_n888_ = new_n751_ & ~new_n887_;
  assign new_n889_ = new_n885_ & new_n888_;
  assign new_n890_ = new_n740_ & ~new_n744_1_;
  assign new_n891_ = ng471 & ~new_n744_1_;
  assign new_n892_ = ~new_n890_ & ~new_n891_;
  assign new_n893_ = ~new_n734_1_ & ~new_n892_;
  assign new_n894_ = new_n885_ & new_n893_;
  assign new_n895_ = ~new_n747_ & ~new_n894_;
  assign new_n896_ = ~new_n751_ & new_n887_;
  assign new_n897_ = ng210 & ng211;
  assign new_n898_ = ~new_n892_ & new_n897_;
  assign new_n899_ = ~new_n734_1_ & new_n898_;
  assign new_n900_ = ~new_n884_ & new_n897_;
  assign new_n901_ = new_n734_1_ & new_n900_;
  assign new_n902_ = ~new_n899_ & ~new_n901_;
  assign new_n903_ = ~new_n751_ & ~new_n902_;
  assign new_n904_ = ~new_n896_ & ~new_n903_;
  assign new_n905_ = ng210 & new_n895_;
  assign new_n906_ = new_n904_ & new_n905_;
  assign new_n907_ = ~ng210 & ng211;
  assign new_n908_ = new_n751_ & new_n907_;
  assign new_n909_ = new_n751_ & ~new_n902_;
  assign new_n910_ = new_n751_ & new_n887_;
  assign new_n911_ = ~new_n908_ & ~new_n909_;
  assign new_n912_ = ~new_n742_ & ~new_n910_;
  assign new_n913_ = new_n911_ & new_n912_;
  assign new_n914_ = ~new_n889_ & ~new_n906_;
  assign new_n915_ = new_n913_ & new_n914_;
  assign new_n916_ = ng211 & new_n895_;
  assign new_n917_ = new_n913_ & new_n916_;
  assign new_n918_ = ~new_n889_ & ~new_n917_;
  assign new_n919_ = new_n904_ & new_n918_;
  assign n244 = new_n915_ | new_n919_;
  assign new_n921_ = new_n627_ & ~new_n919_;
  assign new_n922_ = ng548 & ~new_n627_;
  assign n249 = new_n921_ | new_n922_;
  assign new_n924_ = ng677 & ng276;
  assign new_n925_ = ng691 & ~ng276;
  assign new_n926_ = ~new_n924_ & ~new_n925_;
  assign new_n927_ = ng277 & new_n926_;
  assign new_n928_ = ng692 & ng276;
  assign new_n929_ = ng680 & ~ng276;
  assign new_n930_ = ~new_n928_ & ~new_n929_;
  assign new_n931_ = ~ng277 & new_n930_;
  assign new_n932_ = ~new_n927_ & ~new_n931_;
  assign new_n933_ = ng278 & new_n932_;
  assign new_n934_ = ng694 & ng276;
  assign new_n935_ = ~ng276 & ng682;
  assign new_n936_ = ~new_n934_ & ~new_n935_;
  assign new_n937_ = ng277 & new_n936_;
  assign new_n938_ = ng276 & ng683;
  assign new_n939_ = ~ng276 & ng697;
  assign new_n940_ = ~new_n938_ & ~new_n939_;
  assign new_n941_ = ~ng277 & new_n940_;
  assign new_n942_ = ~new_n937_ & ~new_n941_;
  assign new_n943_ = ~ng278 & new_n942_;
  assign new_n944_ = ~new_n933_ & ~new_n943_;
  assign new_n945_ = ng279 & new_n944_;
  assign new_n946_ = ~ng279 & new_n944_;
  assign new_n947_ = ~new_n945_ & ~new_n946_;
  assign new_n948_ = ng478 & new_n947_;
  assign new_n949_ = new_n947_ & ~new_n948_;
  assign new_n950_ = ng478 & ~new_n948_;
  assign new_n951_ = ~new_n949_ & ~new_n950_;
  assign new_n952_ = ng282 & ~ng283;
  assign new_n953_ = new_n770_ & ~new_n951_;
  assign new_n954_ = new_n952_ & new_n953_;
  assign new_n955_ = new_n787_ & ~new_n954_;
  assign new_n956_ = new_n952_ & new_n955_;
  assign new_n957_ = new_n776_ & ~new_n780_;
  assign new_n958_ = ng478 & ~new_n780_;
  assign new_n959_ = ~new_n957_ & ~new_n958_;
  assign new_n960_ = ~new_n770_ & ~new_n959_;
  assign new_n961_ = new_n952_ & new_n960_;
  assign new_n962_ = ~new_n783_ & ~new_n961_;
  assign new_n963_ = ~new_n787_ & new_n954_;
  assign new_n964_ = ng282 & ng283;
  assign new_n965_ = ~new_n959_ & new_n964_;
  assign new_n966_ = ~new_n770_ & new_n965_;
  assign new_n967_ = ~new_n951_ & new_n964_;
  assign new_n968_ = new_n770_ & new_n967_;
  assign new_n969_ = ~new_n966_ & ~new_n968_;
  assign new_n970_ = ~new_n787_ & ~new_n969_;
  assign new_n971_ = ~new_n963_ & ~new_n970_;
  assign new_n972_ = ng282 & new_n962_;
  assign new_n973_ = new_n971_ & new_n972_;
  assign new_n974_ = ~ng282 & ng283;
  assign new_n975_ = new_n787_ & new_n974_;
  assign new_n976_ = new_n787_ & ~new_n969_;
  assign new_n977_ = new_n787_ & new_n954_;
  assign new_n978_ = ~new_n975_ & ~new_n976_;
  assign new_n979_ = ~new_n778_ & ~new_n977_;
  assign new_n980_ = new_n978_ & new_n979_;
  assign new_n981_ = ~new_n956_ & ~new_n973_;
  assign new_n982_ = new_n980_ & new_n981_;
  assign new_n983_ = ng283 & new_n962_;
  assign new_n984_ = new_n980_ & new_n983_;
  assign new_n985_ = ~new_n956_ & ~new_n984_;
  assign new_n986_ = new_n971_ & new_n985_;
  assign n254 = new_n982_ | new_n986_;
  assign new_n988_ = ng418 & new_n629_1_;
  assign new_n989_ = ng422 & ~new_n629_1_;
  assign n264 = new_n988_ | new_n989_;
  assign new_n991_ = ng677 & new_n815_;
  assign new_n992_ = ng500 & ~new_n815_;
  assign n269 = new_n991_ | new_n992_;
  assign new_n994_ = ng445 & new_n642_;
  assign new_n995_ = ng694 & ng677;
  assign new_n996_ = ng694 & ~ng677;
  assign new_n997_ = ~new_n995_ & ~new_n996_;
  assign new_n998_ = new_n649_1_ & ~new_n997_;
  assign new_n999_ = ng418 & new_n654_1_;
  assign new_n1000_ = ng694 & new_n658_;
  assign new_n1001_ = ~new_n994_ & ~new_n998_;
  assign new_n1002_ = ~new_n999_ & ~new_n1000_;
  assign new_n1003_ = new_n1001_ & new_n1002_;
  assign new_n1004_ = pg560 & new_n667_;
  assign new_n1005_ = ng516 & new_n681_;
  assign new_n1006_ = ~new_n716_ & ~new_n1004_;
  assign new_n1007_ = ~new_n1005_ & new_n1006_;
  assign new_n1008_ = ng694 & new_n701_;
  assign new_n1009_ = ~ng197 & ng694;
  assign new_n1010_ = ng207 & new_n723_;
  assign new_n1011_ = ng208 & new_n1010_;
  assign new_n1012_ = ng208 & ~new_n1011_;
  assign new_n1013_ = new_n1010_ & ~new_n1011_;
  assign new_n1014_ = ~new_n1012_ & ~new_n1013_;
  assign new_n1015_ = ~new_n742_ & new_n1014_;
  assign new_n1016_ = new_n752_ & new_n1015_;
  assign new_n1017_ = ng197 & ~new_n1016_;
  assign n509 = new_n1009_ | new_n1017_;
  assign new_n1019_ = new_n705_ & n509;
  assign new_n1020_ = ng694 & ~ng269;
  assign new_n1021_ = ng279 & new_n759_1_;
  assign new_n1022_ = ng280 & new_n1021_;
  assign new_n1023_ = ng280 & ~new_n1022_;
  assign new_n1024_ = new_n1021_ & ~new_n1022_;
  assign new_n1025_ = ~new_n1023_ & ~new_n1024_;
  assign new_n1026_ = ~new_n778_ & new_n1025_;
  assign new_n1027_ = new_n788_ & new_n1026_;
  assign new_n1028_ = ng269 & ~new_n1027_;
  assign n684 = new_n1020_ | new_n1028_;
  assign new_n1030_ = new_n708_ & n684;
  assign new_n1031_ = new_n710_ & ~new_n997_;
  assign new_n1032_ = ~new_n1008_ & ~new_n1019_;
  assign new_n1033_ = ~new_n1030_ & ~new_n1031_;
  assign new_n1034_ = new_n1032_ & new_n1033_;
  assign new_n1035_ = new_n1003_ & new_n1007_;
  assign n274 = ~new_n1034_ | ~new_n1035_;
  assign new_n1037_ = ~ng677 & new_n814_1_;
  assign new_n1038_ = ng677 & new_n1037_;
  assign new_n1039_ = ng532 & ~new_n1037_;
  assign n279 = new_n1038_ | new_n1039_;
  assign new_n1041_ = ~ng197 & ng683;
  assign new_n1042_ = ng197 & ~new_n915_;
  assign n284 = new_n1041_ | new_n1042_;
  assign new_n1044_ = ng680 & new_n815_;
  assign new_n1045_ = ng512 & ~new_n815_;
  assign n299 = new_n1044_ | new_n1045_;
  assign new_n1047_ = ng691 & new_n1037_;
  assign new_n1048_ = ng465 & ~new_n1037_;
  assign n304 = new_n1047_ | new_n1048_;
  assign new_n1050_ = pg39 & pg40;
  assign new_n1051_ = pg40 & ~new_n1050_;
  assign new_n1052_ = pg39 & ~new_n1050_;
  assign new_n1053_ = ~new_n1051_ & ~new_n1052_;
  assign new_n1054_ = pg38 & pg37;
  assign new_n1055_ = pg38 & ~new_n1054_;
  assign new_n1056_ = pg37 & ~new_n1054_;
  assign new_n1057_ = ~new_n1055_ & ~new_n1056_;
  assign new_n1058_ = pg32 & pg36;
  assign new_n1059_ = pg36 & ~new_n1058_;
  assign new_n1060_ = pg32 & ~new_n1058_;
  assign new_n1061_ = ~new_n1059_ & ~new_n1060_;
  assign new_n1062_ = ~new_n1057_ & ~new_n1061_;
  assign new_n1063_ = ~new_n1057_ & ~new_n1062_;
  assign new_n1064_ = ~new_n1061_ & ~new_n1062_;
  assign new_n1065_ = ~new_n1063_ & ~new_n1064_;
  assign new_n1066_ = ~new_n1053_ & ~new_n1065_;
  assign new_n1067_ = ~new_n1053_ & ~new_n1066_;
  assign new_n1068_ = ~new_n1065_ & ~new_n1066_;
  assign new_n1069_ = ~new_n1067_ & ~new_n1068_;
  assign new_n1070_ = ~new_n510_ & ~new_n1069_;
  assign new_n1071_ = ~new_n1069_ & ~new_n1070_;
  assign new_n1072_ = ~new_n510_ & ~new_n1070_;
  assign new_n1073_ = ~new_n1071_ & ~new_n1072_;
  assign new_n1074_ = ng48 & ~new_n1073_;
  assign new_n1075_ = ng48 & ~new_n1074_;
  assign new_n1076_ = ~new_n1073_ & ~new_n1074_;
  assign n309 = new_n1075_ | new_n1076_;
  assign new_n1078_ = ng622 & ~new_n835_;
  assign new_n1079_ = new_n834_ & ~new_n835_;
  assign new_n1080_ = ~new_n1078_ & ~new_n1079_;
  assign n314 = pg639 & ~new_n1080_;
  assign new_n1082_ = ng692 & ~ng269;
  assign new_n1083_ = ng278 & ~new_n772_;
  assign new_n1084_ = new_n771_ & ~new_n772_;
  assign new_n1085_ = ~new_n1083_ & ~new_n1084_;
  assign new_n1086_ = new_n788_ & ~new_n1085_;
  assign new_n1087_ = ~new_n778_ & new_n1086_;
  assign new_n1088_ = ng269 & new_n1087_;
  assign n319 = new_n1082_ | new_n1088_;
  assign new_n1090_ = ng430 & new_n629_1_;
  assign new_n1091_ = ng461 & ~new_n629_1_;
  assign n324 = new_n1090_ | new_n1091_;
  assign new_n1093_ = ng634 & new_n826_;
  assign new_n1094_ = ng642 & new_n1093_;
  assign new_n1095_ = ng606 & new_n1094_;
  assign new_n1096_ = ng646 & new_n1095_;
  assign new_n1097_ = ng650 & new_n1096_;
  assign new_n1098_ = ng650 & ~new_n1097_;
  assign new_n1099_ = new_n1096_ & ~new_n1097_;
  assign new_n1100_ = ~new_n1098_ & ~new_n1099_;
  assign n329 = ng638 & ~new_n1100_;
  assign new_n1102_ = ~new_n670_ & ~new_n686_;
  assign new_n1103_ = ~new_n667_ & ~new_n677_;
  assign new_n1104_ = new_n1102_ & new_n1103_;
  assign new_n1105_ = ~new_n682_ & ~new_n693_;
  assign new_n1106_ = ~new_n681_ & ~new_n690_;
  assign new_n1107_ = new_n1105_ & new_n1106_;
  assign new_n1108_ = new_n674_1_ & new_n1104_;
  assign new_n1109_ = new_n1107_ & new_n1108_;
  assign new_n1110_ = new_n713_ & new_n1109_;
  assign new_n1111_ = ng672 & new_n686_;
  assign new_n1112_ = ng269 & new_n670_;
  assign new_n1113_ = pg563 & new_n667_;
  assign new_n1114_ = ng548 & new_n677_;
  assign new_n1115_ = ~new_n1111_ & ~new_n1112_;
  assign new_n1116_ = ~new_n1113_ & ~new_n1114_;
  assign new_n1117_ = new_n1115_ & new_n1116_;
  assign new_n1118_ = ng457 & new_n642_;
  assign new_n1119_ = ng691 & ng677;
  assign new_n1120_ = ng691 & ~ng677;
  assign new_n1121_ = ~new_n1119_ & ~new_n1120_;
  assign new_n1122_ = new_n649_1_ & ~new_n1121_;
  assign new_n1123_ = ng406 & new_n654_1_;
  assign new_n1124_ = ng691 & new_n658_;
  assign new_n1125_ = ~new_n1118_ & ~new_n1122_;
  assign new_n1126_ = ~new_n1123_ & ~new_n1124_;
  assign new_n1127_ = new_n1125_ & new_n1126_;
  assign new_n1128_ = ng465 & new_n682_;
  assign new_n1129_ = ng492 & new_n693_;
  assign new_n1130_ = ng504 & new_n681_;
  assign new_n1131_ = ~ng489 & new_n690_;
  assign new_n1132_ = ~new_n1128_ & ~new_n1129_;
  assign new_n1133_ = ~new_n1130_ & ~new_n1131_;
  assign new_n1134_ = new_n1132_ & new_n1133_;
  assign new_n1135_ = ng691 & new_n701_;
  assign new_n1136_ = new_n705_ & n174;
  assign new_n1137_ = ng691 & ~ng269;
  assign new_n1138_ = ng277 & ~new_n771_;
  assign new_n1139_ = ng276 & ~new_n771_;
  assign new_n1140_ = ~new_n1138_ & ~new_n1139_;
  assign new_n1141_ = new_n788_ & ~new_n1140_;
  assign new_n1142_ = ~new_n778_ & new_n1141_;
  assign new_n1143_ = ng269 & new_n1142_;
  assign n369 = new_n1137_ | new_n1143_;
  assign new_n1145_ = new_n708_ & n369;
  assign new_n1146_ = new_n710_ & ~new_n1121_;
  assign new_n1147_ = ~new_n1135_ & ~new_n1136_;
  assign new_n1148_ = ~new_n1145_ & ~new_n1146_;
  assign new_n1149_ = new_n1147_ & new_n1148_;
  assign new_n1150_ = new_n1117_ & new_n1127_;
  assign new_n1151_ = new_n1134_ & new_n1149_;
  assign new_n1152_ = new_n1150_ & new_n1151_;
  assign n334 = new_n1110_ | ~new_n1152_;
  assign new_n1154_ = new_n519_1_ & pg6360;
  assign new_n1155_ = ng25 & ~new_n519_1_;
  assign n339 = new_n1154_ | new_n1155_;
  assign new_n1157_ = ng692 & new_n815_;
  assign new_n1158_ = ng508 & ~new_n815_;
  assign n344 = new_n1157_ | new_n1158_;
  assign new_n1160_ = new_n519_1_ & pg6362;
  assign new_n1161_ = ng29 & ~new_n519_1_;
  assign n364 = new_n1160_ | new_n1161_;
  assign new_n1163_ = ng457 & new_n629_1_;
  assign new_n1164_ = ng453 & ~new_n629_1_;
  assign n374 = new_n1163_ | new_n1164_;
  assign new_n1166_ = ng449 & new_n629_1_;
  assign new_n1167_ = ng445 & ~new_n629_1_;
  assign n379 = new_n1166_ | new_n1167_;
  assign new_n1169_ = new_n519_1_ & pg6368;
  assign new_n1170_ = ng7 & ~new_n519_1_;
  assign n384 = new_n1169_ | new_n1170_;
  assign new_n1172_ = ~ng269 & ng680;
  assign new_n1173_ = ng279 & ~new_n1021_;
  assign new_n1174_ = new_n759_1_ & ~new_n1021_;
  assign new_n1175_ = ~new_n1173_ & ~new_n1174_;
  assign new_n1176_ = new_n788_ & new_n1175_;
  assign new_n1177_ = ~new_n778_ & ~new_n1176_;
  assign new_n1178_ = ng269 & new_n1177_;
  assign n389 = new_n1172_ | new_n1178_;
  assign new_n1180_ = ng594 & ~new_n844_;
  assign new_n1181_ = new_n843_ & ~new_n844_;
  assign new_n1182_ = ~new_n1180_ & ~new_n1181_;
  assign n394 = new_n845_ & ~new_n1182_;
  assign new_n1184_ = ng691 & new_n580_;
  assign new_n1185_ = ng269 & ~new_n580_;
  assign n399 = new_n1184_ | new_n1185_;
  assign new_n1187_ = ng692 & new_n580_;
  assign new_n1188_ = ng293 & ~new_n580_;
  assign n404 = new_n1187_ | new_n1188_;
  assign new_n1190_ = ng628 & ~new_n837_;
  assign new_n1191_ = new_n836_ & ~new_n837_;
  assign new_n1192_ = ~new_n1190_ & ~new_n1191_;
  assign n409 = pg639 & ~new_n1192_;
  assign new_n1194_ = ng574 & ~new_n842_;
  assign new_n1195_ = new_n841_ & ~new_n842_;
  assign new_n1196_ = ~new_n1194_ & ~new_n1195_;
  assign new_n1197_ = new_n845_ & ~new_n1196_;
  assign n424 = ~new_n845_ | new_n1197_;
  assign new_n1199_ = ~pg22 & ~pg41;
  assign new_n1200_ = new_n514_1_ & new_n1199_;
  assign n439 = ng672 | new_n1200_;
  assign new_n1202_ = ~ng197 & ng680;
  assign new_n1203_ = ng207 & ~new_n1010_;
  assign new_n1204_ = new_n723_ & ~new_n1010_;
  assign new_n1205_ = ~new_n1203_ & ~new_n1204_;
  assign new_n1206_ = new_n752_ & new_n1205_;
  assign new_n1207_ = ~new_n742_ & ~new_n1206_;
  assign new_n1208_ = ng197 & new_n1207_;
  assign n449 = new_n1202_ | new_n1208_;
  assign new_n1210_ = ng445 & new_n629_1_;
  assign new_n1211_ = ng441 & ~new_n629_1_;
  assign n454 = new_n1210_ | new_n1211_;
  assign new_n1213_ = new_n519_1_ & pg6370;
  assign new_n1214_ = ng11 & ~new_n519_1_;
  assign n459 = new_n1213_ | new_n1214_;
  assign new_n1216_ = ng616 & ~new_n833_;
  assign new_n1217_ = new_n832_ & ~new_n833_;
  assign new_n1218_ = ~new_n1216_ & ~new_n1217_;
  assign n474 = pg639 & ~new_n1218_;
  assign new_n1220_ = new_n627_ & ~new_n986_;
  assign new_n1221_ = ng554 & ~new_n627_;
  assign n479 = new_n1220_ | new_n1221_;
  assign new_n1223_ = ng625 & ~new_n836_;
  assign new_n1224_ = new_n835_ & ~new_n836_;
  assign new_n1225_ = ~new_n1223_ & ~new_n1224_;
  assign n484 = pg639 & ~new_n1225_;
  assign new_n1227_ = ng422 & new_n629_1_;
  assign new_n1228_ = ng426 & ~new_n629_1_;
  assign n489 = new_n1227_ | new_n1228_;
  assign new_n1230_ = ng465 & ng478;
  assign new_n1231_ = ~ng465 & ng471;
  assign new_n1232_ = ~new_n1230_ & ~new_n1231_;
  assign new_n1233_ = new_n629_1_ & ~new_n1232_;
  assign new_n1234_ = ng402 & ~new_n629_1_;
  assign n494 = new_n1233_ | new_n1234_;
  assign new_n1236_ = ~new_n903_ & ~new_n909_;
  assign n504 = ng496 | ~new_n1236_;
  assign new_n1238_ = ng634 & ~new_n1093_;
  assign new_n1239_ = new_n826_ & ~new_n1093_;
  assign new_n1240_ = ~new_n1238_ & ~new_n1239_;
  assign n514 = ng638 & ~new_n1240_;
  assign new_n1242_ = ng414 & new_n629_1_;
  assign new_n1243_ = ng418 & ~new_n629_1_;
  assign n519 = new_n1242_ | new_n1243_;
  assign new_n1245_ = new_n519_1_ & pg6284;
  assign new_n1246_ = ~new_n519_1_ & new_n560_;
  assign n529 = new_n1245_ | new_n1246_;
  assign new_n1248_ = ng677 & ~ng269;
  assign new_n1249_ = ~ng276 & ~new_n778_;
  assign new_n1250_ = new_n788_ & new_n1249_;
  assign new_n1251_ = ng269 & new_n1250_;
  assign n534 = new_n1248_ | new_n1251_;
  assign new_n1253_ = ng453 & new_n629_1_;
  assign new_n1254_ = ng449 & ~new_n629_1_;
  assign n539 = new_n1253_ | new_n1254_;
  assign new_n1256_ = ng590 & ~new_n843_;
  assign new_n1257_ = new_n842_ & ~new_n843_;
  assign new_n1258_ = ~new_n1256_ & ~new_n1257_;
  assign new_n1259_ = new_n845_ & ~new_n1258_;
  assign n549 = ~new_n845_ | new_n1259_;
  assign new_n1261_ = ng441 & new_n629_1_;
  assign new_n1262_ = ng437 & ~new_n629_1_;
  assign n554 = new_n1261_ | new_n1262_;
  assign new_n1264_ = ng697 & new_n815_;
  assign new_n1265_ = ng528 & ~new_n815_;
  assign n559 = new_n1264_ | new_n1265_;
  assign new_n1267_ = new_n627_ & ~new_n982_;
  assign new_n1268_ = ng551 & ~new_n627_;
  assign n569 = new_n1267_ | new_n1268_;
  assign new_n1270_ = ng426 & new_n629_1_;
  assign new_n1271_ = ng430 & ~new_n629_1_;
  assign n584 = new_n1270_ | new_n1271_;
  assign new_n1273_ = new_n627_ & ~new_n915_;
  assign new_n1274_ = ng545 & ~new_n627_;
  assign n594 = new_n1273_ | new_n1274_;
  assign new_n1276_ = ng669 & new_n686_;
  assign new_n1277_ = ng197 & new_n670_;
  assign new_n1278_ = pg564 & new_n667_;
  assign new_n1279_ = ng545 & new_n677_;
  assign new_n1280_ = ~new_n1276_ & ~new_n1277_;
  assign new_n1281_ = ~new_n1278_ & ~new_n1279_;
  assign new_n1282_ = new_n1280_ & new_n1281_;
  assign new_n1283_ = ng461 & new_n642_;
  assign new_n1284_ = ng677 & new_n649_1_;
  assign new_n1285_ = ng402 & new_n654_1_;
  assign new_n1286_ = ng677 & new_n658_;
  assign new_n1287_ = ~new_n1283_ & ~new_n1284_;
  assign new_n1288_ = ~new_n1285_ & ~new_n1286_;
  assign new_n1289_ = new_n1287_ & new_n1288_;
  assign new_n1290_ = ng532 & new_n682_;
  assign new_n1291_ = ng496 & new_n693_;
  assign new_n1292_ = ng500 & new_n681_;
  assign new_n1293_ = ~ng486 & new_n690_;
  assign new_n1294_ = ~new_n1290_ & ~new_n1291_;
  assign new_n1295_ = ~new_n1292_ & ~new_n1293_;
  assign new_n1296_ = new_n1294_ & new_n1295_;
  assign new_n1297_ = ng677 & new_n701_;
  assign new_n1298_ = new_n705_ & n184;
  assign new_n1299_ = new_n708_ & n534;
  assign new_n1300_ = ng677 & new_n710_;
  assign new_n1301_ = ~new_n1297_ & ~new_n1298_;
  assign new_n1302_ = ~new_n1299_ & ~new_n1300_;
  assign new_n1303_ = new_n1301_ & new_n1302_;
  assign new_n1304_ = new_n1282_ & new_n1289_;
  assign new_n1305_ = new_n1296_ & new_n1303_;
  assign new_n1306_ = new_n1304_ & new_n1305_;
  assign n604 = new_n1110_ | ~new_n1306_;
  assign new_n1308_ = pg561 & new_n667_;
  assign new_n1309_ = ~new_n716_ & ~new_n1308_;
  assign new_n1310_ = ng449 & new_n642_;
  assign new_n1311_ = ng677 & ng680;
  assign new_n1312_ = ~ng677 & ng680;
  assign new_n1313_ = ~new_n1311_ & ~new_n1312_;
  assign new_n1314_ = new_n649_1_ & ~new_n1313_;
  assign new_n1315_ = ng414 & new_n654_1_;
  assign new_n1316_ = ng680 & new_n658_;
  assign new_n1317_ = ~new_n1310_ & ~new_n1314_;
  assign new_n1318_ = ~new_n1315_ & ~new_n1316_;
  assign new_n1319_ = new_n1317_ & new_n1318_;
  assign new_n1320_ = ng297 & new_n670_;
  assign new_n1321_ = ng541 & new_n682_;
  assign new_n1322_ = ng554 & new_n677_;
  assign new_n1323_ = ng512 & new_n681_;
  assign new_n1324_ = ~new_n1320_ & ~new_n1321_;
  assign new_n1325_ = ~new_n1322_ & ~new_n1323_;
  assign new_n1326_ = new_n1324_ & new_n1325_;
  assign new_n1327_ = ng680 & new_n701_;
  assign new_n1328_ = new_n705_ & n449;
  assign new_n1329_ = new_n708_ & n389;
  assign new_n1330_ = new_n710_ & ~new_n1313_;
  assign new_n1331_ = ~new_n1327_ & ~new_n1328_;
  assign new_n1332_ = ~new_n1329_ & ~new_n1330_;
  assign new_n1333_ = new_n1331_ & new_n1332_;
  assign new_n1334_ = new_n1309_ & new_n1319_;
  assign new_n1335_ = new_n1326_ & new_n1333_;
  assign n609 = ~new_n1334_ | ~new_n1335_;
  assign new_n1337_ = ng406 & new_n629_1_;
  assign new_n1338_ = ng410 & ~new_n629_1_;
  assign n614 = new_n1337_ | new_n1338_;
  assign new_n1340_ = ng654 & new_n1097_;
  assign new_n1341_ = ng654 & ~new_n1340_;
  assign new_n1342_ = new_n1097_ & ~new_n1340_;
  assign new_n1343_ = ~new_n1341_ & ~new_n1342_;
  assign n619 = ng638 & ~new_n1343_;
  assign new_n1345_ = pg562 & new_n667_;
  assign new_n1346_ = ~new_n716_ & ~new_n1345_;
  assign new_n1347_ = ng453 & new_n642_;
  assign new_n1348_ = ng677 & ng692;
  assign new_n1349_ = ~ng677 & ng692;
  assign new_n1350_ = ~new_n1348_ & ~new_n1349_;
  assign new_n1351_ = new_n649_1_ & ~new_n1350_;
  assign new_n1352_ = ng410 & new_n654_1_;
  assign new_n1353_ = ng692 & new_n658_;
  assign new_n1354_ = ~new_n1347_ & ~new_n1351_;
  assign new_n1355_ = ~new_n1352_ & ~new_n1353_;
  assign new_n1356_ = new_n1354_ & new_n1355_;
  assign new_n1357_ = ng293 & new_n670_;
  assign new_n1358_ = ng536 & new_n682_;
  assign new_n1359_ = ng551 & new_n677_;
  assign new_n1360_ = ng508 & new_n681_;
  assign new_n1361_ = ~new_n1357_ & ~new_n1358_;
  assign new_n1362_ = ~new_n1359_ & ~new_n1360_;
  assign new_n1363_ = new_n1361_ & new_n1362_;
  assign new_n1364_ = ng692 & new_n701_;
  assign new_n1365_ = ~ng197 & ng692;
  assign new_n1366_ = ng206 & ~new_n736_;
  assign new_n1367_ = new_n735_ & ~new_n736_;
  assign new_n1368_ = ~new_n1366_ & ~new_n1367_;
  assign new_n1369_ = new_n752_ & ~new_n1368_;
  assign new_n1370_ = ~new_n742_ & new_n1369_;
  assign new_n1371_ = ng197 & new_n1370_;
  assign n694 = new_n1365_ | new_n1371_;
  assign new_n1373_ = new_n705_ & n694;
  assign new_n1374_ = new_n708_ & n319;
  assign new_n1375_ = new_n710_ & ~new_n1350_;
  assign new_n1376_ = ~new_n1364_ & ~new_n1373_;
  assign new_n1377_ = ~new_n1374_ & ~new_n1375_;
  assign new_n1378_ = new_n1376_ & new_n1377_;
  assign new_n1379_ = new_n1346_ & new_n1356_;
  assign new_n1380_ = new_n1363_ & new_n1378_;
  assign n629 = ~new_n1379_ | ~new_n1380_;
  assign new_n1382_ = ~ng269 & ng683;
  assign new_n1383_ = ng269 & ~new_n982_;
  assign n634 = new_n1382_ | new_n1383_;
  assign new_n1385_ = ~pg22 & ~n309;
  assign n639 = ng669 | new_n1385_;
  assign new_n1387_ = new_n519_1_ & pg6372;
  assign new_n1388_ = ng15 & ~new_n519_1_;
  assign n649 = new_n1387_ | new_n1388_;
  assign new_n1390_ = ng606 & ~new_n1095_;
  assign new_n1391_ = new_n1094_ & ~new_n1095_;
  assign new_n1392_ = ~new_n1390_ & ~new_n1391_;
  assign n659 = ng638 & ~new_n1392_;
  assign new_n1394_ = ng594 & ng590;
  assign new_n1395_ = ng590 & ~new_n1394_;
  assign new_n1396_ = ng594 & ~new_n1394_;
  assign new_n1397_ = ~new_n1395_ & ~new_n1396_;
  assign new_n1398_ = ng574 & ~ng590;
  assign new_n1399_ = ng594 & new_n1398_;
  assign new_n1400_ = ng582 & new_n1399_;
  assign new_n1401_ = ng578 & new_n1400_;
  assign new_n1402_ = ng586 & new_n1401_;
  assign new_n1403_ = ~new_n1397_ & ~new_n1402_;
  assign new_n1404_ = ng578 & ng677;
  assign new_n1405_ = ~ng578 & ng691;
  assign new_n1406_ = ~new_n1404_ & ~new_n1405_;
  assign new_n1407_ = ng582 & new_n1406_;
  assign new_n1408_ = ng578 & ng692;
  assign new_n1409_ = ~ng578 & ng680;
  assign new_n1410_ = ~new_n1408_ & ~new_n1409_;
  assign new_n1411_ = ~ng582 & new_n1410_;
  assign new_n1412_ = ~new_n1407_ & ~new_n1411_;
  assign new_n1413_ = ng586 & new_n1412_;
  assign new_n1414_ = ng578 & ng694;
  assign new_n1415_ = ~ng578 & ng682;
  assign new_n1416_ = ~new_n1414_ & ~new_n1415_;
  assign new_n1417_ = ng582 & new_n1416_;
  assign new_n1418_ = ng578 & ng683;
  assign new_n1419_ = ~ng578 & ng697;
  assign new_n1420_ = ~new_n1418_ & ~new_n1419_;
  assign new_n1421_ = ~ng582 & new_n1420_;
  assign new_n1422_ = ~new_n1417_ & ~new_n1421_;
  assign new_n1423_ = ~ng586 & new_n1422_;
  assign new_n1424_ = ~new_n1413_ & ~new_n1423_;
  assign new_n1425_ = ng574 & new_n1424_;
  assign new_n1426_ = ~ng574 & new_n1424_;
  assign new_n1427_ = ~new_n1425_ & ~new_n1426_;
  assign new_n1428_ = ~new_n1402_ & new_n1427_;
  assign n664 = new_n1403_ | new_n1428_;
  assign new_n1430_ = ng682 & new_n815_;
  assign new_n1431_ = ng520 & ~new_n815_;
  assign n669 = new_n1430_ | new_n1431_;
  assign new_n1433_ = ng680 & new_n580_;
  assign new_n1434_ = ng297 & ~new_n580_;
  assign n674 = new_n1433_ | new_n1434_;
  assign new_n1436_ = new_n519_1_ & pg6374;
  assign new_n1437_ = ng19 & ~new_n519_1_;
  assign n679 = new_n1436_ | new_n1437_;
  assign new_n1439_ = ng646 & ~new_n1096_;
  assign new_n1440_ = new_n1095_ & ~new_n1096_;
  assign new_n1441_ = ~new_n1439_ & ~new_n1440_;
  assign n689 = ng638 & ~new_n1441_;
  assign new_n1443_ = ~ng197 & ng697;
  assign new_n1444_ = ng197 & ~new_n919_;
  assign n699 = new_n1443_ | new_n1444_;
  assign new_n1446_ = ng680 & new_n1037_;
  assign new_n1447_ = ng465 & new_n787_;
  assign new_n1448_ = ~ng465 & new_n751_;
  assign new_n1449_ = ~new_n1447_ & ~new_n1448_;
  assign new_n1450_ = ~ng536 & ~new_n1449_;
  assign new_n1451_ = new_n627_ & new_n1450_;
  assign new_n1452_ = ~ng541 & ~new_n1451_;
  assign new_n1453_ = ~new_n1037_ & ~new_n1452_;
  assign n704 = new_n1446_ | new_n1453_;
  assign new_n1455_ = ~ng269 & ng697;
  assign new_n1456_ = ng269 & ~new_n986_;
  assign n709 = new_n1455_ | new_n1456_;
  assign new_n1458_ = ng642 & ~new_n1094_;
  assign new_n1459_ = new_n1093_ & ~new_n1094_;
  assign new_n1460_ = ~new_n1458_ & ~new_n1459_;
  assign n714 = ng638 & ~new_n1460_;
  assign new_n1462_ = ng610 & ~new_n831_;
  assign new_n1463_ = ng602 & ~new_n831_;
  assign new_n1464_ = ~new_n1462_ & ~new_n1463_;
  assign n719 = pg639 & ~new_n1464_;
  assign new_n1466_ = ng619 & ~new_n834_;
  assign new_n1467_ = new_n833_ & ~new_n834_;
  assign new_n1468_ = ~new_n1466_ & ~new_n1467_;
  assign n724 = pg639 & ~new_n1468_;
  assign new_n1470_ = ng586 & ~new_n841_;
  assign new_n1471_ = new_n840_ & ~new_n841_;
  assign new_n1472_ = ~new_n1470_ & ~new_n1471_;
  assign n734 = new_n845_ & ~new_n1472_;
  assign new_n1474_ = ng691 & new_n815_;
  assign new_n1475_ = ng504 & ~new_n815_;
  assign n739 = new_n1474_ | new_n1475_;
  assign new_n1477_ = ng613 & ~new_n832_;
  assign new_n1478_ = new_n831_ & ~new_n832_;
  assign new_n1479_ = ~new_n1477_ & ~new_n1478_;
  assign new_n1480_ = pg639 & ~new_n1479_;
  assign n744 = ~pg639 | new_n1480_;
  assign n749 = pg639 & ~ng602;
  assign new_n1483_ = ng631 & ~new_n838_;
  assign new_n1484_ = new_n837_ & ~new_n838_;
  assign new_n1485_ = ~new_n1483_ & ~new_n1484_;
  assign n759 = pg639 & ~new_n1485_;
  assign new_n1487_ = ng571 & new_n1340_;
  assign new_n1488_ = ng571 & ~new_n1487_;
  assign new_n1489_ = new_n1340_ & ~new_n1487_;
  assign new_n1490_ = ~new_n1488_ & ~new_n1489_;
  assign n769 = ng638 & ~new_n1490_;
  assign new_n1492_ = ng692 & new_n1037_;
  assign new_n1493_ = ng465 & ~new_n775_;
  assign new_n1494_ = ~ng465 & ~new_n739_1_;
  assign new_n1495_ = ~new_n1493_ & ~new_n1494_;
  assign new_n1496_ = new_n627_ & new_n1495_;
  assign new_n1497_ = ng536 & ~new_n1496_;
  assign new_n1498_ = ~new_n1037_ & new_n1497_;
  assign n774 = new_n1492_ | new_n1498_;
  assign new_n1500_ = new_n519_1_ & pg6366;
  assign new_n1501_ = ng33 & ~new_n519_1_;
  assign n779 = new_n1500_ | new_n1501_;
  assign new_n1503_ = ng461 & new_n629_1_;
  assign new_n1504_ = ng457 & ~new_n629_1_;
  assign n794 = new_n1503_ | new_n1504_;
  assign new_n1506_ = ng434 & new_n642_;
  assign new_n1507_ = ng677 & ng697;
  assign new_n1508_ = ~ng677 & ng697;
  assign new_n1509_ = ~new_n1507_ & ~new_n1508_;
  assign new_n1510_ = new_n649_1_ & ~new_n1509_;
  assign new_n1511_ = ng430 & new_n654_1_;
  assign new_n1512_ = ng697 & new_n658_;
  assign new_n1513_ = ~new_n1506_ & ~new_n1510_;
  assign new_n1514_ = ~new_n1511_ & ~new_n1512_;
  assign new_n1515_ = new_n1513_ & new_n1514_;
  assign new_n1516_ = pg557 & new_n667_;
  assign new_n1517_ = ng528 & new_n681_;
  assign new_n1518_ = ~new_n716_ & ~new_n1516_;
  assign new_n1519_ = ~new_n1517_ & new_n1518_;
  assign new_n1520_ = ng697 & new_n701_;
  assign new_n1521_ = new_n705_ & n699;
  assign new_n1522_ = new_n708_ & n709;
  assign new_n1523_ = new_n710_ & ~new_n1509_;
  assign new_n1524_ = ~new_n1520_ & ~new_n1521_;
  assign new_n1525_ = ~new_n1522_ & ~new_n1523_;
  assign new_n1526_ = new_n1524_ & new_n1525_;
  assign new_n1527_ = new_n1515_ & new_n1519_;
  assign n799 = ~new_n1526_ | ~new_n1527_;
  assign new_n1529_ = ng437 & new_n642_;
  assign new_n1530_ = ng677 & ng683;
  assign new_n1531_ = ~ng677 & ng683;
  assign new_n1532_ = ~new_n1530_ & ~new_n1531_;
  assign new_n1533_ = new_n649_1_ & ~new_n1532_;
  assign new_n1534_ = ng426 & new_n654_1_;
  assign new_n1535_ = ng683 & new_n658_;
  assign new_n1536_ = ~new_n1529_ & ~new_n1533_;
  assign new_n1537_ = ~new_n1534_ & ~new_n1535_;
  assign new_n1538_ = new_n1536_ & new_n1537_;
  assign new_n1539_ = pg558 & new_n667_;
  assign new_n1540_ = ng524 & new_n681_;
  assign new_n1541_ = ~new_n716_ & ~new_n1539_;
  assign new_n1542_ = ~new_n1540_ & new_n1541_;
  assign new_n1543_ = ng683 & new_n701_;
  assign new_n1544_ = new_n705_ & n284;
  assign new_n1545_ = new_n708_ & n634;
  assign new_n1546_ = new_n710_ & ~new_n1532_;
  assign new_n1547_ = ~new_n1543_ & ~new_n1544_;
  assign new_n1548_ = ~new_n1545_ & ~new_n1546_;
  assign new_n1549_ = new_n1547_ & new_n1548_;
  assign new_n1550_ = new_n1538_ & new_n1542_;
  assign n804 = ~new_n1549_ | ~new_n1550_;
  assign new_n1552_ = ng694 & new_n815_;
  assign new_n1553_ = ng516 & ~new_n815_;
  assign n809 = new_n1552_ | new_n1553_;
  assign new_n1555_ = ~new_n970_ & ~new_n976_;
  assign n819 = ng492 | ~new_n1555_;
  assign pg5692 = 1'b0;
  assign pg6728 = 1'b0;
  assign n194 = ~pg47;
  assign n444 = ~ng691;
  assign n564 = ~ng677;
  assign n764 = ~ng266;
  assign pg4098 = pg23;
  assign pg4108 = pg45;
  assign pg4109 = pg46;
  assign pg4307 = ng485;
  assign pg5137 = ng43;
  assign pg1293 = ng699;
  assign pg3222 = pg705;
  assign pg4104 = pg22;
  assign pg4105 = pg40;
  assign pg5469 = ng668;
  assign pg4106 = pg42;
  assign pg4107 = pg44;
  assign pg4422 = pg564;
  assign pg3600 = ng43;
  assign pg4100 = pg36;
  assign pg1290 = ng666;
  assign pg4099 = pg32;
  assign pg4101 = pg37;
  assign pg4110 = pg41;
  assign pg4321 = ng668;
  assign pg4102 = pg38;
  assign pg5468 = ng485;
  assign pg4103 = pg39;
  assign pg4112 = pg47;
  assign n154 = ng642;
  assign n204 = pg46;
  assign n239 = ng2;
  assign n259 = ng14;
  assign n289 = ng606;
  assign n294 = ng1;
  assign n349 = ng571;
  assign n354 = pg39;
  assign n359 = ng6;
  assign n414 = pg45;
  assign n419 = ng634;
  assign n429 = pg37;
  assign n434 = ng654;
  assign n464 = ng650;
  assign n469 = ng10;
  assign n499 = ng598;
  assign n524 = ng646;
  assign n544 = ng478;
  assign n574 = pg32;
  assign n589 = pg40;
  assign n599 = ng18;
  assign n624 = ng24;
  assign n644 = pg567;
  assign n654 = pg42;
  assign n729 = ng28;
  assign n784 = ng667;
  assign n789 = pg702;
  assign n814 = pg38;
  assign n824 = ng663;
  always @ (posedge clock) begin
    ng230 <= n154;
    ng197 <= n159;
    ng434 <= n164;
    ng25 <= n169;
    ng205 <= n174;
    ng266 <= n179;
    ng204 <= n184;
    ng524 <= n189;
    ng699 <= n194;
    ng658 <= n199;
    ng666 <= n204;
    ng414 <= n209;
    ng1 <= n214;
    ng598 <= n219;
    ng578 <= n224;
    ng406 <= n229;
    ng582 <= n234;
    ng691 <= n239;
    ng668 <= n244;
    ng548 <= n249;
    ng485 <= n254;
    ng694 <= n259;
    ng422 <= n264;
    ng500 <= n269;
    ng19 <= n274;
    ng532 <= n279;
    ng210 <= n284;
    ng236 <= n289;
    ng677 <= n294;
    ng512 <= n299;
    ng465 <= n304;
    ng676 <= n309;
    ng622 <= n314;
    ng278 <= n319;
    ng461 <= n324;
    ng650 <= n329;
    ng7 <= n334;
    ng18 <= n339;
    ng508 <= n344;
    ng260 <= n349;
    ng689 <= n354;
    ng692 <= n359;
    ng24 <= n364;
    ng277 <= n369;
    ng453 <= n374;
    ng445 <= n379;
    ng2 <= n384;
    ng279 <= n389;
    ng594 <= n394;
    ng269 <= n399;
    ng293 <= n404;
    ng628 <= n409;
    ng667 <= n414;
    ng286 <= n419;
    ng574 <= n424;
    ng687 <= n429;
    ng254 <= n434;
    ng672 <= n439;
    ng489 <= n444;
    ng207 <= n449;
    ng441 <= n454;
    ng6 <= n459;
    ng290 <= n464;
    ng680 <= n469;
    ng616 <= n474;
    ng554 <= n479;
    ng625 <= n484;
    ng426 <= n489;
    ng402 <= n494;
    ng218 <= n499;
    ng496 <= n504;
    ng208 <= n509;
    ng634 <= n514;
    ng418 <= n519;
    ng242 <= n524;
    ng48 <= n529;
    ng276 <= n534;
    ng449 <= n539;
    ng471 <= n544;
    ng590 <= n549;
    ng437 <= n554;
    ng528 <= n559;
    ng486 <= n564;
    ng551 <= n569;
    ng685 <= n574;
    ng281 <= n579;
    ng430 <= n584;
    ng698 <= n589;
    ng545 <= n594;
    ng682 <= n599;
    ng3 <= n604;
    ng15 <= n609;
    ng410 <= n614;
    ng654 <= n619;
    ng683 <= n624;
    ng11 <= n629;
    ng282 <= n634;
    ng669 <= n639;
    ng212 <= n644;
    ng10 <= n649;
    ng663 <= n654;
    ng606 <= n659;
    ng43 <= n664;
    ng520 <= n669;
    ng297 <= n674;
    ng14 <= n679;
    ng280 <= n684;
    ng646 <= n689;
    ng206 <= n694;
    ng211 <= n699;
    ng541 <= n704;
    ng283 <= n709;
    ng642 <= n714;
    ng610 <= n719;
    ng619 <= n724;
    ng697 <= n729;
    ng586 <= n734;
    ng504 <= n739;
    ng613 <= n744;
    ng602 <= n749;
    ng209 <= n754;
    ng631 <= n759;
    ng662 <= n764;
    ng571 <= n769;
    ng536 <= n774;
    ng28 <= n779;
    ng638 <= n784;
    ng675 <= n789;
    ng457 <= n794;
    ng33 <= n799;
    ng29 <= n804;
    ng516 <= n809;
    ng688 <= n814;
    ng492 <= n819;
    ng478 <= n824;
  end
endmodule

