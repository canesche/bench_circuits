module top ( clock, 
    c_6, c_5, c_4, c_19, c_3, c_29, c_2, c_1, c_0, ck, c_13, c_24, c_14,
    c_23, c_11, c_22, c_12, c_21, c_17, c_28, c_31, c_18, c_27, c_32, c_15,
    c_26, c_16, c_25, clear, c_30, c_20, c_10, x, c_9, c_8, c_7,
    w, z  );
  input  clock;
  input  c_6, c_5, c_4, c_19, c_3, c_29, c_2, c_1, c_0, ck, c_13, c_24,
    c_14, c_23, c_11, c_22, c_12, c_21, c_17, c_28, c_31, c_18, c_27, c_32,
    c_15, c_26, c_16, c_25, clear, c_30, c_20, c_10, x, c_9, c_8, c_7;
  output w, z;
  reg ny_4, ny_9, ny_22, ny_16, ny_23, ny_15, ny_28, ny_29, ny_14, ny_21,
    ny_8, ny_31, ny_1, ny_30, ny_2, ny_11, ny_24, ny_3, ny_10, ny_17,
    ny_12, ny_5, ny_6, ny_7, ny_13, ny_26, ny_20, ny_27, ny_19, ny_32,
    ny_18, ny_25;
  wire new_n135_, new_n136_, new_n138_1_, new_n139_, new_n140_, new_n141_,
    new_n142_, new_n143_1_, new_n144_, new_n145_, new_n146_, new_n147_,
    new_n148_1_, new_n149_, new_n150_, new_n151_, new_n152_, new_n153_1_,
    new_n154_, new_n155_, new_n156_, new_n157_, new_n158_1_, new_n159_,
    new_n160_, new_n161_, new_n162_, new_n163_1_, new_n164_, new_n165_,
    new_n166_, new_n167_, new_n168_1_, new_n169_, new_n170_, new_n171_,
    new_n172_, new_n173_1_, new_n174_, new_n175_, new_n176_, new_n177_,
    new_n178_1_, new_n179_, new_n180_, new_n181_, new_n182_, new_n183_1_,
    new_n184_, new_n185_, new_n186_, new_n187_, new_n188_1_, new_n189_,
    new_n190_, new_n191_, new_n192_, new_n193_1_, new_n194_, new_n195_,
    new_n196_, new_n197_, new_n198_1_, new_n199_, new_n200_, new_n201_,
    new_n202_, new_n203_1_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_1_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_1_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_1_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_1_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_1_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_1_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n266_, new_n267_, new_n268_,
    new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_,
    new_n276_, new_n277_, new_n278_, new_n279_, new_n281_, new_n282_,
    new_n283_, new_n284_, new_n286_, new_n287_, new_n288_, new_n290_,
    new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n309_, new_n310_,
    new_n311_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_,
    new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_,
    new_n325_, new_n326_, new_n329_, new_n330_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n348_,
    new_n349_, new_n351_, new_n352_, new_n354_, new_n355_, new_n356_,
    new_n357_, new_n358_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n365_, new_n366_, new_n367_, new_n369_, new_n370_, new_n372_,
    new_n373_, new_n375_, new_n376_, new_n377_, new_n378_, new_n381_,
    new_n382_, new_n384_, new_n385_, new_n386_, new_n389_, new_n390_,
    new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_,
    new_n399_, new_n400_, new_n401_, new_n403_, new_n404_, new_n405_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n412_, new_n413_, n78,
    n83, n88, n93, n98, n103, n108, n113, n118, n123, n128, n133, n138,
    n143, n148, n153, n158, n163, n168, n173, n178, n183, n188, n193, n198,
    n203, n208, n213, n218, n223, n228, n233;
  assign new_n135_ = ny_29 & ny_30;
  assign new_n136_ = ny_31 & new_n135_;
  assign w = ny_32 & new_n136_;
  assign new_n138_1_ = x & ~ny_1;
  assign new_n139_ = ~ny_2 & new_n138_1_;
  assign new_n140_ = ~ny_3 & new_n139_;
  assign new_n141_ = ~ny_4 & new_n140_;
  assign new_n142_ = ~ny_5 & new_n141_;
  assign new_n143_1_ = ~ny_6 & new_n142_;
  assign new_n144_ = ~ny_7 & new_n143_1_;
  assign new_n145_ = ~ny_8 & new_n144_;
  assign new_n146_ = ~ny_9 & new_n145_;
  assign new_n147_ = ~ny_10 & new_n146_;
  assign new_n148_1_ = ~ny_11 & new_n147_;
  assign new_n149_ = ny_12 & new_n148_1_;
  assign new_n150_ = c_12 & new_n149_;
  assign new_n151_ = ~ny_12 & new_n148_1_;
  assign new_n152_ = ~ny_13 & new_n151_;
  assign new_n153_1_ = ~ny_14 & new_n152_;
  assign new_n154_ = ~ny_15 & new_n153_1_;
  assign new_n155_ = ~ny_16 & new_n154_;
  assign new_n156_ = ~ny_17 & new_n155_;
  assign new_n157_ = ~ny_18 & new_n156_;
  assign new_n158_1_ = ~ny_19 & new_n157_;
  assign new_n159_ = ~ny_20 & new_n158_1_;
  assign new_n160_ = ~ny_21 & new_n159_;
  assign new_n161_ = ~ny_22 & new_n160_;
  assign new_n162_ = ~ny_23 & new_n161_;
  assign new_n163_1_ = ~ny_24 & new_n162_;
  assign new_n164_ = ~ny_25 & new_n163_1_;
  assign new_n165_ = ~ny_26 & new_n164_;
  assign new_n166_ = ny_27 & new_n165_;
  assign new_n167_ = c_27 & new_n166_;
  assign new_n168_1_ = ny_8 & new_n144_;
  assign new_n169_ = c_8 & new_n168_1_;
  assign new_n170_ = ~ny_27 & new_n165_;
  assign new_n171_ = ~ny_28 & new_n170_;
  assign new_n172_ = ny_29 & new_n171_;
  assign new_n173_1_ = c_29 & new_n172_;
  assign new_n174_ = ny_19 & new_n157_;
  assign new_n175_ = c_19 & new_n174_;
  assign new_n176_ = ~new_n173_1_ & ~new_n175_;
  assign new_n177_ = ny_7 & new_n143_1_;
  assign new_n178_1_ = c_7 & new_n177_;
  assign new_n179_ = new_n176_ & ~new_n178_1_;
  assign new_n180_ = ~new_n167_ & ~new_n169_;
  assign new_n181_ = new_n179_ & new_n180_;
  assign new_n182_ = ny_6 & new_n142_;
  assign new_n183_1_ = c_6 & new_n182_;
  assign new_n184_ = ny_21 & new_n159_;
  assign new_n185_ = c_21 & new_n184_;
  assign new_n186_ = ~new_n150_ & new_n181_;
  assign new_n187_ = ~new_n183_1_ & new_n186_;
  assign new_n188_1_ = ~new_n185_ & new_n187_;
  assign new_n189_ = c_0 & x;
  assign new_n190_ = ny_25 & new_n163_1_;
  assign new_n191_ = c_25 & new_n190_;
  assign new_n192_ = ~new_n189_ & ~new_n191_;
  assign new_n193_1_ = ny_2 & new_n138_1_;
  assign new_n194_ = c_2 & new_n193_1_;
  assign new_n195_ = ny_26 & new_n164_;
  assign new_n196_ = c_26 & new_n195_;
  assign new_n197_ = ~ny_29 & new_n171_;
  assign new_n198_1_ = ~ny_30 & new_n197_;
  assign new_n199_ = ~ny_31 & new_n198_1_;
  assign new_n200_ = ny_32 & new_n199_;
  assign new_n201_ = c_32 & new_n200_;
  assign new_n202_ = ny_24 & new_n162_;
  assign new_n203_1_ = c_24 & new_n202_;
  assign new_n204_ = ~new_n201_ & ~new_n203_1_;
  assign new_n205_ = ny_23 & new_n161_;
  assign new_n206_ = c_23 & new_n205_;
  assign new_n207_ = new_n204_ & ~new_n206_;
  assign new_n208_1_ = ny_14 & new_n152_;
  assign new_n209_ = c_14 & new_n208_1_;
  assign new_n210_ = new_n207_ & ~new_n209_;
  assign new_n211_ = ~new_n194_ & ~new_n196_;
  assign new_n212_ = new_n210_ & new_n211_;
  assign new_n213_1_ = ny_5 & new_n141_;
  assign new_n214_ = c_5 & new_n213_1_;
  assign new_n215_ = ny_16 & new_n154_;
  assign new_n216_ = c_16 & new_n215_;
  assign new_n217_ = ny_18 & new_n156_;
  assign new_n218_1_ = c_18 & new_n217_;
  assign new_n219_ = ny_20 & new_n158_1_;
  assign new_n220_ = c_20 & new_n219_;
  assign new_n221_ = ~new_n218_1_ & ~new_n220_;
  assign new_n222_ = ~new_n214_ & ~new_n216_;
  assign new_n223_1_ = new_n221_ & new_n222_;
  assign new_n224_ = ny_17 & new_n155_;
  assign new_n225_ = c_17 & new_n224_;
  assign new_n226_ = new_n192_ & new_n212_;
  assign new_n227_ = new_n223_1_ & new_n226_;
  assign new_n228_1_ = ~new_n225_ & new_n227_;
  assign new_n229_ = ny_9 & new_n145_;
  assign new_n230_ = c_9 & new_n229_;
  assign new_n231_ = ny_13 & new_n151_;
  assign new_n232_ = c_13 & new_n231_;
  assign new_n233_1_ = ny_30 & new_n197_;
  assign new_n234_ = c_30 & new_n233_1_;
  assign new_n235_ = ny_31 & new_n198_1_;
  assign new_n236_ = c_31 & new_n235_;
  assign new_n237_ = ~new_n234_ & ~new_n236_;
  assign new_n238_ = x & ny_1;
  assign new_n239_ = c_1 & new_n238_;
  assign new_n240_ = ny_4 & new_n140_;
  assign new_n241_ = c_4 & new_n240_;
  assign new_n242_ = ny_22 & new_n160_;
  assign new_n243_ = c_22 & new_n242_;
  assign new_n244_ = new_n237_ & ~new_n239_;
  assign new_n245_ = ~new_n241_ & new_n244_;
  assign new_n246_ = ~new_n243_ & new_n245_;
  assign new_n247_ = ~new_n230_ & ~new_n232_;
  assign new_n248_ = new_n246_ & new_n247_;
  assign new_n249_ = ny_3 & new_n139_;
  assign new_n250_ = c_3 & new_n249_;
  assign new_n251_ = ny_10 & new_n146_;
  assign new_n252_ = c_10 & new_n251_;
  assign new_n253_ = ny_11 & new_n147_;
  assign new_n254_ = c_11 & new_n253_;
  assign new_n255_ = ny_28 & new_n170_;
  assign new_n256_ = c_28 & new_n255_;
  assign new_n257_ = ny_15 & new_n153_1_;
  assign new_n258_ = c_15 & new_n257_;
  assign new_n259_ = ~new_n254_ & ~new_n256_;
  assign new_n260_ = ~new_n258_ & new_n259_;
  assign new_n261_ = ~new_n250_ & ~new_n252_;
  assign new_n262_ = new_n260_ & new_n261_;
  assign new_n263_ = new_n188_1_ & new_n228_1_;
  assign new_n264_ = new_n248_ & new_n263_;
  assign z = ~new_n262_ | ~new_n264_;
  assign new_n266_ = ~clear & x;
  assign new_n267_ = ny_1 & new_n266_;
  assign new_n268_ = ny_2 & new_n267_;
  assign new_n269_ = ~ny_4 & ny_3;
  assign new_n270_ = new_n268_ & new_n269_;
  assign new_n271_ = ny_1 & ny_2;
  assign new_n272_ = ny_3 & new_n271_;
  assign new_n273_ = new_n266_ & ~new_n272_;
  assign new_n274_ = ny_4 & new_n273_;
  assign n78 = new_n270_ | new_n274_;
  assign new_n276_ = ny_5 & ny_6;
  assign new_n277_ = ny_7 & new_n276_;
  assign new_n278_ = ny_8 & new_n277_;
  assign new_n279_ = ~clear & new_n278_;
  assign n83 = ~ny_9 & new_n279_;
  assign new_n281_ = ny_17 & ny_18;
  assign new_n282_ = ny_19 & new_n281_;
  assign new_n283_ = ny_20 & new_n282_;
  assign new_n284_ = ~clear & new_n283_;
  assign n123 = ~ny_21 & new_n284_;
  assign new_n286_ = ny_22 & n123;
  assign new_n287_ = ny_21 & new_n284_;
  assign new_n288_ = ~ny_22 & new_n287_;
  assign n88 = new_n286_ | new_n288_;
  assign new_n290_ = ny_9 & ny_10;
  assign new_n291_ = ny_11 & new_n290_;
  assign new_n292_ = ny_12 & new_n291_;
  assign new_n293_ = ~clear & new_n292_;
  assign new_n294_ = ny_13 & new_n293_;
  assign new_n295_ = ny_14 & new_n294_;
  assign new_n296_ = ~ny_16 & ny_15;
  assign new_n297_ = new_n295_ & new_n296_;
  assign new_n298_ = ny_14 & ny_13;
  assign new_n299_ = ny_15 & new_n298_;
  assign new_n300_ = new_n293_ & ~new_n299_;
  assign new_n301_ = ny_16 & new_n300_;
  assign n93 = new_n297_ | new_n301_;
  assign new_n303_ = ny_22 & ny_21;
  assign new_n304_ = new_n284_ & ~new_n303_;
  assign new_n305_ = ny_23 & new_n304_;
  assign new_n306_ = ny_22 & new_n287_;
  assign new_n307_ = ~ny_23 & new_n306_;
  assign n98 = new_n305_ | new_n307_;
  assign new_n309_ = new_n293_ & ~new_n298_;
  assign new_n310_ = ny_15 & new_n309_;
  assign new_n311_ = ~ny_15 & new_n295_;
  assign n103 = new_n310_ | new_n311_;
  assign new_n313_ = ny_23 & new_n303_;
  assign new_n314_ = ny_24 & new_n313_;
  assign new_n315_ = ~clear & new_n314_;
  assign new_n316_ = ny_25 & new_n315_;
  assign new_n317_ = ny_26 & new_n316_;
  assign new_n318_ = ~ny_28 & ny_27;
  assign new_n319_ = new_n317_ & new_n318_;
  assign new_n320_ = ny_26 & ny_25;
  assign new_n321_ = ny_27 & new_n320_;
  assign new_n322_ = new_n315_ & ~new_n321_;
  assign new_n323_ = ny_28 & new_n322_;
  assign n108 = new_n319_ | new_n323_;
  assign new_n325_ = ny_28 & new_n321_;
  assign new_n326_ = ~clear & new_n325_;
  assign n113 = ~ny_29 & new_n326_;
  assign n198 = ~ny_13 & new_n293_;
  assign new_n329_ = ny_14 & n198;
  assign new_n330_ = ~ny_14 & new_n294_;
  assign n118 = new_n329_ | new_n330_;
  assign new_n332_ = ny_4 & new_n272_;
  assign new_n333_ = ~clear & new_n332_;
  assign new_n334_ = ny_5 & new_n333_;
  assign new_n335_ = ny_6 & new_n334_;
  assign new_n336_ = ~ny_8 & ny_7;
  assign new_n337_ = new_n335_ & new_n336_;
  assign new_n338_ = ~new_n277_ & new_n333_;
  assign new_n339_ = ny_8 & new_n338_;
  assign n128 = new_n337_ | new_n339_;
  assign new_n341_ = ~new_n135_ & new_n326_;
  assign new_n342_ = ny_31 & new_n341_;
  assign new_n343_ = ny_29 & new_n326_;
  assign new_n344_ = ny_30 & new_n343_;
  assign new_n345_ = ~ny_31 & new_n344_;
  assign n133 = new_n342_ | new_n345_;
  assign n138 = ~ny_1 & new_n266_;
  assign new_n348_ = ny_30 & n113;
  assign new_n349_ = ~ny_30 & new_n343_;
  assign n143 = new_n348_ | new_n349_;
  assign new_n351_ = ny_2 & n138;
  assign new_n352_ = ~ny_2 & new_n267_;
  assign n148 = new_n351_ | new_n352_;
  assign new_n354_ = new_n279_ & ~new_n290_;
  assign new_n355_ = ny_11 & new_n354_;
  assign new_n356_ = ny_9 & new_n279_;
  assign new_n357_ = ny_10 & new_n356_;
  assign new_n358_ = ~ny_11 & new_n357_;
  assign n153 = new_n355_ | new_n358_;
  assign new_n360_ = ny_23 & ~ny_24;
  assign new_n361_ = new_n306_ & new_n360_;
  assign new_n362_ = new_n284_ & ~new_n313_;
  assign new_n363_ = ny_24 & new_n362_;
  assign n158 = new_n361_ | new_n363_;
  assign new_n365_ = new_n266_ & ~new_n271_;
  assign new_n366_ = ny_3 & new_n365_;
  assign new_n367_ = ~ny_3 & new_n268_;
  assign n163 = new_n366_ | new_n367_;
  assign new_n369_ = ny_10 & n83;
  assign new_n370_ = ~ny_10 & new_n356_;
  assign n168 = new_n369_ | new_n370_;
  assign new_n372_ = ny_16 & new_n299_;
  assign new_n373_ = ~clear & new_n372_;
  assign n173 = ~ny_17 & new_n373_;
  assign new_n375_ = ny_11 & ~ny_12;
  assign new_n376_ = new_n357_ & new_n375_;
  assign new_n377_ = new_n279_ & ~new_n291_;
  assign new_n378_ = ny_12 & new_n377_;
  assign n178 = new_n376_ | new_n378_;
  assign n183 = ~ny_5 & new_n333_;
  assign new_n381_ = ny_6 & n183;
  assign new_n382_ = ~ny_6 & new_n334_;
  assign n188 = new_n381_ | new_n382_;
  assign new_n384_ = ~new_n276_ & new_n333_;
  assign new_n385_ = ny_7 & new_n384_;
  assign new_n386_ = ~ny_7 & new_n335_;
  assign n193 = new_n385_ | new_n386_;
  assign n233 = ~ny_25 & new_n315_;
  assign new_n389_ = ny_26 & n233;
  assign new_n390_ = ~ny_26 & new_n316_;
  assign n203 = new_n389_ | new_n390_;
  assign new_n392_ = ny_17 & new_n373_;
  assign new_n393_ = ny_18 & new_n392_;
  assign new_n394_ = ~ny_20 & ny_19;
  assign new_n395_ = new_n393_ & new_n394_;
  assign new_n396_ = ~new_n282_ & new_n373_;
  assign new_n397_ = ny_20 & new_n396_;
  assign n208 = new_n395_ | new_n397_;
  assign new_n399_ = new_n315_ & ~new_n320_;
  assign new_n400_ = ny_27 & new_n399_;
  assign new_n401_ = ~ny_27 & new_n317_;
  assign n213 = new_n400_ | new_n401_;
  assign new_n403_ = ~new_n281_ & new_n373_;
  assign new_n404_ = ny_19 & new_n403_;
  assign new_n405_ = ~ny_19 & new_n393_;
  assign n218 = new_n404_ | new_n405_;
  assign new_n407_ = ny_31 & ~ny_32;
  assign new_n408_ = new_n344_ & new_n407_;
  assign new_n409_ = ~new_n136_ & new_n326_;
  assign new_n410_ = ny_32 & new_n409_;
  assign n223 = new_n408_ | new_n410_;
  assign new_n412_ = ny_18 & n173;
  assign new_n413_ = ~ny_18 & new_n392_;
  assign n228 = new_n412_ | new_n413_;
  always @ (posedge clock) begin
    ny_4 <= n78;
    ny_9 <= n83;
    ny_22 <= n88;
    ny_16 <= n93;
    ny_23 <= n98;
    ny_15 <= n103;
    ny_28 <= n108;
    ny_29 <= n113;
    ny_14 <= n118;
    ny_21 <= n123;
    ny_8 <= n128;
    ny_31 <= n133;
    ny_1 <= n138;
    ny_30 <= n143;
    ny_2 <= n148;
    ny_11 <= n153;
    ny_24 <= n158;
    ny_3 <= n163;
    ny_10 <= n168;
    ny_17 <= n173;
    ny_12 <= n178;
    ny_5 <= n183;
    ny_6 <= n188;
    ny_7 <= n193;
    ny_13 <= n198;
    ny_26 <= n203;
    ny_20 <= n208;
    ny_27 <= n213;
    ny_19 <= n218;
    ny_32 <= n223;
    ny_18 <= n228;
    ny_25 <= n233;
  end
endmodule

