module f51m ( 
    \1 , 2, 3, 4, 5, 6, 7, 8,
    44, 45, 46, 47, 48, 49, 50, 51  );
  input  \1 , 2, 3, 4, 5, 6, 7, 8;
  output 44, 45, 46, 47, 48, 49, 50, 51;
  wire new_n17_, new_n18_, new_n19_, new_n20_, new_n21_, new_n22_, new_n23_,
    new_n24_, new_n25_, new_n26_, new_n27_, new_n28_, new_n29_, new_n30_,
    new_n31_, new_n32_, new_n33_, new_n34_, new_n35_, new_n36_, new_n37_,
    new_n38_, new_n39_, new_n40_, new_n41_, new_n42_, new_n43_, new_n44_,
    new_n45_, new_n46_, new_n47_, new_n48_, new_n49_, new_n50_, new_n51_,
    new_n52_, new_n53_, new_n54_, new_n55_, new_n56_, new_n57_, new_n58_,
    new_n59_, new_n60_, new_n61_, new_n62_, new_n63_, new_n64_, new_n65_,
    new_n67_, new_n68_, new_n69_, new_n70_, new_n71_, new_n72_, new_n73_,
    new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_, new_n80_,
    new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_, new_n87_,
    new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_, new_n94_,
    new_n95_, new_n96_, new_n97_, new_n98_, new_n100_, new_n101_,
    new_n102_, new_n103_, new_n104_, new_n105_, new_n106_, new_n107_,
    new_n108_, new_n109_, new_n110_, new_n111_, new_n112_, new_n113_,
    new_n114_, new_n115_, new_n116_, new_n117_, new_n118_, new_n119_,
    new_n120_, new_n121_, new_n122_, new_n123_, new_n124_, new_n125_,
    new_n126_, new_n127_, new_n128_, new_n130_, new_n131_, new_n132_,
    new_n133_, new_n134_, new_n135_, new_n136_, new_n137_, new_n138_,
    new_n139_, new_n140_, new_n141_, new_n142_, new_n144_, new_n145_,
    new_n146_, new_n147_, new_n148_, new_n149_, new_n150_, new_n152_,
    new_n153_;
  assign new_n17_ = 2 & 6;
  assign new_n18_ = ~4 & ~new_n17_;
  assign new_n19_ = ~3 & 5;
  assign new_n20_ = ~\1  & new_n19_;
  assign new_n21_ = 3 & 8;
  assign new_n22_ = \1  & new_n21_;
  assign new_n23_ = ~new_n20_ & ~new_n22_;
  assign new_n24_ = ~new_n18_ & ~new_n23_;
  assign new_n25_ = 7 & new_n24_;
  assign new_n26_ = 6 & 8;
  assign new_n27_ = 5 & new_n26_;
  assign new_n28_ = ~4 & ~new_n27_;
  assign new_n29_ = 2 & ~new_n28_;
  assign new_n30_ = 5 & 6;
  assign new_n31_ = 4 & new_n30_;
  assign new_n32_ = ~new_n29_ & ~new_n31_;
  assign new_n33_ = ~3 & ~new_n32_;
  assign new_n34_ = 7 & 8;
  assign new_n35_ = ~2 & ~6;
  assign new_n36_ = 4 & ~new_n35_;
  assign new_n37_ = ~new_n34_ & ~new_n36_;
  assign new_n38_ = ~4 & ~6;
  assign new_n39_ = ~new_n37_ & ~new_n38_;
  assign new_n40_ = ~5 & ~new_n39_;
  assign new_n41_ = ~2 & ~4;
  assign new_n42_ = ~new_n40_ & ~new_n41_;
  assign new_n43_ = 3 & ~new_n42_;
  assign new_n44_ = ~new_n33_ & ~new_n43_;
  assign new_n45_ = ~\1  & ~new_n44_;
  assign new_n46_ = ~4 & ~5;
  assign new_n47_ = 2 & ~new_n46_;
  assign new_n48_ = ~5 & ~6;
  assign new_n49_ = 4 & ~new_n48_;
  assign new_n50_ = ~new_n47_ & ~new_n49_;
  assign new_n51_ = 3 & ~new_n50_;
  assign new_n52_ = 2 & 4;
  assign new_n53_ = ~5 & ~new_n52_;
  assign new_n54_ = ~6 & ~7;
  assign new_n55_ = 4 & ~new_n54_;
  assign new_n56_ = ~2 & ~new_n55_;
  assign new_n57_ = ~7 & ~8;
  assign new_n58_ = 6 & ~new_n57_;
  assign new_n59_ = ~4 & ~new_n58_;
  assign new_n60_ = ~new_n56_ & ~new_n59_;
  assign new_n61_ = ~new_n53_ & new_n60_;
  assign new_n62_ = ~3 & ~new_n61_;
  assign new_n63_ = ~new_n51_ & ~new_n62_;
  assign new_n64_ = \1  & ~new_n63_;
  assign new_n65_ = ~new_n45_ & ~new_n64_;
  assign 44 = new_n25_ | ~new_n65_;
  assign new_n67_ = 6 & new_n34_;
  assign new_n68_ = ~5 & ~new_n67_;
  assign new_n69_ = 3 & ~new_n68_;
  assign new_n70_ = 5 & new_n58_;
  assign new_n71_ = ~new_n69_ & ~new_n70_;
  assign new_n72_ = ~2 & ~new_n71_;
  assign new_n73_ = ~3 & ~8;
  assign new_n74_ = 5 & ~new_n73_;
  assign new_n75_ = ~7 & ~new_n74_;
  assign new_n76_ = ~3 & ~new_n30_;
  assign new_n77_ = ~5 & ~8;
  assign new_n78_ = ~new_n76_ & ~new_n77_;
  assign new_n79_ = ~new_n75_ & new_n78_;
  assign new_n80_ = 2 & ~new_n79_;
  assign new_n81_ = ~new_n72_ & ~new_n80_;
  assign new_n82_ = ~4 & ~new_n81_;
  assign new_n83_ = 3 & ~new_n48_;
  assign new_n84_ = 5 & ~new_n54_;
  assign new_n85_ = ~new_n83_ & ~new_n84_;
  assign new_n86_ = 2 & ~new_n85_;
  assign new_n87_ = ~3 & ~new_n84_;
  assign new_n88_ = ~6 & ~new_n34_;
  assign new_n89_ = ~5 & new_n88_;
  assign new_n90_ = ~new_n87_ & ~new_n89_;
  assign new_n91_ = ~2 & ~new_n90_;
  assign new_n92_ = ~new_n86_ & ~new_n91_;
  assign new_n93_ = 4 & ~new_n92_;
  assign new_n94_ = 3 & ~5;
  assign new_n95_ = 2 & new_n94_;
  assign new_n96_ = ~6 & new_n34_;
  assign new_n97_ = new_n95_ & new_n96_;
  assign new_n98_ = ~new_n93_ & ~new_n97_;
  assign 45 = new_n82_ | ~new_n98_;
  assign new_n100_ = 3 & 5;
  assign new_n101_ = ~5 & 8;
  assign new_n102_ = ~3 & new_n101_;
  assign new_n103_ = ~new_n100_ & ~new_n102_;
  assign new_n104_ = ~new_n38_ & ~new_n103_;
  assign new_n105_ = 7 & new_n104_;
  assign new_n106_ = 4 & 5;
  assign new_n107_ = ~7 & 8;
  assign new_n108_ = ~4 & new_n107_;
  assign new_n109_ = ~new_n106_ & ~new_n108_;
  assign new_n110_ = 3 & ~new_n109_;
  assign new_n111_ = 4 & ~5;
  assign new_n112_ = ~3 & new_n111_;
  assign new_n113_ = ~new_n110_ & ~new_n112_;
  assign new_n114_ = 6 & ~new_n113_;
  assign new_n115_ = ~5 & ~new_n26_;
  assign new_n116_ = 3 & new_n115_;
  assign new_n117_ = 5 & ~new_n58_;
  assign new_n118_ = ~3 & new_n117_;
  assign new_n119_ = ~new_n116_ & ~new_n118_;
  assign new_n120_ = ~4 & ~new_n119_;
  assign new_n121_ = ~5 & ~new_n34_;
  assign new_n122_ = 3 & new_n121_;
  assign new_n123_ = 5 & ~7;
  assign new_n124_ = ~3 & new_n123_;
  assign new_n125_ = ~new_n122_ & ~new_n124_;
  assign new_n126_ = ~6 & ~new_n125_;
  assign new_n127_ = ~new_n120_ & ~new_n126_;
  assign new_n128_ = ~new_n114_ & new_n127_;
  assign 46 = new_n105_ | ~new_n128_;
  assign new_n130_ = 6 & 7;
  assign new_n131_ = ~new_n107_ & ~new_n130_;
  assign new_n132_ = 5 & ~new_n131_;
  assign new_n133_ = 7 & ~new_n77_;
  assign new_n134_ = ~6 & ~new_n133_;
  assign new_n135_ = ~new_n67_ & ~new_n134_;
  assign new_n136_ = ~new_n132_ & new_n135_;
  assign new_n137_ = 4 & ~new_n136_;
  assign new_n138_ = ~new_n57_ & ~new_n121_;
  assign new_n139_ = 6 & ~new_n138_;
  assign new_n140_ = ~6 & new_n133_;
  assign new_n141_ = ~new_n139_ & ~new_n140_;
  assign new_n142_ = ~4 & ~new_n141_;
  assign 47 = new_n137_ | new_n142_;
  assign new_n144_ = 6 & new_n107_;
  assign new_n145_ = 7 & ~8;
  assign new_n146_ = ~new_n144_ & ~new_n145_;
  assign new_n147_ = ~5 & ~new_n146_;
  assign new_n148_ = ~7 & ~new_n26_;
  assign new_n149_ = ~new_n34_ & ~new_n148_;
  assign new_n150_ = 5 & ~new_n149_;
  assign 48 = new_n147_ | new_n150_;
  assign new_n152_ = 6 & ~new_n107_;
  assign new_n153_ = ~6 & new_n107_;
  assign 49 = new_n152_ | new_n153_;
  assign 50 = new_n107_ | new_n145_;
  assign 51 = ~8;
endmodule

